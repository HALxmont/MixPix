magic
tech sky130A
magscale 1 2
timestamp 1668295095
<< viali >>
rect 1961 57545 1995 57579
rect 3893 57545 3927 57579
rect 5089 57545 5123 57579
rect 6653 57545 6687 57579
rect 8217 57545 8251 57579
rect 9781 57545 9815 57579
rect 11621 57545 11655 57579
rect 12909 57545 12943 57579
rect 14473 57545 14507 57579
rect 16773 57545 16807 57579
rect 17693 57545 17727 57579
rect 19441 57545 19475 57579
rect 20821 57545 20855 57579
rect 22385 57545 22419 57579
rect 24593 57545 24627 57579
rect 25513 57545 25547 57579
rect 27169 57545 27203 57579
rect 28641 57545 28675 57579
rect 30205 57545 30239 57579
rect 32321 57545 32355 57579
rect 33333 57545 33367 57579
rect 34897 57545 34931 57579
rect 36461 57545 36495 57579
rect 38025 57545 38059 57579
rect 40049 57545 40083 57579
rect 41153 57545 41187 57579
rect 42717 57545 42751 57579
rect 44281 57545 44315 57579
rect 45845 57545 45879 57579
rect 47777 57545 47811 57579
rect 2145 57409 2179 57443
rect 4077 57409 4111 57443
rect 5273 57409 5307 57443
rect 6837 57409 6871 57443
rect 8401 57409 8435 57443
rect 9965 57409 9999 57443
rect 11805 57409 11839 57443
rect 13093 57409 13127 57443
rect 14657 57409 14691 57443
rect 16957 57409 16991 57443
rect 17509 57409 17543 57443
rect 19257 57409 19291 57443
rect 20637 57409 20671 57443
rect 22201 57409 22235 57443
rect 24409 57409 24443 57443
rect 25329 57409 25363 57443
rect 26985 57409 27019 57443
rect 28457 57409 28491 57443
rect 30021 57409 30055 57443
rect 32137 57409 32171 57443
rect 33149 57409 33183 57443
rect 34713 57409 34747 57443
rect 36277 57409 36311 57443
rect 37841 57409 37875 57443
rect 39865 57409 39899 57443
rect 40969 57409 41003 57443
rect 42533 57409 42567 57443
rect 44097 57409 44131 57443
rect 45661 57409 45695 57443
rect 47593 57409 47627 57443
rect 48789 57409 48823 57443
rect 50353 57409 50387 57443
rect 51917 57409 51951 57443
rect 53481 57409 53515 57443
rect 56609 57409 56643 57443
rect 57989 57409 58023 57443
rect 55321 57341 55355 57375
rect 2697 57205 2731 57239
rect 18705 57205 18739 57239
rect 20085 57205 20119 57239
rect 18705 57001 18739 57035
rect 19533 57001 19567 57035
rect 19993 57001 20027 57035
rect 57529 57001 57563 57035
rect 1409 56797 1443 56831
rect 17509 56797 17543 56831
rect 18521 56797 18555 56831
rect 19349 56797 19383 56831
rect 20177 56797 20211 56831
rect 58173 56797 58207 56831
rect 18061 56729 18095 56763
rect 42349 56729 42383 56763
rect 20729 56661 20763 56695
rect 40785 56661 40819 56695
rect 13553 56457 13587 56491
rect 15761 56457 15795 56491
rect 17509 56457 17543 56491
rect 18797 56457 18831 56491
rect 21281 56457 21315 56491
rect 22753 56457 22787 56491
rect 24685 56457 24719 56491
rect 25329 56457 25363 56491
rect 26433 56457 26467 56491
rect 27169 56457 27203 56491
rect 28733 56457 28767 56491
rect 31309 56457 31343 56491
rect 32321 56457 32355 56491
rect 35725 56457 35759 56491
rect 44005 56457 44039 56491
rect 46305 56457 46339 56491
rect 17049 56389 17083 56423
rect 13737 56321 13771 56355
rect 15945 56321 15979 56355
rect 17693 56321 17727 56355
rect 18337 56321 18371 56355
rect 18981 56321 19015 56355
rect 19625 56321 19659 56355
rect 20269 56321 20303 56355
rect 21097 56321 21131 56355
rect 21925 56321 21959 56355
rect 22569 56321 22603 56355
rect 23213 56321 23247 56355
rect 23857 56321 23891 56355
rect 24501 56321 24535 56355
rect 25145 56321 25179 56355
rect 26249 56321 26283 56355
rect 26985 56321 27019 56355
rect 28549 56321 28583 56355
rect 29193 56321 29227 56355
rect 30481 56321 30515 56355
rect 31125 56321 31159 56355
rect 32137 56321 32171 56355
rect 32781 56321 32815 56355
rect 35541 56321 35575 56355
rect 36185 56321 36219 56355
rect 43821 56321 43855 56355
rect 44465 56321 44499 56355
rect 46121 56321 46155 56355
rect 58173 56321 58207 56355
rect 18153 56185 18187 56219
rect 19441 56185 19475 56219
rect 22109 56185 22143 56219
rect 29929 56185 29963 56219
rect 30665 56185 30699 56219
rect 14197 56117 14231 56151
rect 20085 56117 20119 56151
rect 23397 56117 23431 56151
rect 24041 56117 24075 56151
rect 27997 56117 28031 56151
rect 29377 56117 29411 56151
rect 46765 56117 46799 56151
rect 17509 55845 17543 55879
rect 18521 55845 18555 55879
rect 19625 55845 19659 55879
rect 22385 55777 22419 55811
rect 1409 55709 1443 55743
rect 17693 55709 17727 55743
rect 18705 55709 18739 55743
rect 19809 55709 19843 55743
rect 16129 55573 16163 55607
rect 17049 55573 17083 55607
rect 20269 55573 20303 55607
rect 20913 55573 20947 55607
rect 21741 55573 21775 55607
rect 23029 55573 23063 55607
rect 23765 55573 23799 55607
rect 24409 55573 24443 55607
rect 25053 55573 25087 55607
rect 26065 55573 26099 55607
rect 26801 55573 26835 55607
rect 29561 55573 29595 55607
rect 30941 55573 30975 55607
rect 17785 55301 17819 55335
rect 18797 55301 18831 55335
rect 19809 55301 19843 55335
rect 58173 55097 58207 55131
rect 1409 54621 1443 54655
rect 58173 53941 58207 53975
rect 1409 53533 1443 53567
rect 1409 52445 1443 52479
rect 58173 52445 58207 52479
rect 1409 51357 1443 51391
rect 58173 51357 58207 51391
rect 1409 50269 1443 50303
rect 58173 49725 58207 49759
rect 1409 49181 1443 49215
rect 58173 48501 58207 48535
rect 1409 48093 1443 48127
rect 58173 47005 58207 47039
rect 58173 45917 58207 45951
rect 58173 44217 58207 44251
rect 58173 43061 58207 43095
rect 16589 42517 16623 42551
rect 16681 42177 16715 42211
rect 16865 42177 16899 42211
rect 17049 41973 17083 42007
rect 17785 41973 17819 42007
rect 18613 41701 18647 41735
rect 14381 41565 14415 41599
rect 14473 41565 14507 41599
rect 14565 41565 14599 41599
rect 14749 41565 14783 41599
rect 15853 41565 15887 41599
rect 16037 41565 16071 41599
rect 16129 41565 16163 41599
rect 16221 41565 16255 41599
rect 16957 41565 16991 41599
rect 17141 41565 17175 41599
rect 17233 41565 17267 41599
rect 17325 41565 17359 41599
rect 19441 41565 19475 41599
rect 58173 41565 58207 41599
rect 12817 41497 12851 41531
rect 13001 41497 13035 41531
rect 19257 41497 19291 41531
rect 19625 41497 19659 41531
rect 10333 41429 10367 41463
rect 12633 41429 12667 41463
rect 13553 41429 13587 41463
rect 14105 41429 14139 41463
rect 15301 41429 15335 41463
rect 16497 41429 16531 41463
rect 17601 41429 17635 41463
rect 20085 41429 20119 41463
rect 17049 41225 17083 41259
rect 20821 41225 20855 41259
rect 10241 41157 10275 41191
rect 15209 41157 15243 41191
rect 16681 41157 16715 41191
rect 20177 41157 20211 41191
rect 6653 41089 6687 41123
rect 6742 41092 6776 41126
rect 6858 41089 6892 41123
rect 7021 41089 7055 41123
rect 10425 41089 10459 41123
rect 12909 41089 12943 41123
rect 13001 41089 13035 41123
rect 13093 41089 13127 41123
rect 13277 41089 13311 41123
rect 14013 41089 14047 41123
rect 14105 41089 14139 41123
rect 14197 41089 14231 41123
rect 14381 41089 14415 41123
rect 15025 41089 15059 41123
rect 16865 41089 16899 41123
rect 17785 41089 17819 41123
rect 17969 41089 18003 41123
rect 18061 41089 18095 41123
rect 18153 41089 18187 41123
rect 18889 41089 18923 41123
rect 19073 41089 19107 41123
rect 19165 41092 19199 41126
rect 19257 41089 19291 41123
rect 20361 41089 20395 41123
rect 14841 41021 14875 41055
rect 19993 41021 20027 41055
rect 22661 40953 22695 40987
rect 6377 40885 6411 40919
rect 7573 40885 7607 40919
rect 10609 40885 10643 40919
rect 12633 40885 12667 40919
rect 13737 40885 13771 40919
rect 15669 40885 15703 40919
rect 18429 40885 18463 40919
rect 19533 40885 19567 40919
rect 23213 40885 23247 40919
rect 13553 40681 13587 40715
rect 18613 40681 18647 40715
rect 10701 40545 10735 40579
rect 14381 40545 14415 40579
rect 3801 40477 3835 40511
rect 6101 40477 6135 40511
rect 6368 40477 6402 40511
rect 9873 40477 9907 40511
rect 9962 40474 9996 40508
rect 10057 40477 10091 40511
rect 10241 40477 10275 40511
rect 10968 40477 11002 40511
rect 13369 40477 13403 40511
rect 14105 40477 14139 40511
rect 16129 40477 16163 40511
rect 16396 40477 16430 40511
rect 19257 40477 19291 40511
rect 19524 40477 19558 40511
rect 22109 40477 22143 40511
rect 22201 40477 22235 40511
rect 22293 40477 22327 40511
rect 22477 40477 22511 40511
rect 23213 40477 23247 40511
rect 27353 40477 27387 40511
rect 31217 40477 31251 40511
rect 58173 40477 58207 40511
rect 3985 40409 4019 40443
rect 13185 40409 13219 40443
rect 23029 40409 23063 40443
rect 27620 40409 27654 40443
rect 31484 40409 31518 40443
rect 4169 40341 4203 40375
rect 7481 40341 7515 40375
rect 9597 40341 9631 40375
rect 12081 40341 12115 40375
rect 12633 40341 12667 40375
rect 17509 40341 17543 40375
rect 20637 40341 20671 40375
rect 21833 40341 21867 40375
rect 23397 40341 23431 40375
rect 28733 40341 28767 40375
rect 32597 40341 32631 40375
rect 3985 40137 4019 40171
rect 8769 40137 8803 40171
rect 12173 40137 12207 40171
rect 12817 40137 12851 40171
rect 16681 40137 16715 40171
rect 19901 40137 19935 40171
rect 27629 40137 27663 40171
rect 6929 40069 6963 40103
rect 9496 40069 9530 40103
rect 18766 40069 18800 40103
rect 20913 40069 20947 40103
rect 28917 40069 28951 40103
rect 29101 40069 29135 40103
rect 2872 40001 2906 40035
rect 6561 40001 6595 40035
rect 6745 40001 6779 40035
rect 7389 40001 7423 40035
rect 7656 40001 7690 40035
rect 11529 40001 11563 40035
rect 11713 40001 11747 40035
rect 11808 40001 11842 40035
rect 11897 40001 11931 40035
rect 13941 40001 13975 40035
rect 17794 40001 17828 40035
rect 21097 40001 21131 40035
rect 21281 40001 21315 40035
rect 22477 40001 22511 40035
rect 22661 40001 22695 40035
rect 22753 40001 22787 40035
rect 22891 40001 22925 40035
rect 24694 40001 24728 40035
rect 27859 40001 27893 40035
rect 27997 40001 28031 40035
rect 28110 40001 28144 40035
rect 28273 40001 28307 40035
rect 2605 39933 2639 39967
rect 9229 39933 9263 39967
rect 14197 39933 14231 39967
rect 18061 39933 18095 39967
rect 18521 39933 18555 39967
rect 23121 39933 23155 39967
rect 24961 39933 24995 39967
rect 28733 39933 28767 39967
rect 10609 39797 10643 39831
rect 14657 39797 14691 39831
rect 23581 39797 23615 39831
rect 27077 39797 27111 39831
rect 3801 39593 3835 39627
rect 11437 39593 11471 39627
rect 12173 39593 12207 39627
rect 31493 39593 31527 39627
rect 4905 39525 4939 39559
rect 32321 39525 32355 39559
rect 5549 39457 5583 39491
rect 13553 39457 13587 39491
rect 22385 39457 22419 39491
rect 4077 39389 4111 39423
rect 4169 39389 4203 39423
rect 4261 39389 4295 39423
rect 4445 39389 4479 39423
rect 7389 39389 7423 39423
rect 7665 39389 7699 39423
rect 9229 39389 9263 39423
rect 11069 39389 11103 39423
rect 11253 39389 11287 39423
rect 14105 39389 14139 39423
rect 14381 39389 14415 39423
rect 23029 39389 23063 39423
rect 23213 39389 23247 39423
rect 23305 39389 23339 39423
rect 23397 39389 23431 39423
rect 24409 39389 24443 39423
rect 27261 39389 27295 39423
rect 30849 39389 30883 39423
rect 31028 39386 31062 39420
rect 31125 39389 31159 39423
rect 31263 39389 31297 39423
rect 5816 39321 5850 39355
rect 9496 39321 9530 39355
rect 13308 39321 13342 39355
rect 22118 39321 22152 39355
rect 23673 39321 23707 39355
rect 24654 39321 24688 39355
rect 27528 39321 27562 39355
rect 31953 39321 31987 39355
rect 32137 39321 32171 39355
rect 6929 39253 6963 39287
rect 10609 39253 10643 39287
rect 16865 39253 16899 39287
rect 21005 39253 21039 39287
rect 25789 39253 25823 39287
rect 28641 39253 28675 39287
rect 30389 39253 30423 39287
rect 9965 39049 9999 39083
rect 13093 39049 13127 39083
rect 18337 39049 18371 39083
rect 22845 39049 22879 39083
rect 27537 39049 27571 39083
rect 2688 38981 2722 39015
rect 4261 38981 4295 39015
rect 5457 38981 5491 39015
rect 11529 38981 11563 39015
rect 23213 38981 23247 39015
rect 2421 38913 2455 38947
rect 4491 38913 4525 38947
rect 4629 38913 4663 38947
rect 4742 38913 4776 38947
rect 4905 38913 4939 38947
rect 6377 38913 6411 38947
rect 6561 38913 6595 38947
rect 10221 38913 10255 38947
rect 10346 38916 10380 38950
rect 10446 38913 10480 38947
rect 10609 38913 10643 38947
rect 12909 38913 12943 38947
rect 17049 38913 17083 38947
rect 23029 38913 23063 38947
rect 26985 38913 27019 38947
rect 27793 38913 27827 38947
rect 27905 38913 27939 38947
rect 27997 38913 28031 38947
rect 28181 38913 28215 38947
rect 7849 38845 7883 38879
rect 8125 38845 8159 38879
rect 58173 38777 58207 38811
rect 3801 38709 3835 38743
rect 6745 38709 6779 38743
rect 8585 38709 8619 38743
rect 23857 38709 23891 38743
rect 29653 38709 29687 38743
rect 4169 38505 4203 38539
rect 6101 38505 6135 38539
rect 28089 38505 28123 38539
rect 16313 38437 16347 38471
rect 30941 38369 30975 38403
rect 2881 38301 2915 38335
rect 2973 38301 3007 38335
rect 3065 38301 3099 38335
rect 3249 38301 3283 38335
rect 6357 38301 6391 38335
rect 6466 38301 6500 38335
rect 6561 38301 6595 38335
rect 6745 38301 6779 38335
rect 15761 38301 15795 38335
rect 16037 38301 16071 38335
rect 16129 38301 16163 38335
rect 16773 38301 16807 38335
rect 17049 38301 17083 38335
rect 17141 38301 17175 38335
rect 19349 38301 19383 38335
rect 19442 38301 19476 38335
rect 19855 38301 19889 38335
rect 24593 38301 24627 38335
rect 28273 38301 28307 38335
rect 31585 38301 31619 38335
rect 3801 38233 3835 38267
rect 3985 38233 4019 38267
rect 9321 38233 9355 38267
rect 15945 38233 15979 38267
rect 16957 38233 16991 38267
rect 19625 38233 19659 38267
rect 19717 38233 19751 38267
rect 24838 38233 24872 38267
rect 28457 38233 28491 38267
rect 30674 38233 30708 38267
rect 31769 38233 31803 38267
rect 2605 38165 2639 38199
rect 7297 38165 7331 38199
rect 10609 38165 10643 38199
rect 17325 38165 17359 38199
rect 19993 38165 20027 38199
rect 25973 38165 26007 38199
rect 29561 38165 29595 38199
rect 31401 38165 31435 38199
rect 32321 38165 32355 38199
rect 3065 37961 3099 37995
rect 8309 37961 8343 37995
rect 10241 37961 10275 37995
rect 24409 37961 24443 37995
rect 25881 37961 25915 37995
rect 3433 37893 3467 37927
rect 10425 37893 10459 37927
rect 10609 37893 10643 37927
rect 11713 37893 11747 37927
rect 11805 37893 11839 37927
rect 17601 37893 17635 37927
rect 17693 37893 17727 37927
rect 25697 37893 25731 37927
rect 3249 37825 3283 37859
rect 8493 37825 8527 37859
rect 11529 37825 11563 37859
rect 11897 37825 11931 37859
rect 17325 37825 17359 37859
rect 17418 37825 17452 37859
rect 17831 37825 17865 37859
rect 18429 37825 18463 37859
rect 18685 37825 18719 37859
rect 20269 37825 20303 37859
rect 20453 37825 20487 37859
rect 24685 37825 24719 37859
rect 24777 37825 24811 37859
rect 24869 37825 24903 37859
rect 25053 37825 25087 37859
rect 25513 37825 25547 37859
rect 27813 37825 27847 37859
rect 30297 37825 30331 37859
rect 30481 37825 30515 37859
rect 30573 37825 30607 37859
rect 30665 37825 30699 37859
rect 31401 37825 31435 37859
rect 32588 37825 32622 37859
rect 32321 37757 32355 37791
rect 12081 37689 12115 37723
rect 3985 37621 4019 37655
rect 9137 37621 9171 37655
rect 17969 37621 18003 37655
rect 19809 37621 19843 37655
rect 20637 37621 20671 37655
rect 23305 37621 23339 37655
rect 23949 37621 23983 37655
rect 29101 37621 29135 37655
rect 30941 37621 30975 37655
rect 33701 37621 33735 37655
rect 34621 37621 34655 37655
rect 58173 37621 58207 37655
rect 16773 37417 16807 37451
rect 18245 37417 18279 37451
rect 20453 37417 20487 37451
rect 7021 37349 7055 37383
rect 24409 37349 24443 37383
rect 33701 37349 33735 37383
rect 1869 37213 1903 37247
rect 5641 37213 5675 37247
rect 7481 37213 7515 37247
rect 7757 37213 7791 37247
rect 7849 37213 7883 37247
rect 14105 37213 14139 37247
rect 15393 37213 15427 37247
rect 17607 37213 17641 37247
rect 17785 37213 17819 37247
rect 17877 37213 17911 37247
rect 17989 37213 18023 37247
rect 19349 37213 19383 37247
rect 19442 37213 19476 37247
rect 19717 37213 19751 37247
rect 19855 37213 19889 37247
rect 21833 37213 21867 37247
rect 23029 37213 23063 37247
rect 23121 37213 23155 37247
rect 23397 37213 23431 37247
rect 24961 37213 24995 37247
rect 30573 37213 30607 37247
rect 32413 37213 32447 37247
rect 34713 37213 34747 37247
rect 34897 37213 34931 37247
rect 34989 37213 35023 37247
rect 35081 37213 35115 37247
rect 2136 37145 2170 37179
rect 5908 37145 5942 37179
rect 7665 37145 7699 37179
rect 14289 37145 14323 37179
rect 15638 37145 15672 37179
rect 19625 37145 19659 37179
rect 21566 37145 21600 37179
rect 23213 37145 23247 37179
rect 25206 37145 25240 37179
rect 30840 37145 30874 37179
rect 3249 37077 3283 37111
rect 8033 37077 8067 37111
rect 14473 37077 14507 37111
rect 19993 37077 20027 37111
rect 22293 37077 22327 37111
rect 22845 37077 22879 37111
rect 26341 37077 26375 37111
rect 28917 37077 28951 37111
rect 29653 37077 29687 37111
rect 31953 37077 31987 37111
rect 35357 37077 35391 37111
rect 14565 36873 14599 36907
rect 15485 36873 15519 36907
rect 18153 36873 18187 36907
rect 18705 36873 18739 36907
rect 20453 36873 20487 36907
rect 24961 36873 24995 36907
rect 29929 36873 29963 36907
rect 32597 36873 32631 36907
rect 36277 36873 36311 36907
rect 3157 36805 3191 36839
rect 6837 36805 6871 36839
rect 7757 36805 7791 36839
rect 16865 36805 16899 36839
rect 17969 36805 18003 36839
rect 23673 36805 23707 36839
rect 25973 36805 26007 36839
rect 34437 36805 34471 36839
rect 35142 36805 35176 36839
rect 4905 36737 4939 36771
rect 6561 36737 6595 36771
rect 6745 36737 6779 36771
rect 6929 36737 6963 36771
rect 7941 36737 7975 36771
rect 12081 36737 12115 36771
rect 13185 36737 13219 36771
rect 13452 36737 13486 36771
rect 15741 36737 15775 36771
rect 15853 36737 15887 36771
rect 15945 36740 15979 36774
rect 16129 36737 16163 36771
rect 17049 36737 17083 36771
rect 17785 36737 17819 36771
rect 19809 36737 19843 36771
rect 19993 36737 20027 36771
rect 20085 36737 20119 36771
rect 20177 36737 20211 36771
rect 20913 36737 20947 36771
rect 22845 36737 22879 36771
rect 22937 36737 22971 36771
rect 23029 36737 23063 36771
rect 23213 36737 23247 36771
rect 27445 36737 27479 36771
rect 27701 36737 27735 36771
rect 29285 36737 29319 36771
rect 29469 36737 29503 36771
rect 29561 36737 29595 36771
rect 29653 36737 29687 36771
rect 31125 36737 31159 36771
rect 32873 36737 32907 36771
rect 32965 36737 32999 36771
rect 33057 36737 33091 36771
rect 33241 36737 33275 36771
rect 33793 36737 33827 36771
rect 33977 36737 34011 36771
rect 34069 36737 34103 36771
rect 34161 36737 34195 36771
rect 34897 36737 34931 36771
rect 31401 36669 31435 36703
rect 5457 36601 5491 36635
rect 16681 36601 16715 36635
rect 7113 36533 7147 36567
rect 7573 36533 7607 36567
rect 12173 36533 12207 36567
rect 19349 36533 19383 36567
rect 22201 36533 22235 36567
rect 22661 36533 22695 36567
rect 28825 36533 28859 36567
rect 5181 36329 5215 36363
rect 7021 36329 7055 36363
rect 9689 36329 9723 36363
rect 12541 36329 12575 36363
rect 14105 36329 14139 36363
rect 15209 36329 15243 36363
rect 16313 36329 16347 36363
rect 27077 36329 27111 36363
rect 27537 36329 27571 36363
rect 29561 36329 29595 36363
rect 34161 36329 34195 36363
rect 35081 36329 35115 36363
rect 25145 36261 25179 36295
rect 3801 36193 3835 36227
rect 26525 36193 26559 36227
rect 28641 36193 28675 36227
rect 35633 36193 35667 36227
rect 7297 36125 7331 36159
rect 7386 36119 7420 36153
rect 7481 36125 7515 36159
rect 7665 36125 7699 36159
rect 9505 36125 9539 36159
rect 10149 36125 10183 36159
rect 14381 36125 14415 36159
rect 14473 36125 14507 36159
rect 14565 36125 14599 36159
rect 14749 36125 14783 36159
rect 22293 36125 22327 36159
rect 22661 36125 22695 36159
rect 23489 36125 23523 36159
rect 23673 36125 23707 36159
rect 27813 36125 27847 36159
rect 27905 36125 27939 36159
rect 27997 36125 28031 36159
rect 28181 36125 28215 36159
rect 29009 36125 29043 36159
rect 31953 36125 31987 36159
rect 32229 36125 32263 36159
rect 34713 36125 34747 36159
rect 35889 36125 35923 36159
rect 58173 36125 58207 36159
rect 4068 36057 4102 36091
rect 10416 36057 10450 36091
rect 12633 36057 12667 36091
rect 13369 36057 13403 36091
rect 22385 36057 22419 36091
rect 22477 36057 22511 36091
rect 23857 36057 23891 36091
rect 26258 36057 26292 36091
rect 28825 36057 28859 36091
rect 29745 36057 29779 36091
rect 29929 36057 29963 36091
rect 33793 36057 33827 36091
rect 33977 36057 34011 36091
rect 34897 36057 34931 36091
rect 6561 35989 6595 36023
rect 11529 35989 11563 36023
rect 13461 35989 13495 36023
rect 22109 35989 22143 36023
rect 24409 35989 24443 36023
rect 30389 35989 30423 36023
rect 31401 35989 31435 36023
rect 33333 35989 33367 36023
rect 37013 35989 37047 36023
rect 12725 35785 12759 35819
rect 25145 35785 25179 35819
rect 33333 35785 33367 35819
rect 4537 35717 4571 35751
rect 11529 35717 11563 35751
rect 13185 35717 13219 35751
rect 23489 35717 23523 35751
rect 33517 35717 33551 35751
rect 4353 35649 4387 35683
rect 7490 35649 7524 35683
rect 7757 35649 7791 35683
rect 11713 35649 11747 35683
rect 13369 35649 13403 35683
rect 17417 35649 17451 35683
rect 17601 35649 17635 35683
rect 23673 35649 23707 35683
rect 24501 35649 24535 35683
rect 24685 35649 24719 35683
rect 24796 35655 24830 35689
rect 24915 35649 24949 35683
rect 25605 35649 25639 35683
rect 32229 35649 32263 35683
rect 33701 35649 33735 35683
rect 9045 35581 9079 35615
rect 9321 35581 9355 35615
rect 9781 35581 9815 35615
rect 10057 35581 10091 35615
rect 23857 35581 23891 35615
rect 27169 35513 27203 35547
rect 34161 35513 34195 35547
rect 4721 35445 4755 35479
rect 5273 35445 5307 35479
rect 6377 35445 6411 35479
rect 11897 35445 11931 35479
rect 13921 35445 13955 35479
rect 17785 35445 17819 35479
rect 22385 35445 22419 35479
rect 23029 35445 23063 35479
rect 32413 35445 32447 35479
rect 4261 35241 4295 35275
rect 7205 35241 7239 35275
rect 8401 35241 8435 35275
rect 11989 35241 12023 35275
rect 19441 35241 19475 35275
rect 25053 35241 25087 35275
rect 6745 35173 6779 35207
rect 9873 35105 9907 35139
rect 10609 35105 10643 35139
rect 17141 35105 17175 35139
rect 21649 35105 21683 35139
rect 4537 35037 4571 35071
rect 4629 35037 4663 35071
rect 4721 35037 4755 35071
rect 4905 35037 4939 35071
rect 7461 35037 7495 35071
rect 7573 35037 7607 35071
rect 7665 35037 7699 35071
rect 7849 35037 7883 35071
rect 10149 35037 10183 35071
rect 13021 35037 13055 35071
rect 13369 35037 13403 35071
rect 22109 35037 22143 35071
rect 24409 35037 24443 35071
rect 24593 35037 24627 35071
rect 24685 35037 24719 35071
rect 24823 35037 24857 35071
rect 31493 35037 31527 35071
rect 31769 35037 31803 35071
rect 58173 35037 58207 35071
rect 6377 34969 6411 35003
rect 6561 34969 6595 35003
rect 10876 34969 10910 35003
rect 13185 34969 13219 35003
rect 13277 34969 13311 35003
rect 17386 34969 17420 35003
rect 21382 34969 21416 35003
rect 30297 34969 30331 35003
rect 30481 34969 30515 35003
rect 5457 34901 5491 34935
rect 13553 34901 13587 34935
rect 18521 34901 18555 34935
rect 20269 34901 20303 34935
rect 23857 34901 23891 34935
rect 25513 34901 25547 34935
rect 30113 34901 30147 34935
rect 33701 34901 33735 34935
rect 3985 34697 4019 34731
rect 9045 34697 9079 34731
rect 10333 34697 10367 34731
rect 12449 34697 12483 34731
rect 13645 34697 13679 34731
rect 17141 34697 17175 34731
rect 20269 34697 20303 34731
rect 20821 34697 20855 34731
rect 31585 34697 31619 34731
rect 2872 34629 2906 34663
rect 4445 34629 4479 34663
rect 8769 34629 8803 34663
rect 9505 34629 9539 34663
rect 11897 34629 11931 34663
rect 13369 34629 13403 34663
rect 18981 34629 19015 34663
rect 27905 34629 27939 34663
rect 29101 34629 29135 34663
rect 30450 34629 30484 34663
rect 2605 34561 2639 34595
rect 4721 34561 4755 34595
rect 4810 34561 4844 34595
rect 4905 34561 4939 34595
rect 5089 34561 5123 34595
rect 7849 34561 7883 34595
rect 8401 34561 8435 34595
rect 8494 34561 8528 34595
rect 8677 34561 8711 34595
rect 8907 34561 8941 34595
rect 9689 34561 9723 34595
rect 10589 34561 10623 34595
rect 10682 34561 10716 34595
rect 10793 34561 10827 34595
rect 10977 34561 11011 34595
rect 11529 34561 11563 34595
rect 11713 34561 11747 34595
rect 13093 34561 13127 34595
rect 13277 34561 13311 34595
rect 13461 34561 13495 34595
rect 17417 34561 17451 34595
rect 17509 34561 17543 34595
rect 17601 34561 17635 34595
rect 17785 34561 17819 34595
rect 18797 34561 18831 34595
rect 19625 34561 19659 34595
rect 19809 34561 19843 34595
rect 19901 34561 19935 34595
rect 19993 34561 20027 34595
rect 22201 34561 22235 34595
rect 22364 34561 22398 34595
rect 22480 34564 22514 34598
rect 22569 34561 22603 34595
rect 28089 34561 28123 34595
rect 29377 34561 29411 34595
rect 29469 34561 29503 34595
rect 29561 34561 29595 34595
rect 29745 34561 29779 34595
rect 33793 34561 33827 34595
rect 33977 34561 34011 34595
rect 34072 34564 34106 34598
rect 34161 34561 34195 34595
rect 19165 34493 19199 34527
rect 28549 34493 28583 34527
rect 30205 34493 30239 34527
rect 34437 34493 34471 34527
rect 16037 34425 16071 34459
rect 5549 34357 5583 34391
rect 22845 34357 22879 34391
rect 24777 34357 24811 34391
rect 27721 34357 27755 34391
rect 33333 34357 33367 34391
rect 5733 34153 5767 34187
rect 11069 34153 11103 34187
rect 14565 34153 14599 34187
rect 18521 34153 18555 34187
rect 21833 34153 21867 34187
rect 25881 34153 25915 34187
rect 35081 34153 35115 34187
rect 13553 34085 13587 34119
rect 22293 34017 22327 34051
rect 30205 34017 30239 34051
rect 33057 34017 33091 34051
rect 4077 33949 4111 33983
rect 4169 33949 4203 33983
rect 4261 33949 4295 33983
rect 4445 33949 4479 33983
rect 10425 33949 10459 33983
rect 10588 33949 10622 33983
rect 10701 33949 10735 33983
rect 10839 33949 10873 33983
rect 11529 33949 11563 33983
rect 13369 33949 13403 33983
rect 16865 33949 16899 33983
rect 17601 33949 17635 33983
rect 17693 33949 17727 33983
rect 17785 33949 17819 33983
rect 17969 33949 18003 33983
rect 19349 33949 19383 33983
rect 19442 33949 19476 33983
rect 19814 33949 19848 33983
rect 22560 33949 22594 33983
rect 24869 33949 24903 33983
rect 26985 33949 27019 33983
rect 29009 33949 29043 33983
rect 29929 33949 29963 33983
rect 32689 33949 32723 33983
rect 33517 33949 33551 33983
rect 33701 33949 33735 33983
rect 33793 33949 33827 33983
rect 33885 33949 33919 33983
rect 34897 33949 34931 33983
rect 4905 33881 4939 33915
rect 5089 33881 5123 33915
rect 5273 33881 5307 33915
rect 14657 33881 14691 33915
rect 16609 33881 16643 33915
rect 17325 33881 17359 33915
rect 19625 33881 19659 33915
rect 19717 33881 19751 33915
rect 21465 33881 21499 33915
rect 21649 33881 21683 33915
rect 25053 33881 25087 33915
rect 27252 33881 27286 33915
rect 31217 33881 31251 33915
rect 31401 33881 31435 33915
rect 32873 33881 32907 33915
rect 34713 33881 34747 33915
rect 3801 33813 3835 33847
rect 7573 33813 7607 33847
rect 15485 33813 15519 33847
rect 19993 33813 20027 33847
rect 23673 33813 23707 33847
rect 25237 33813 25271 33847
rect 28365 33813 28399 33847
rect 31585 33813 31619 33847
rect 34161 33813 34195 33847
rect 4445 33609 4479 33643
rect 5273 33609 5307 33643
rect 8033 33609 8067 33643
rect 17049 33609 17083 33643
rect 27261 33609 27295 33643
rect 34529 33609 34563 33643
rect 2872 33541 2906 33575
rect 4629 33541 4663 33575
rect 14136 33541 14170 33575
rect 14841 33541 14875 33575
rect 16865 33541 16899 33575
rect 19165 33541 19199 33575
rect 22100 33541 22134 33575
rect 23949 33541 23983 33575
rect 31401 33541 31435 33575
rect 35642 33541 35676 33575
rect 2605 33473 2639 33507
rect 4813 33473 4847 33507
rect 6920 33473 6954 33507
rect 12449 33473 12483 33507
rect 15117 33473 15151 33507
rect 15209 33473 15243 33507
rect 15301 33473 15335 33507
rect 15485 33473 15519 33507
rect 16681 33473 16715 33507
rect 17877 33473 17911 33507
rect 18521 33473 18555 33507
rect 19349 33473 19383 33507
rect 21833 33473 21867 33507
rect 24225 33473 24259 33507
rect 24317 33473 24351 33507
rect 24409 33473 24443 33507
rect 24593 33473 24627 33507
rect 25053 33473 25087 33507
rect 25237 33473 25271 33507
rect 25329 33473 25363 33507
rect 25467 33473 25501 33507
rect 27537 33473 27571 33507
rect 27629 33473 27663 33507
rect 27721 33473 27755 33507
rect 27905 33473 27939 33507
rect 30389 33473 30423 33507
rect 30481 33473 30515 33507
rect 30573 33473 30607 33507
rect 30757 33473 30791 33507
rect 32689 33473 32723 33507
rect 32956 33473 32990 33507
rect 6653 33405 6687 33439
rect 14381 33405 14415 33439
rect 35909 33405 35943 33439
rect 12265 33337 12299 33371
rect 18337 33337 18371 33371
rect 25697 33337 25731 33371
rect 31217 33337 31251 33371
rect 58173 33337 58207 33371
rect 3985 33269 4019 33303
rect 11529 33269 11563 33303
rect 13001 33269 13035 33303
rect 19993 33269 20027 33303
rect 23213 33269 23247 33303
rect 26341 33269 26375 33303
rect 29561 33269 29595 33303
rect 30113 33269 30147 33303
rect 34069 33269 34103 33303
rect 5549 33065 5583 33099
rect 6745 33065 6779 33099
rect 13553 33065 13587 33099
rect 23857 33065 23891 33099
rect 27721 33065 27755 33099
rect 7849 32929 7883 32963
rect 9689 32929 9723 32963
rect 14381 32929 14415 32963
rect 24409 32929 24443 32963
rect 24685 32929 24719 32963
rect 32321 32929 32355 32963
rect 32597 32929 32631 32963
rect 7021 32861 7055 32895
rect 7113 32861 7147 32895
rect 7205 32861 7239 32895
rect 7389 32861 7423 32895
rect 8033 32861 8067 32895
rect 10333 32861 10367 32895
rect 13185 32861 13219 32895
rect 14105 32861 14139 32895
rect 16221 32861 16255 32895
rect 16314 32861 16348 32895
rect 16727 32861 16761 32895
rect 17693 32861 17727 32895
rect 18245 32861 18279 32895
rect 23489 32861 23523 32895
rect 26902 32861 26936 32895
rect 27169 32861 27203 32895
rect 30297 32861 30331 32895
rect 31493 32861 31527 32895
rect 35826 32861 35860 32895
rect 36093 32861 36127 32895
rect 8217 32793 8251 32827
rect 9505 32793 9539 32827
rect 10149 32793 10183 32827
rect 13369 32793 13403 32827
rect 16497 32793 16531 32827
rect 16589 32793 16623 32827
rect 18429 32793 18463 32827
rect 18613 32793 18647 32827
rect 23673 32793 23707 32827
rect 31677 32793 31711 32827
rect 6193 32725 6227 32759
rect 10517 32725 10551 32759
rect 11069 32725 11103 32759
rect 15485 32725 15519 32759
rect 16865 32725 16899 32759
rect 22109 32725 22143 32759
rect 25789 32725 25823 32759
rect 29745 32725 29779 32759
rect 30481 32725 30515 32759
rect 31861 32725 31895 32759
rect 34713 32725 34747 32759
rect 5181 32521 5215 32555
rect 5641 32521 5675 32555
rect 14013 32521 14047 32555
rect 20085 32521 20119 32555
rect 25329 32521 25363 32555
rect 30573 32521 30607 32555
rect 32873 32521 32907 32555
rect 6653 32453 6687 32487
rect 18245 32453 18279 32487
rect 18950 32453 18984 32487
rect 28457 32453 28491 32487
rect 2493 32385 2527 32419
rect 5825 32385 5859 32419
rect 6837 32385 6871 32419
rect 9597 32385 9631 32419
rect 10609 32385 10643 32419
rect 10701 32385 10735 32419
rect 10793 32385 10827 32419
rect 10977 32385 11011 32419
rect 11621 32385 11655 32419
rect 17601 32385 17635 32419
rect 17785 32385 17819 32419
rect 17877 32385 17911 32419
rect 17969 32385 18003 32419
rect 22201 32385 22235 32419
rect 24317 32385 24351 32419
rect 28365 32385 28399 32419
rect 28549 32385 28583 32419
rect 28733 32385 28767 32419
rect 30389 32385 30423 32419
rect 32229 32385 32263 32419
rect 32413 32385 32447 32419
rect 32505 32385 32539 32419
rect 32597 32385 32631 32419
rect 38402 32385 38436 32419
rect 2237 32317 2271 32351
rect 8309 32317 8343 32351
rect 8585 32317 8619 32351
rect 9873 32317 9907 32351
rect 18705 32317 18739 32351
rect 38669 32317 38703 32351
rect 24501 32249 24535 32283
rect 3617 32181 3651 32215
rect 7021 32181 7055 32215
rect 10333 32181 10367 32215
rect 22385 32181 22419 32215
rect 28181 32181 28215 32215
rect 37289 32181 37323 32215
rect 58173 32181 58207 32215
rect 2145 31977 2179 32011
rect 7205 31977 7239 32011
rect 10885 31977 10919 32011
rect 13369 31977 13403 32011
rect 30941 31977 30975 32011
rect 32137 31977 32171 32011
rect 36645 31977 36679 32011
rect 8125 31909 8159 31943
rect 28089 31909 28123 31943
rect 35449 31909 35483 31943
rect 9505 31841 9539 31875
rect 16313 31841 16347 31875
rect 22845 31841 22879 31875
rect 25053 31841 25087 31875
rect 29561 31841 29595 31875
rect 2375 31773 2409 31807
rect 2494 31770 2528 31804
rect 2605 31773 2639 31807
rect 2789 31773 2823 31807
rect 5089 31773 5123 31807
rect 5181 31773 5215 31807
rect 5273 31773 5307 31807
rect 5457 31773 5491 31807
rect 5917 31773 5951 31807
rect 9772 31773 9806 31807
rect 13001 31773 13035 31807
rect 14361 31773 14395 31807
rect 14470 31773 14504 31807
rect 14565 31770 14599 31804
rect 14749 31773 14783 31807
rect 16773 31773 16807 31807
rect 21465 31773 21499 31807
rect 22569 31773 22603 31807
rect 24777 31773 24811 31807
rect 28273 31773 28307 31807
rect 28365 31773 28399 31807
rect 28641 31773 28675 31807
rect 29828 31773 29862 31807
rect 36001 31773 36035 31807
rect 36185 31773 36219 31807
rect 36280 31767 36314 31801
rect 36389 31773 36423 31807
rect 13185 31705 13219 31739
rect 16129 31705 16163 31739
rect 28457 31705 28491 31739
rect 4813 31637 4847 31671
rect 14105 31637 14139 31671
rect 15301 31637 15335 31671
rect 18061 31637 18095 31671
rect 26065 31637 26099 31671
rect 32597 31637 32631 31671
rect 37565 31637 37599 31671
rect 2421 31433 2455 31467
rect 5457 31433 5491 31467
rect 8309 31433 8343 31467
rect 12265 31433 12299 31467
rect 16773 31433 16807 31467
rect 25237 31433 25271 31467
rect 26065 31433 26099 31467
rect 32137 31433 32171 31467
rect 36185 31433 36219 31467
rect 5825 31365 5859 31399
rect 13400 31365 13434 31399
rect 15209 31365 15243 31399
rect 15301 31365 15335 31399
rect 31125 31365 31159 31399
rect 32965 31365 32999 31399
rect 2605 31297 2639 31331
rect 2789 31297 2823 31331
rect 5641 31297 5675 31331
rect 6653 31297 6687 31331
rect 6742 31300 6776 31334
rect 6842 31297 6876 31331
rect 7021 31297 7055 31331
rect 9597 31297 9631 31331
rect 14933 31297 14967 31331
rect 15026 31297 15060 31331
rect 15398 31297 15432 31331
rect 17785 31297 17819 31331
rect 19708 31297 19742 31331
rect 22477 31297 22511 31331
rect 22661 31297 22695 31331
rect 23949 31297 23983 31331
rect 25421 31297 25455 31331
rect 25881 31297 25915 31331
rect 30389 31297 30423 31331
rect 31033 31297 31067 31331
rect 31217 31297 31251 31331
rect 31401 31297 31435 31331
rect 32321 31297 32355 31331
rect 32413 31297 32447 31331
rect 33149 31297 33183 31331
rect 35817 31297 35851 31331
rect 36001 31297 36035 31331
rect 37657 31297 37691 31331
rect 13645 31229 13679 31263
rect 17509 31229 17543 31263
rect 19441 31229 19475 31263
rect 23305 31229 23339 31263
rect 24685 31229 24719 31263
rect 3341 31093 3375 31127
rect 6377 31093 6411 31127
rect 10149 31093 10183 31127
rect 15577 31093 15611 31127
rect 20821 31093 20855 31127
rect 22845 31093 22879 31127
rect 24041 31093 24075 31127
rect 28089 31093 28123 31127
rect 29101 31093 29135 31127
rect 30849 31093 30883 31127
rect 33333 31093 33367 31127
rect 38945 31093 38979 31127
rect 8217 30889 8251 30923
rect 13369 30889 13403 30923
rect 15117 30889 15151 30923
rect 21741 30889 21775 30923
rect 39313 30889 39347 30923
rect 18705 30821 18739 30855
rect 28549 30821 28583 30855
rect 33241 30821 33275 30855
rect 1869 30753 1903 30787
rect 26801 30753 26835 30787
rect 30389 30753 30423 30787
rect 4537 30685 4571 30719
rect 6377 30685 6411 30719
rect 12817 30685 12851 30719
rect 13093 30685 13127 30719
rect 13185 30685 13219 30719
rect 14289 30685 14323 30719
rect 14473 30685 14507 30719
rect 16497 30685 16531 30719
rect 17325 30685 17359 30719
rect 22569 30685 22603 30719
rect 22661 30685 22695 30719
rect 22753 30685 22787 30719
rect 22937 30685 22971 30719
rect 24501 30685 24535 30719
rect 30113 30685 30147 30719
rect 31493 30685 31527 30719
rect 32045 30685 32079 30719
rect 32229 30685 32263 30719
rect 32321 30685 32355 30719
rect 32413 30685 32447 30719
rect 33425 30685 33459 30719
rect 33517 30685 33551 30719
rect 33793 30685 33827 30719
rect 35357 30685 35391 30719
rect 36001 30685 36035 30719
rect 36185 30685 36219 30719
rect 36280 30685 36314 30719
rect 36369 30685 36403 30719
rect 37105 30685 37139 30719
rect 37933 30685 37967 30719
rect 58173 30685 58207 30719
rect 2136 30617 2170 30651
rect 4804 30617 4838 30651
rect 6644 30617 6678 30651
rect 13001 30617 13035 30651
rect 16230 30617 16264 30651
rect 17592 30617 17626 30651
rect 24685 30617 24719 30651
rect 26534 30617 26568 30651
rect 27261 30617 27295 30651
rect 33609 30617 33643 30651
rect 35173 30617 35207 30651
rect 35541 30617 35575 30651
rect 36645 30617 36679 30651
rect 38178 30617 38212 30651
rect 3249 30549 3283 30583
rect 5917 30549 5951 30583
rect 7757 30549 7791 30583
rect 9965 30549 9999 30583
rect 14657 30549 14691 30583
rect 19349 30549 19383 30583
rect 20269 30549 20303 30583
rect 22293 30549 22327 30583
rect 24869 30549 24903 30583
rect 25421 30549 25455 30583
rect 29653 30549 29687 30583
rect 32689 30549 32723 30583
rect 2145 30345 2179 30379
rect 7389 30345 7423 30379
rect 3617 30277 3651 30311
rect 7941 30277 7975 30311
rect 8125 30277 8159 30311
rect 10241 30277 10275 30311
rect 10609 30277 10643 30311
rect 11621 30277 11655 30311
rect 15669 30277 15703 30311
rect 18061 30277 18095 30311
rect 19809 30277 19843 30311
rect 24225 30277 24259 30311
rect 25789 30277 25823 30311
rect 29285 30277 29319 30311
rect 31033 30277 31067 30311
rect 31125 30277 31159 30311
rect 33710 30277 33744 30311
rect 35449 30277 35483 30311
rect 2401 30209 2435 30243
rect 2494 30209 2528 30243
rect 2605 30209 2639 30243
rect 2789 30209 2823 30243
rect 3433 30209 3467 30243
rect 9413 30209 9447 30243
rect 9505 30209 9539 30243
rect 9597 30209 9631 30243
rect 9781 30209 9815 30243
rect 10425 30209 10459 30243
rect 11805 30209 11839 30243
rect 15025 30209 15059 30243
rect 15209 30209 15243 30243
rect 15304 30209 15338 30243
rect 15393 30209 15427 30243
rect 16865 30209 16899 30243
rect 18337 30209 18371 30243
rect 18429 30209 18463 30243
rect 18521 30209 18555 30243
rect 18705 30209 18739 30243
rect 19165 30209 19199 30243
rect 19349 30209 19383 30243
rect 19441 30209 19475 30243
rect 19533 30209 19567 30243
rect 21005 30209 21039 30243
rect 22376 30209 22410 30243
rect 24133 30209 24167 30243
rect 24317 30209 24351 30243
rect 24501 30209 24535 30243
rect 25145 30209 25179 30243
rect 25329 30209 25363 30243
rect 25421 30209 25455 30243
rect 25513 30209 25547 30243
rect 29101 30209 29135 30243
rect 30941 30209 30975 30243
rect 31309 30209 31343 30243
rect 35081 30209 35115 30243
rect 35265 30209 35299 30243
rect 35909 30209 35943 30243
rect 36072 30209 36106 30243
rect 36185 30209 36219 30243
rect 36277 30209 36311 30243
rect 37289 30209 37323 30243
rect 3249 30141 3283 30175
rect 11989 30141 12023 30175
rect 17049 30141 17083 30175
rect 21281 30141 21315 30175
rect 22109 30141 22143 30175
rect 33977 30141 34011 30175
rect 23489 30073 23523 30107
rect 26341 30073 26375 30107
rect 9137 30005 9171 30039
rect 12541 30005 12575 30039
rect 16681 30005 16715 30039
rect 17509 30005 17543 30039
rect 23949 30005 23983 30039
rect 28917 30005 28951 30039
rect 30757 30005 30791 30039
rect 32597 30005 32631 30039
rect 36553 30005 36587 30039
rect 2881 29801 2915 29835
rect 10977 29801 11011 29835
rect 11897 29801 11931 29835
rect 19257 29801 19291 29835
rect 20177 29801 20211 29835
rect 27813 29801 27847 29835
rect 29561 29801 29595 29835
rect 39313 29801 39347 29835
rect 15853 29733 15887 29767
rect 21281 29733 21315 29767
rect 9137 29665 9171 29699
rect 11345 29665 11379 29699
rect 37940 29665 37974 29699
rect 4353 29597 4387 29631
rect 4629 29597 4663 29631
rect 4721 29597 4755 29631
rect 9393 29597 9427 29631
rect 11161 29597 11195 29631
rect 18061 29597 18095 29631
rect 19441 29597 19475 29631
rect 20361 29597 20395 29631
rect 22569 29597 22603 29631
rect 22661 29597 22695 29631
rect 22937 29597 22971 29631
rect 23857 29597 23891 29631
rect 24869 29597 24903 29631
rect 25053 29597 25087 29631
rect 25145 29597 25179 29631
rect 25237 29597 25271 29631
rect 27353 29597 27387 29631
rect 28641 29597 28675 29631
rect 28733 29597 28767 29631
rect 28825 29597 28859 29631
rect 29009 29597 29043 29631
rect 30941 29597 30975 29631
rect 33701 29597 33735 29631
rect 33793 29597 33827 29631
rect 34069 29597 34103 29631
rect 38189 29597 38223 29631
rect 58173 29597 58207 29631
rect 4537 29529 4571 29563
rect 18245 29529 18279 29563
rect 19625 29529 19659 29563
rect 20545 29529 20579 29563
rect 21097 29529 21131 29563
rect 22753 29529 22787 29563
rect 25513 29529 25547 29563
rect 27086 29529 27120 29563
rect 28365 29529 28399 29563
rect 30674 29529 30708 29563
rect 33885 29529 33919 29563
rect 35817 29529 35851 29563
rect 36001 29529 36035 29563
rect 4905 29461 4939 29495
rect 10517 29461 10551 29495
rect 16865 29461 16899 29495
rect 17417 29461 17451 29495
rect 21741 29461 21775 29495
rect 22385 29461 22419 29495
rect 23673 29461 23707 29495
rect 25973 29461 26007 29495
rect 31953 29461 31987 29495
rect 33517 29461 33551 29495
rect 36185 29461 36219 29495
rect 3709 29257 3743 29291
rect 12817 29257 12851 29291
rect 15669 29257 15703 29291
rect 23857 29257 23891 29291
rect 24685 29257 24719 29291
rect 25237 29257 25271 29291
rect 25973 29257 26007 29291
rect 30573 29257 30607 29291
rect 36461 29257 36495 29291
rect 39313 29257 39347 29291
rect 4537 29189 4571 29223
rect 7941 29189 7975 29223
rect 10793 29189 10827 29223
rect 10977 29189 11011 29223
rect 13737 29189 13771 29223
rect 14841 29189 14875 29223
rect 17877 29189 17911 29223
rect 18797 29189 18831 29223
rect 20085 29189 20119 29223
rect 22109 29189 22143 29223
rect 22201 29189 22235 29223
rect 24501 29189 24535 29223
rect 29469 29189 29503 29223
rect 33793 29189 33827 29223
rect 33885 29189 33919 29223
rect 2789 29121 2823 29155
rect 2881 29121 2915 29155
rect 2973 29121 3007 29155
rect 3157 29121 3191 29155
rect 4261 29121 4295 29155
rect 4445 29121 4479 29155
rect 4629 29121 4663 29155
rect 7665 29121 7699 29155
rect 7849 29121 7883 29155
rect 9781 29121 9815 29155
rect 9870 29124 9904 29158
rect 9965 29121 9999 29155
rect 10149 29121 10183 29155
rect 13369 29121 13403 29155
rect 13462 29121 13496 29155
rect 13645 29121 13679 29155
rect 13834 29121 13868 29155
rect 14657 29121 14691 29155
rect 19901 29121 19935 29155
rect 20173 29121 20207 29155
rect 20269 29121 20303 29155
rect 22017 29121 22051 29155
rect 22385 29121 22419 29155
rect 22937 29121 22971 29155
rect 24317 29121 24351 29155
rect 25421 29121 25455 29155
rect 26157 29121 26191 29155
rect 26985 29121 27019 29155
rect 29377 29121 29411 29155
rect 29561 29121 29595 29155
rect 29745 29121 29779 29155
rect 30389 29121 30423 29155
rect 30573 29121 30607 29155
rect 31033 29121 31067 29155
rect 33701 29121 33735 29155
rect 34069 29121 34103 29155
rect 34529 29121 34563 29155
rect 38189 29121 38223 29155
rect 9045 29053 9079 29087
rect 10609 29053 10643 29087
rect 35173 29053 35207 29087
rect 35449 29053 35483 29087
rect 37933 29053 37967 29087
rect 4813 28985 4847 29019
rect 11529 28985 11563 29019
rect 14013 28985 14047 29019
rect 19349 28985 19383 29019
rect 20453 28985 20487 29019
rect 23121 28985 23155 29019
rect 29193 28985 29227 29019
rect 33517 28985 33551 29019
rect 34713 28985 34747 29019
rect 2513 28917 2547 28951
rect 8401 28917 8435 28951
rect 9505 28917 9539 28951
rect 15025 28917 15059 28951
rect 20913 28917 20947 28951
rect 21833 28917 21867 28951
rect 2973 28713 3007 28747
rect 26893 28713 26927 28747
rect 29653 28713 29687 28747
rect 36645 28713 36679 28747
rect 16037 28645 16071 28679
rect 24593 28645 24627 28679
rect 12449 28577 12483 28611
rect 30757 28577 30791 28611
rect 33517 28577 33551 28611
rect 2605 28509 2639 28543
rect 4629 28509 4663 28543
rect 4905 28509 4939 28543
rect 4997 28509 5031 28543
rect 9229 28509 9263 28543
rect 9496 28509 9530 28543
rect 12081 28509 12115 28543
rect 13185 28509 13219 28543
rect 13277 28509 13311 28543
rect 13369 28509 13403 28543
rect 13553 28509 13587 28543
rect 14657 28509 14691 28543
rect 14841 28509 14875 28543
rect 14933 28509 14967 28543
rect 15025 28509 15059 28543
rect 15853 28509 15887 28543
rect 24409 28509 24443 28543
rect 26249 28509 26283 28543
rect 26709 28509 26743 28543
rect 29561 28509 29595 28543
rect 29745 28509 29779 28543
rect 31033 28509 31067 28543
rect 33793 28509 33827 28543
rect 34897 28509 34931 28543
rect 34989 28509 35023 28543
rect 35265 28509 35299 28543
rect 36001 28509 36035 28543
rect 36185 28506 36219 28540
rect 36280 28509 36314 28543
rect 36415 28509 36449 28543
rect 37105 28509 37139 28543
rect 2789 28441 2823 28475
rect 4813 28441 4847 28475
rect 12265 28441 12299 28475
rect 14197 28441 14231 28475
rect 17509 28441 17543 28475
rect 18061 28441 18095 28475
rect 23489 28441 23523 28475
rect 25237 28441 25271 28475
rect 35081 28441 35115 28475
rect 37289 28441 37323 28475
rect 5181 28373 5215 28407
rect 10609 28373 10643 28407
rect 12909 28373 12943 28407
rect 15301 28373 15335 28407
rect 16957 28373 16991 28407
rect 18153 28373 18187 28407
rect 29009 28373 29043 28407
rect 31493 28373 31527 28407
rect 34713 28373 34747 28407
rect 37473 28373 37507 28407
rect 3801 28169 3835 28203
rect 8585 28169 8619 28203
rect 9413 28169 9447 28203
rect 11529 28169 11563 28203
rect 13093 28169 13127 28203
rect 13921 28169 13955 28203
rect 14381 28169 14415 28203
rect 30297 28169 30331 28203
rect 35541 28169 35575 28203
rect 2666 28101 2700 28135
rect 5365 28101 5399 28135
rect 6745 28101 6779 28135
rect 12725 28101 12759 28135
rect 15494 28101 15528 28135
rect 22293 28101 22327 28135
rect 34529 28101 34563 28135
rect 36737 28101 36771 28135
rect 38494 28101 38528 28135
rect 4997 28033 5031 28067
rect 5090 28033 5124 28067
rect 5273 28033 5307 28067
rect 5503 28033 5537 28067
rect 6377 28033 6411 28067
rect 6525 28033 6559 28067
rect 6653 28033 6687 28067
rect 6881 28033 6915 28067
rect 8401 28033 8435 28067
rect 8585 28033 8619 28067
rect 9229 28033 9263 28067
rect 9413 28033 9447 28067
rect 11713 28033 11747 28067
rect 11805 28033 11839 28067
rect 12541 28033 12575 28067
rect 12817 28033 12851 28067
rect 12909 28033 12943 28067
rect 15761 28033 15795 28067
rect 17141 28033 17175 28067
rect 18521 28033 18555 28067
rect 30113 28033 30147 28067
rect 31309 28033 31343 28067
rect 31585 28033 31619 28067
rect 32137 28033 32171 28067
rect 33701 28033 33735 28067
rect 34345 28033 34379 28067
rect 34437 28033 34471 28067
rect 34713 28033 34747 28067
rect 36093 28033 36127 28067
rect 36277 28033 36311 28067
rect 36369 28033 36403 28067
rect 36507 28033 36541 28067
rect 38761 28033 38795 28067
rect 2421 27965 2455 27999
rect 7941 27965 7975 27999
rect 18245 27965 18279 27999
rect 19533 27965 19567 27999
rect 19809 27965 19843 27999
rect 29929 27965 29963 27999
rect 33425 27965 33459 27999
rect 37381 27897 37415 27931
rect 58173 27897 58207 27931
rect 5641 27829 5675 27863
rect 7021 27829 7055 27863
rect 9873 27829 9907 27863
rect 17233 27829 17267 27863
rect 22385 27829 22419 27863
rect 24317 27829 24351 27863
rect 29377 27829 29411 27863
rect 34161 27829 34195 27863
rect 11713 27625 11747 27659
rect 13553 27625 13587 27659
rect 5549 27557 5583 27591
rect 17141 27557 17175 27591
rect 21097 27557 21131 27591
rect 30665 27489 30699 27523
rect 4905 27421 4939 27455
rect 4998 27421 5032 27455
rect 5181 27421 5215 27455
rect 5273 27421 5307 27455
rect 5411 27421 5445 27455
rect 6653 27421 6687 27455
rect 6746 27421 6780 27455
rect 7021 27421 7055 27455
rect 7118 27421 7152 27455
rect 7941 27421 7975 27455
rect 9229 27421 9263 27455
rect 9413 27421 9447 27455
rect 10885 27421 10919 27455
rect 11161 27421 11195 27455
rect 12173 27421 12207 27455
rect 12440 27421 12474 27455
rect 16489 27421 16523 27455
rect 16681 27421 16715 27455
rect 20453 27421 20487 27455
rect 20913 27421 20947 27455
rect 26433 27421 26467 27455
rect 30389 27421 30423 27455
rect 33149 27421 33183 27455
rect 6929 27353 6963 27387
rect 7757 27353 7791 27387
rect 16589 27353 16623 27387
rect 21649 27353 21683 27387
rect 21833 27353 21867 27387
rect 26678 27353 26712 27387
rect 32965 27353 32999 27387
rect 7297 27285 7331 27319
rect 8125 27285 8159 27319
rect 9321 27285 9355 27319
rect 17693 27285 17727 27319
rect 22017 27285 22051 27319
rect 24409 27285 24443 27319
rect 27813 27285 27847 27319
rect 29929 27285 29963 27319
rect 33333 27285 33367 27319
rect 6837 27081 6871 27115
rect 25421 27081 25455 27115
rect 3617 27013 3651 27047
rect 26065 27013 26099 27047
rect 32873 27013 32907 27047
rect 33885 27013 33919 27047
rect 34805 27013 34839 27047
rect 3433 26945 3467 26979
rect 7950 26945 7984 26979
rect 8217 26945 8251 26979
rect 10057 26945 10091 26979
rect 11897 26945 11931 26979
rect 13185 26945 13219 26979
rect 16957 26945 16991 26979
rect 17224 26945 17258 26979
rect 19165 26945 19199 26979
rect 19421 26945 19455 26979
rect 23498 26945 23532 26979
rect 23765 26945 23799 26979
rect 24777 26945 24811 26979
rect 24940 26951 24974 26985
rect 25056 26945 25090 26979
rect 25191 26945 25225 26979
rect 26249 26945 26283 26979
rect 27905 26945 27939 26979
rect 28161 26945 28195 26979
rect 31033 26945 31067 26979
rect 32781 26945 32815 26979
rect 32965 26945 32999 26979
rect 33149 26945 33183 26979
rect 33793 26945 33827 26979
rect 33977 26945 34011 26979
rect 34161 26945 34195 26979
rect 34621 26945 34655 26979
rect 39885 26945 39919 26979
rect 9781 26877 9815 26911
rect 11621 26877 11655 26911
rect 12909 26877 12943 26911
rect 30757 26877 30791 26911
rect 40141 26877 40175 26911
rect 8769 26809 8803 26843
rect 30205 26809 30239 26843
rect 3801 26741 3835 26775
rect 9229 26741 9263 26775
rect 18337 26741 18371 26775
rect 20545 26741 20579 26775
rect 22385 26741 22419 26775
rect 24225 26741 24259 26775
rect 25881 26741 25915 26775
rect 29285 26741 29319 26775
rect 32597 26741 32631 26775
rect 33609 26741 33643 26775
rect 34989 26741 35023 26775
rect 38761 26741 38795 26775
rect 58173 26741 58207 26775
rect 7205 26537 7239 26571
rect 7757 26537 7791 26571
rect 11897 26537 11931 26571
rect 12725 26537 12759 26571
rect 18705 26537 18739 26571
rect 27813 26537 27847 26571
rect 2881 26469 2915 26503
rect 11069 26401 11103 26435
rect 17141 26401 17175 26435
rect 25605 26401 25639 26435
rect 29009 26401 29043 26435
rect 29561 26401 29595 26435
rect 29837 26401 29871 26435
rect 3065 26333 3099 26367
rect 3249 26333 3283 26367
rect 4077 26333 4111 26367
rect 4169 26333 4203 26367
rect 4261 26333 4295 26367
rect 4445 26333 4479 26367
rect 8033 26333 8067 26367
rect 8125 26333 8159 26367
rect 8217 26333 8251 26367
rect 8401 26333 8435 26367
rect 11989 26333 12023 26367
rect 16313 26333 16347 26367
rect 16773 26333 16807 26367
rect 16957 26333 16991 26367
rect 18061 26333 18095 26367
rect 18224 26333 18258 26367
rect 18337 26333 18371 26367
rect 18475 26333 18509 26367
rect 21005 26333 21039 26367
rect 22753 26333 22787 26367
rect 23213 26333 23247 26367
rect 24501 26333 24535 26367
rect 24685 26333 24719 26367
rect 24777 26333 24811 26367
rect 24869 26333 24903 26367
rect 33471 26333 33505 26367
rect 33609 26333 33643 26367
rect 33701 26333 33735 26367
rect 33885 26333 33919 26367
rect 34713 26333 34747 26367
rect 34897 26333 34931 26367
rect 34989 26333 35023 26367
rect 35081 26333 35115 26367
rect 35817 26333 35851 26367
rect 40233 26333 40267 26367
rect 9321 26265 9355 26299
rect 12633 26265 12667 26299
rect 19349 26265 19383 26299
rect 25872 26265 25906 26299
rect 27445 26265 27479 26299
rect 27629 26265 27663 26299
rect 31033 26265 31067 26299
rect 32781 26265 32815 26299
rect 35357 26265 35391 26299
rect 40049 26265 40083 26299
rect 40877 26265 40911 26299
rect 41061 26265 41095 26299
rect 3801 26197 3835 26231
rect 4905 26197 4939 26231
rect 25145 26197 25179 26231
rect 26985 26197 27019 26231
rect 33241 26197 33275 26231
rect 40417 26197 40451 26231
rect 41245 26197 41279 26231
rect 3893 25993 3927 26027
rect 7481 25993 7515 26027
rect 8401 25993 8435 26027
rect 17509 25993 17543 26027
rect 18889 25993 18923 26027
rect 25145 25993 25179 26027
rect 26249 25993 26283 26027
rect 30849 25993 30883 26027
rect 32689 25993 32723 26027
rect 34989 25993 35023 26027
rect 40601 25993 40635 26027
rect 2780 25925 2814 25959
rect 5457 25925 5491 25959
rect 5641 25925 5675 25959
rect 8861 25925 8895 25959
rect 9045 25925 9079 25959
rect 14289 25925 14323 25959
rect 19073 25925 19107 25959
rect 20913 25925 20947 25959
rect 21281 25925 21315 25959
rect 26985 25925 27019 25959
rect 33394 25925 33428 25959
rect 36102 25925 36136 25959
rect 2513 25857 2547 25891
rect 6607 25857 6641 25891
rect 6726 25860 6760 25894
rect 6842 25857 6876 25891
rect 7021 25857 7055 25891
rect 9873 25857 9907 25891
rect 11713 25857 11747 25891
rect 13829 25857 13863 25891
rect 14473 25857 14507 25891
rect 15853 25857 15887 25891
rect 16865 25857 16899 25891
rect 17785 25857 17819 25891
rect 17874 25860 17908 25894
rect 17969 25857 18003 25891
rect 18153 25857 18187 25891
rect 19257 25857 19291 25891
rect 19901 25857 19935 25891
rect 20085 25857 20119 25891
rect 21097 25857 21131 25891
rect 22569 25857 22603 25891
rect 22753 25857 22787 25891
rect 22845 25857 22879 25891
rect 22937 25857 22971 25891
rect 23673 25857 23707 25891
rect 25605 25857 25639 25891
rect 25784 25857 25818 25891
rect 25881 25857 25915 25891
rect 26019 25857 26053 25891
rect 29294 25857 29328 25891
rect 29561 25857 29595 25891
rect 33149 25857 33183 25891
rect 39885 25857 39919 25891
rect 40141 25857 40175 25891
rect 40877 25857 40911 25891
rect 40969 25857 41003 25891
rect 41061 25857 41095 25891
rect 41245 25857 41279 25891
rect 5825 25789 5859 25823
rect 9597 25789 9631 25823
rect 11989 25789 12023 25823
rect 15577 25789 15611 25823
rect 19717 25789 19751 25823
rect 36369 25789 36403 25823
rect 4629 25653 4663 25687
rect 6377 25653 6411 25687
rect 13093 25653 13127 25687
rect 16681 25653 16715 25687
rect 23213 25653 23247 25687
rect 28181 25653 28215 25687
rect 34529 25653 34563 25687
rect 38761 25653 38795 25687
rect 5365 25449 5399 25483
rect 7205 25449 7239 25483
rect 25605 25449 25639 25483
rect 38117 25449 38151 25483
rect 40049 25449 40083 25483
rect 9137 25381 9171 25415
rect 11161 25381 11195 25415
rect 6745 25313 6779 25347
rect 18153 25313 18187 25347
rect 18429 25313 18463 25347
rect 22937 25313 22971 25347
rect 32321 25313 32355 25347
rect 4077 25245 4111 25279
rect 4169 25245 4203 25279
rect 4261 25245 4295 25279
rect 4445 25245 4479 25279
rect 6478 25245 6512 25279
rect 9321 25245 9355 25279
rect 9873 25245 9907 25279
rect 15301 25245 15335 25279
rect 22681 25245 22715 25279
rect 25789 25245 25823 25279
rect 37381 25245 37415 25279
rect 40325 25245 40359 25279
rect 40417 25245 40451 25279
rect 40509 25245 40543 25279
rect 40693 25245 40727 25279
rect 58173 25245 58207 25279
rect 10057 25177 10091 25211
rect 10977 25177 11011 25211
rect 15117 25177 15151 25211
rect 16037 25177 16071 25211
rect 16221 25177 16255 25211
rect 16957 25177 16991 25211
rect 17141 25177 17175 25211
rect 25973 25177 26007 25211
rect 29653 25177 29687 25211
rect 29837 25177 29871 25211
rect 32054 25177 32088 25211
rect 37136 25177 37170 25211
rect 3801 25109 3835 25143
rect 10241 25109 10275 25143
rect 13461 25109 13495 25143
rect 14381 25109 14415 25143
rect 14933 25109 14967 25143
rect 21557 25109 21591 25143
rect 30021 25109 30055 25143
rect 30941 25109 30975 25143
rect 36001 25109 36035 25143
rect 39221 25109 39255 25143
rect 41153 25109 41187 25143
rect 4721 24905 4755 24939
rect 10977 24905 11011 24939
rect 12633 24905 12667 24939
rect 15761 24905 15795 24939
rect 21281 24837 21315 24871
rect 28641 24837 28675 24871
rect 38301 24837 38335 24871
rect 3626 24769 3660 24803
rect 5273 24769 5307 24803
rect 10057 24769 10091 24803
rect 10149 24769 10183 24803
rect 10241 24769 10275 24803
rect 10425 24769 10459 24803
rect 11621 24769 11655 24803
rect 12863 24769 12897 24803
rect 13001 24769 13035 24803
rect 13093 24772 13127 24806
rect 13277 24769 13311 24803
rect 14637 24769 14671 24803
rect 16957 24769 16991 24803
rect 17601 24769 17635 24803
rect 17764 24769 17798 24803
rect 17877 24769 17911 24803
rect 18015 24769 18049 24803
rect 18705 24769 18739 24803
rect 18961 24769 18995 24803
rect 21821 24769 21855 24803
rect 22012 24769 22046 24803
rect 22109 24769 22143 24803
rect 22221 24769 22255 24803
rect 22937 24769 22971 24803
rect 23030 24769 23064 24803
rect 23213 24769 23247 24803
rect 23305 24769 23339 24803
rect 23402 24769 23436 24803
rect 28457 24769 28491 24803
rect 30398 24769 30432 24803
rect 30665 24769 30699 24803
rect 3893 24701 3927 24735
rect 14381 24701 14415 24735
rect 18245 24701 18279 24735
rect 9229 24633 9263 24667
rect 16773 24633 16807 24667
rect 25605 24633 25639 24667
rect 29285 24633 29319 24667
rect 2513 24565 2547 24599
rect 7297 24565 7331 24599
rect 9781 24565 9815 24599
rect 12081 24565 12115 24599
rect 13829 24565 13863 24599
rect 20085 24565 20119 24599
rect 22477 24565 22511 24599
rect 23581 24565 23615 24599
rect 26249 24565 26283 24599
rect 28825 24565 28859 24599
rect 37381 24565 37415 24599
rect 39589 24565 39623 24599
rect 5457 24361 5491 24395
rect 8033 24361 8067 24395
rect 19257 24361 19291 24395
rect 28365 24361 28399 24395
rect 30757 24361 30791 24395
rect 37289 24361 37323 24395
rect 14289 24293 14323 24327
rect 8953 24225 8987 24259
rect 17785 24225 17819 24259
rect 36461 24225 36495 24259
rect 6929 24157 6963 24191
rect 7205 24157 7239 24191
rect 9220 24157 9254 24191
rect 11299 24157 11333 24191
rect 11437 24157 11471 24191
rect 11529 24157 11563 24191
rect 11713 24157 11747 24191
rect 12173 24157 12207 24191
rect 14545 24157 14579 24191
rect 14638 24157 14672 24191
rect 14749 24154 14783 24188
rect 14933 24157 14967 24191
rect 16681 24157 16715 24191
rect 17509 24157 17543 24191
rect 19441 24157 19475 24191
rect 20821 24157 20855 24191
rect 20914 24157 20948 24191
rect 21189 24157 21223 24191
rect 21327 24157 21361 24191
rect 22065 24157 22099 24191
rect 22421 24157 22455 24191
rect 22569 24157 22603 24191
rect 24685 24157 24719 24191
rect 24848 24157 24882 24191
rect 24961 24157 24995 24191
rect 25099 24157 25133 24191
rect 26065 24157 26099 24191
rect 26157 24157 26191 24191
rect 26249 24157 26283 24191
rect 26433 24157 26467 24191
rect 27905 24157 27939 24191
rect 28641 24157 28675 24191
rect 28733 24157 28767 24191
rect 28825 24157 28859 24191
rect 29009 24157 29043 24191
rect 30113 24157 30147 24191
rect 30297 24157 30331 24191
rect 30389 24157 30423 24191
rect 30481 24157 30515 24191
rect 36645 24157 36679 24191
rect 37565 24157 37599 24191
rect 37657 24157 37691 24191
rect 37749 24157 37783 24191
rect 37933 24157 37967 24191
rect 40509 24157 40543 24191
rect 41337 24157 41371 24191
rect 58173 24157 58207 24191
rect 4169 24089 4203 24123
rect 12440 24089 12474 24123
rect 16221 24089 16255 24123
rect 19625 24089 19659 24123
rect 21097 24089 21131 24123
rect 22201 24089 22235 24123
rect 22293 24089 22327 24123
rect 36829 24089 36863 24123
rect 40325 24089 40359 24123
rect 41153 24089 41187 24123
rect 10333 24021 10367 24055
rect 11069 24021 11103 24055
rect 13553 24021 13587 24055
rect 15577 24021 15611 24055
rect 21465 24021 21499 24055
rect 21925 24021 21959 24055
rect 25329 24021 25363 24055
rect 25789 24021 25823 24055
rect 27261 24021 27295 24055
rect 29561 24021 29595 24055
rect 31309 24021 31343 24055
rect 40693 24021 40727 24055
rect 41521 24021 41555 24055
rect 6469 23817 6503 23851
rect 9781 23817 9815 23851
rect 13369 23817 13403 23851
rect 14473 23817 14507 23851
rect 18705 23817 18739 23851
rect 26985 23817 27019 23851
rect 29469 23817 29503 23851
rect 41705 23817 41739 23851
rect 8668 23749 8702 23783
rect 10241 23749 10275 23783
rect 12642 23749 12676 23783
rect 15209 23749 15243 23783
rect 16037 23749 16071 23783
rect 22753 23749 22787 23783
rect 24501 23749 24535 23783
rect 27169 23749 27203 23783
rect 28825 23749 28859 23783
rect 29009 23749 29043 23783
rect 36001 23749 36035 23783
rect 2145 23681 2179 23715
rect 2329 23681 2363 23715
rect 7849 23681 7883 23715
rect 8401 23681 8435 23715
rect 10517 23681 10551 23715
rect 10606 23681 10640 23715
rect 10701 23684 10735 23718
rect 10885 23681 10919 23715
rect 13553 23681 13587 23715
rect 13737 23681 13771 23715
rect 14933 23681 14967 23715
rect 15117 23681 15151 23715
rect 15301 23681 15335 23715
rect 18061 23681 18095 23715
rect 22477 23681 22511 23715
rect 22570 23681 22604 23715
rect 22845 23681 22879 23715
rect 22983 23681 23017 23715
rect 25053 23681 25087 23715
rect 25320 23681 25354 23715
rect 27353 23681 27387 23715
rect 28641 23681 28675 23715
rect 29725 23681 29759 23715
rect 29818 23681 29852 23715
rect 29929 23681 29963 23715
rect 30113 23681 30147 23715
rect 35909 23681 35943 23715
rect 36093 23681 36127 23715
rect 36277 23681 36311 23715
rect 37473 23681 37507 23715
rect 37657 23681 37691 23715
rect 39885 23681 39919 23715
rect 40141 23681 40175 23715
rect 40877 23681 40911 23715
rect 40969 23681 41003 23715
rect 41061 23681 41095 23715
rect 41245 23681 41279 23715
rect 7573 23613 7607 23647
rect 12909 23613 12943 23647
rect 40601 23613 40635 23647
rect 18245 23545 18279 23579
rect 26433 23545 26467 23579
rect 30573 23545 30607 23579
rect 38761 23545 38795 23579
rect 2513 23477 2547 23511
rect 11529 23477 11563 23511
rect 15485 23477 15519 23511
rect 23121 23477 23155 23511
rect 35725 23477 35759 23511
rect 37289 23477 37323 23511
rect 3893 23273 3927 23307
rect 4813 23273 4847 23307
rect 10241 23273 10275 23307
rect 11897 23273 11931 23307
rect 22661 23273 22695 23307
rect 36185 23273 36219 23307
rect 39221 23273 39255 23307
rect 7849 23205 7883 23239
rect 11345 23205 11379 23239
rect 14473 23137 14507 23171
rect 23765 23137 23799 23171
rect 34161 23137 34195 23171
rect 2605 23069 2639 23103
rect 2697 23069 2731 23103
rect 2789 23069 2823 23103
rect 2973 23069 3007 23103
rect 5365 23069 5399 23103
rect 5549 23069 5583 23103
rect 5641 23069 5675 23103
rect 5733 23069 5767 23103
rect 6469 23069 6503 23103
rect 10057 23069 10091 23103
rect 11253 23069 11287 23103
rect 11437 23069 11471 23103
rect 16773 23069 16807 23103
rect 18521 23069 18555 23103
rect 22753 23069 22787 23103
rect 22845 23069 22879 23103
rect 24869 23069 24903 23103
rect 25605 23069 25639 23103
rect 25872 23069 25906 23103
rect 31769 23069 31803 23103
rect 31953 23069 31987 23103
rect 32137 23069 32171 23103
rect 35357 23069 35391 23103
rect 35725 23069 35759 23103
rect 37565 23069 37599 23103
rect 40601 23069 40635 23103
rect 40693 23069 40727 23103
rect 40785 23069 40819 23103
rect 40969 23069 41003 23103
rect 6009 23001 6043 23035
rect 6714 23001 6748 23035
rect 9873 23001 9907 23035
rect 12081 23001 12115 23035
rect 12265 23001 12299 23035
rect 18705 23001 18739 23035
rect 25053 23001 25087 23035
rect 32045 23001 32079 23035
rect 33894 23001 33928 23035
rect 35449 23001 35483 23035
rect 35541 23001 35575 23035
rect 37298 23001 37332 23035
rect 2329 22933 2363 22967
rect 15485 22933 15519 22967
rect 18337 22933 18371 22967
rect 22477 22933 22511 22967
rect 26985 22933 27019 22967
rect 29561 22933 29595 22967
rect 32321 22933 32355 22967
rect 32781 22933 32815 22967
rect 35173 22933 35207 22967
rect 40325 22933 40359 22967
rect 1593 22729 1627 22763
rect 5733 22729 5767 22763
rect 6377 22729 6411 22763
rect 7205 22729 7239 22763
rect 10149 22729 10183 22763
rect 11621 22729 11655 22763
rect 15301 22729 15335 22763
rect 19625 22729 19659 22763
rect 26341 22729 26375 22763
rect 33333 22729 33367 22763
rect 35725 22729 35759 22763
rect 37289 22729 37323 22763
rect 1961 22661 1995 22695
rect 2666 22661 2700 22695
rect 6561 22661 6595 22695
rect 14565 22661 14599 22695
rect 14657 22661 14691 22695
rect 16773 22661 16807 22695
rect 26157 22661 26191 22695
rect 34805 22661 34839 22695
rect 36001 22661 36035 22695
rect 1777 22593 1811 22627
rect 2421 22593 2455 22627
rect 4537 22593 4571 22627
rect 4629 22593 4663 22627
rect 4721 22593 4755 22627
rect 4905 22593 4939 22627
rect 6745 22593 6779 22627
rect 7389 22593 7423 22627
rect 14473 22593 14507 22627
rect 14841 22593 14875 22627
rect 18512 22593 18546 22627
rect 21189 22593 21223 22627
rect 21281 22593 21315 22627
rect 21833 22593 21867 22627
rect 22017 22593 22051 22627
rect 24133 22593 24167 22627
rect 25973 22593 26007 22627
rect 27988 22593 28022 22627
rect 32689 22593 32723 22627
rect 32873 22593 32907 22627
rect 32965 22593 32999 22627
rect 33057 22593 33091 22627
rect 33977 22593 34011 22627
rect 34069 22593 34103 22627
rect 34207 22593 34241 22627
rect 34345 22593 34379 22627
rect 35081 22593 35115 22627
rect 35909 22593 35943 22627
rect 36093 22593 36127 22627
rect 36277 22593 36311 22627
rect 37565 22593 37599 22627
rect 37657 22593 37691 22627
rect 37749 22593 37783 22627
rect 37933 22593 37967 22627
rect 39885 22593 39919 22627
rect 40141 22593 40175 22627
rect 18245 22525 18279 22559
rect 23857 22525 23891 22559
rect 27721 22525 27755 22559
rect 34897 22525 34931 22559
rect 3801 22457 3835 22491
rect 7941 22457 7975 22491
rect 35265 22457 35299 22491
rect 38761 22457 38795 22491
rect 58173 22457 58207 22491
rect 4261 22389 4295 22423
rect 14289 22389 14323 22423
rect 15853 22389 15887 22423
rect 17693 22389 17727 22423
rect 20913 22389 20947 22423
rect 21097 22389 21131 22423
rect 21833 22389 21867 22423
rect 22201 22389 22235 22423
rect 22661 22389 22695 22423
rect 23305 22389 23339 22423
rect 29101 22389 29135 22423
rect 32137 22389 32171 22423
rect 33793 22389 33827 22423
rect 34805 22389 34839 22423
rect 9321 22185 9355 22219
rect 19993 22185 20027 22219
rect 33517 22185 33551 22219
rect 37473 22185 37507 22219
rect 7389 22117 7423 22151
rect 18521 22117 18555 22151
rect 21833 22117 21867 22151
rect 6009 22049 6043 22083
rect 16773 22049 16807 22083
rect 19901 22049 19935 22083
rect 1869 21981 1903 22015
rect 3801 21981 3835 22015
rect 9873 21981 9907 22015
rect 10241 21981 10275 22015
rect 11253 21981 11287 22015
rect 11529 21981 11563 22015
rect 11621 21981 11655 22015
rect 15577 21981 15611 22015
rect 15761 21981 15795 22015
rect 17049 21981 17083 22015
rect 17877 21981 17911 22015
rect 18061 21981 18095 22015
rect 18153 21981 18187 22015
rect 18245 21981 18279 22015
rect 19993 21981 20027 22015
rect 23029 21981 23063 22015
rect 23118 21975 23152 22009
rect 23213 21981 23247 22015
rect 23397 21981 23431 22015
rect 24501 21981 24535 22015
rect 28457 21981 28491 22015
rect 32045 21981 32079 22015
rect 32229 21981 32263 22015
rect 32413 21981 32447 22015
rect 33241 21981 33275 22015
rect 33333 21981 33367 22015
rect 33517 21981 33551 22015
rect 2136 21913 2170 21947
rect 4068 21913 4102 21947
rect 6276 21913 6310 21947
rect 9229 21913 9263 21947
rect 10057 21913 10091 21947
rect 10149 21913 10183 21947
rect 11437 21913 11471 21947
rect 15393 21913 15427 21947
rect 20545 21913 20579 21947
rect 28273 21913 28307 21947
rect 32321 21913 32355 21947
rect 3249 21845 3283 21879
rect 5181 21845 5215 21879
rect 10425 21845 10459 21879
rect 11805 21845 11839 21879
rect 14933 21845 14967 21879
rect 19625 21845 19659 21879
rect 22753 21845 22787 21879
rect 24685 21845 24719 21879
rect 28641 21845 28675 21879
rect 32597 21845 32631 21879
rect 33057 21845 33091 21879
rect 36921 21845 36955 21879
rect 40325 21845 40359 21879
rect 2237 21641 2271 21675
rect 4169 21641 4203 21675
rect 6377 21641 6411 21675
rect 7481 21641 7515 21675
rect 12173 21641 12207 21675
rect 21097 21641 21131 21675
rect 23765 21641 23799 21675
rect 28089 21641 28123 21675
rect 32597 21641 32631 21675
rect 33057 21641 33091 21675
rect 3985 21573 4019 21607
rect 5641 21573 5675 21607
rect 5825 21573 5859 21607
rect 10241 21573 10275 21607
rect 15301 21573 15335 21607
rect 18521 21573 18555 21607
rect 24133 21573 24167 21607
rect 30389 21573 30423 21607
rect 32413 21573 32447 21607
rect 33517 21573 33551 21607
rect 39712 21573 39746 21607
rect 40417 21573 40451 21607
rect 2513 21505 2547 21539
rect 2605 21505 2639 21539
rect 2697 21505 2731 21539
rect 2881 21505 2915 21539
rect 3801 21505 3835 21539
rect 5457 21505 5491 21539
rect 6607 21505 6641 21539
rect 6745 21505 6779 21539
rect 6837 21505 6871 21539
rect 7021 21505 7055 21539
rect 9965 21505 9999 21539
rect 10149 21505 10183 21539
rect 10333 21505 10367 21539
rect 12265 21505 12299 21539
rect 14841 21505 14875 21539
rect 15485 21505 15519 21539
rect 16948 21505 16982 21539
rect 18705 21505 18739 21539
rect 21189 21505 21223 21539
rect 22661 21505 22695 21539
rect 22845 21505 22879 21539
rect 22937 21505 22971 21539
rect 23029 21505 23063 21539
rect 23949 21505 23983 21539
rect 26433 21505 26467 21539
rect 28319 21505 28353 21539
rect 28454 21505 28488 21539
rect 28570 21511 28604 21545
rect 28733 21505 28767 21539
rect 30113 21505 30147 21539
rect 32229 21505 32263 21539
rect 33241 21505 33275 21539
rect 40693 21505 40727 21539
rect 40785 21505 40819 21539
rect 40877 21505 40911 21539
rect 41061 21505 41095 21539
rect 15669 21437 15703 21471
rect 16681 21437 16715 21471
rect 22201 21437 22235 21471
rect 29193 21437 29227 21471
rect 30297 21437 30331 21471
rect 33425 21437 33459 21471
rect 39957 21437 39991 21471
rect 10517 21369 10551 21403
rect 18061 21369 18095 21403
rect 20361 21369 20395 21403
rect 29929 21369 29963 21403
rect 8953 21301 8987 21335
rect 14197 21301 14231 21335
rect 14657 21301 14691 21335
rect 18889 21301 18923 21335
rect 19809 21301 19843 21335
rect 23305 21301 23339 21335
rect 25145 21301 25179 21335
rect 26985 21301 27019 21335
rect 27629 21301 27663 21335
rect 30113 21301 30147 21335
rect 33241 21301 33275 21335
rect 38577 21301 38611 21335
rect 58173 21301 58207 21335
rect 10885 21097 10919 21131
rect 14657 21097 14691 21131
rect 16589 21097 16623 21131
rect 17049 21097 17083 21131
rect 30113 21097 30147 21131
rect 36553 21097 36587 21131
rect 40601 21097 40635 21131
rect 11621 21029 11655 21063
rect 16037 21029 16071 21063
rect 21373 21029 21407 21063
rect 10241 20893 10275 20927
rect 10793 20893 10827 20927
rect 11437 20893 11471 20927
rect 12817 20893 12851 20927
rect 15393 20893 15427 20927
rect 15486 20893 15520 20927
rect 15669 20893 15703 20927
rect 15899 20893 15933 20927
rect 17305 20893 17339 20927
rect 17398 20887 17432 20921
rect 17509 20893 17543 20927
rect 17693 20893 17727 20927
rect 20131 20893 20165 20927
rect 20489 20893 20523 20927
rect 20637 20893 20671 20927
rect 21189 20893 21223 20927
rect 22477 20893 22511 20927
rect 26157 20893 26191 20927
rect 29561 20893 29595 20927
rect 29929 20893 29963 20927
rect 36737 20893 36771 20927
rect 37105 20893 37139 20927
rect 39313 20893 39347 20927
rect 40233 20893 40267 20927
rect 40417 20893 40451 20927
rect 13001 20825 13035 20859
rect 14565 20825 14599 20859
rect 15761 20825 15795 20859
rect 20269 20825 20303 20859
rect 20361 20825 20395 20859
rect 22744 20825 22778 20859
rect 25973 20825 26007 20859
rect 29745 20825 29779 20859
rect 29837 20825 29871 20859
rect 36829 20825 36863 20859
rect 36921 20825 36955 20859
rect 39068 20825 39102 20859
rect 3065 20757 3099 20791
rect 12173 20757 12207 20791
rect 13185 20757 13219 20791
rect 19993 20757 20027 20791
rect 22017 20757 22051 20791
rect 23857 20757 23891 20791
rect 26341 20757 26375 20791
rect 27261 20757 27295 20791
rect 32413 20757 32447 20791
rect 37933 20757 37967 20791
rect 7757 20553 7791 20587
rect 13645 20553 13679 20587
rect 15669 20553 15703 20587
rect 33609 20553 33643 20587
rect 40509 20553 40543 20587
rect 20269 20485 20303 20519
rect 23296 20485 23330 20519
rect 33149 20485 33183 20519
rect 34722 20485 34756 20519
rect 40049 20485 40083 20519
rect 7849 20417 7883 20451
rect 8401 20417 8435 20451
rect 9597 20417 9631 20451
rect 12532 20417 12566 20451
rect 14381 20417 14415 20451
rect 15577 20417 15611 20451
rect 17693 20417 17727 20451
rect 17785 20417 17819 20451
rect 20039 20417 20073 20451
rect 20177 20417 20211 20451
rect 20397 20417 20431 20451
rect 20545 20417 20579 20451
rect 23029 20417 23063 20451
rect 25329 20417 25363 20451
rect 26065 20417 26099 20451
rect 26157 20417 26191 20451
rect 26249 20417 26283 20451
rect 26433 20417 26467 20451
rect 27537 20417 27571 20451
rect 28641 20417 28675 20451
rect 29101 20417 29135 20451
rect 30113 20417 30147 20451
rect 32505 20417 32539 20451
rect 32689 20417 32723 20451
rect 32781 20417 32815 20451
rect 32873 20417 32907 20451
rect 36185 20417 36219 20451
rect 40785 20417 40819 20451
rect 40877 20417 40911 20451
rect 40969 20417 41003 20451
rect 41153 20417 41187 20451
rect 9505 20349 9539 20383
rect 12265 20349 12299 20383
rect 14105 20349 14139 20383
rect 29837 20349 29871 20383
rect 34989 20349 35023 20383
rect 35909 20349 35943 20383
rect 27721 20281 27755 20315
rect 9229 20213 9263 20247
rect 9413 20213 9447 20247
rect 10149 20213 10183 20247
rect 11621 20213 11655 20247
rect 17417 20213 17451 20247
rect 17601 20213 17635 20247
rect 19901 20213 19935 20247
rect 24409 20213 24443 20247
rect 25789 20213 25823 20247
rect 29285 20213 29319 20247
rect 11989 20009 12023 20043
rect 12541 20009 12575 20043
rect 14933 20009 14967 20043
rect 19533 20009 19567 20043
rect 23305 20009 23339 20043
rect 26985 20009 27019 20043
rect 29883 20009 29917 20043
rect 33149 20009 33183 20043
rect 36415 20009 36449 20043
rect 40601 20009 40635 20043
rect 8401 19805 8435 19839
rect 12817 19805 12851 19839
rect 12909 19805 12943 19839
rect 13001 19805 13035 19839
rect 13185 19805 13219 19839
rect 14841 19805 14875 19839
rect 14933 19805 14967 19839
rect 19712 19805 19746 19839
rect 20084 19805 20118 19839
rect 20177 19805 20211 19839
rect 23489 19805 23523 19839
rect 25605 19805 25639 19839
rect 25872 19805 25906 19839
rect 28457 19805 28491 19839
rect 28733 19805 28767 19839
rect 28825 19805 28859 19839
rect 29653 19805 29687 19839
rect 31125 19805 31159 19839
rect 31493 19805 31527 19839
rect 32965 19805 32999 19839
rect 35357 19805 35391 19839
rect 35725 19805 35759 19839
rect 36185 19805 36219 19839
rect 39313 19805 39347 19839
rect 40233 19805 40267 19839
rect 40417 19805 40451 19839
rect 58173 19805 58207 19839
rect 6469 19737 6503 19771
rect 8134 19737 8168 19771
rect 19809 19737 19843 19771
rect 19901 19737 19935 19771
rect 23673 19737 23707 19771
rect 28641 19737 28675 19771
rect 31217 19737 31251 19771
rect 31309 19737 31343 19771
rect 32781 19737 32815 19771
rect 35449 19737 35483 19771
rect 35541 19737 35575 19771
rect 39068 19737 39102 19771
rect 4629 19669 4663 19703
rect 5917 19669 5951 19703
rect 7021 19669 7055 19703
rect 14565 19669 14599 19703
rect 27445 19669 27479 19703
rect 29009 19669 29043 19703
rect 30941 19669 30975 19703
rect 35173 19669 35207 19703
rect 37933 19669 37967 19703
rect 6561 19465 6595 19499
rect 7849 19465 7883 19499
rect 14105 19465 14139 19499
rect 18061 19465 18095 19499
rect 22017 19465 22051 19499
rect 25973 19465 26007 19499
rect 26985 19465 27019 19499
rect 35909 19465 35943 19499
rect 39313 19465 39347 19499
rect 40601 19465 40635 19499
rect 6469 19397 6503 19431
rect 14657 19397 14691 19431
rect 25605 19397 25639 19431
rect 27445 19397 27479 19431
rect 29745 19397 29779 19431
rect 31033 19397 31067 19431
rect 36277 19397 36311 19431
rect 2421 19329 2455 19363
rect 4629 19329 4663 19363
rect 5457 19329 5491 19363
rect 7113 19329 7147 19363
rect 7297 19329 7331 19363
rect 7665 19329 7699 19363
rect 8677 19329 8711 19363
rect 14013 19329 14047 19363
rect 14197 19329 14231 19363
rect 16681 19329 16715 19363
rect 16937 19329 16971 19363
rect 21925 19329 21959 19363
rect 22109 19329 22143 19363
rect 25421 19329 25455 19363
rect 25697 19329 25731 19363
rect 25789 19329 25823 19363
rect 27169 19329 27203 19363
rect 29561 19329 29595 19363
rect 29837 19329 29871 19363
rect 29929 19329 29963 19363
rect 30757 19329 30791 19363
rect 33342 19329 33376 19363
rect 33609 19329 33643 19363
rect 36093 19329 36127 19363
rect 36185 19329 36219 19363
rect 36461 19329 36495 19363
rect 37565 19329 37599 19363
rect 38025 19329 38059 19363
rect 40877 19329 40911 19363
rect 40969 19329 41003 19363
rect 41061 19329 41095 19363
rect 41245 19329 41279 19363
rect 7389 19261 7423 19295
rect 7481 19261 7515 19295
rect 8585 19261 8619 19295
rect 9229 19261 9263 19295
rect 22569 19261 22603 19295
rect 27261 19261 27295 19295
rect 30849 19261 30883 19295
rect 32229 19193 32263 19227
rect 2237 19125 2271 19159
rect 5365 19125 5399 19159
rect 8309 19125 8343 19159
rect 8493 19125 8527 19159
rect 10885 19125 10919 19159
rect 11529 19125 11563 19159
rect 27353 19125 27387 19159
rect 30113 19125 30147 19159
rect 30573 19125 30607 19159
rect 31033 19125 31067 19159
rect 5641 18921 5675 18955
rect 6377 18921 6411 18955
rect 15853 18921 15887 18955
rect 16405 18921 16439 18955
rect 20637 18921 20671 18955
rect 30113 18921 30147 18955
rect 30757 18921 30791 18955
rect 32781 18921 32815 18955
rect 37289 18921 37323 18955
rect 40233 18921 40267 18955
rect 3249 18853 3283 18887
rect 4261 18785 4295 18819
rect 4445 18785 4479 18819
rect 11437 18785 11471 18819
rect 17601 18785 17635 18819
rect 21925 18785 21959 18819
rect 23305 18785 23339 18819
rect 1869 18717 1903 18751
rect 2136 18717 2170 18751
rect 5365 18717 5399 18751
rect 5457 18717 5491 18751
rect 6929 18717 6963 18751
rect 7113 18717 7147 18751
rect 7205 18717 7239 18751
rect 7297 18717 7331 18751
rect 7481 18717 7515 18751
rect 8125 18717 8159 18751
rect 9597 18717 9631 18751
rect 9864 18717 9898 18751
rect 11713 18717 11747 18751
rect 11805 18717 11839 18751
rect 11897 18717 11931 18751
rect 12081 18717 12115 18751
rect 16681 18717 16715 18751
rect 16773 18717 16807 18751
rect 16865 18717 16899 18751
rect 17049 18717 17083 18751
rect 18061 18717 18095 18751
rect 18245 18717 18279 18751
rect 18337 18717 18371 18751
rect 18429 18717 18463 18751
rect 19257 18717 19291 18751
rect 21649 18717 21683 18751
rect 23029 18717 23063 18751
rect 29837 18717 29871 18751
rect 29929 18717 29963 18751
rect 30113 18717 30147 18751
rect 30757 18717 30791 18751
rect 30849 18717 30883 18751
rect 32125 18717 32159 18751
rect 32300 18717 32334 18751
rect 32416 18717 32450 18751
rect 32505 18717 32539 18751
rect 37473 18717 37507 18751
rect 37565 18717 37599 18751
rect 37841 18717 37875 18751
rect 40049 18717 40083 18751
rect 58173 18717 58207 18751
rect 6285 18649 6319 18683
rect 12541 18649 12575 18683
rect 19502 18649 19536 18683
rect 27353 18649 27387 18683
rect 31033 18649 31067 18683
rect 37657 18649 37691 18683
rect 39865 18649 39899 18683
rect 3801 18581 3835 18615
rect 4169 18581 4203 18615
rect 4997 18581 5031 18615
rect 7665 18581 7699 18615
rect 10977 18581 11011 18615
rect 18705 18581 18739 18615
rect 26709 18581 26743 18615
rect 27445 18581 27479 18615
rect 29653 18581 29687 18615
rect 30573 18581 30607 18615
rect 31677 18581 31711 18615
rect 40693 18581 40727 18615
rect 41521 18581 41555 18615
rect 2329 18377 2363 18411
rect 5181 18377 5215 18411
rect 11897 18377 11931 18411
rect 14933 18377 14967 18411
rect 17049 18377 17083 18411
rect 18981 18377 19015 18411
rect 32505 18377 32539 18411
rect 38025 18377 38059 18411
rect 3709 18309 3743 18343
rect 4537 18309 4571 18343
rect 7858 18309 7892 18343
rect 11713 18309 11747 18343
rect 32137 18309 32171 18343
rect 32965 18309 32999 18343
rect 33149 18309 33183 18343
rect 36553 18309 36587 18343
rect 38117 18309 38151 18343
rect 1685 18241 1719 18275
rect 2513 18241 2547 18275
rect 4905 18241 4939 18275
rect 10609 18241 10643 18275
rect 10701 18241 10735 18275
rect 10793 18241 10827 18275
rect 10977 18241 11011 18275
rect 11529 18241 11563 18275
rect 12633 18241 12667 18275
rect 13185 18241 13219 18275
rect 13369 18241 13403 18275
rect 13461 18241 13495 18275
rect 13553 18241 13587 18275
rect 14289 18241 14323 18275
rect 14382 18241 14416 18275
rect 14565 18241 14599 18275
rect 14657 18241 14691 18275
rect 14754 18241 14788 18275
rect 17233 18241 17267 18275
rect 17417 18241 17451 18275
rect 19165 18241 19199 18275
rect 19349 18241 19383 18275
rect 21189 18241 21223 18275
rect 22017 18241 22051 18275
rect 23397 18241 23431 18275
rect 24501 18241 24535 18275
rect 24685 18241 24719 18275
rect 24777 18241 24811 18275
rect 24869 18241 24903 18275
rect 29101 18241 29135 18275
rect 29653 18241 29687 18275
rect 32321 18241 32355 18275
rect 36369 18241 36403 18275
rect 36461 18241 36495 18275
rect 36737 18241 36771 18275
rect 40069 18241 40103 18275
rect 40325 18241 40359 18275
rect 41061 18241 41095 18275
rect 41153 18241 41187 18275
rect 41245 18241 41279 18275
rect 41429 18241 41463 18275
rect 2697 18173 2731 18207
rect 3801 18173 3835 18207
rect 3985 18173 4019 18207
rect 4997 18173 5031 18207
rect 8125 18173 8159 18207
rect 22201 18173 22235 18207
rect 22661 18173 22695 18207
rect 40785 18173 40819 18207
rect 5825 18105 5859 18139
rect 9873 18105 9907 18139
rect 21005 18105 21039 18139
rect 21833 18105 21867 18139
rect 36185 18105 36219 18139
rect 1869 18037 1903 18071
rect 3341 18037 3375 18071
rect 6745 18037 6779 18071
rect 9229 18037 9263 18071
rect 10333 18037 10367 18071
rect 13829 18037 13863 18071
rect 23489 18037 23523 18071
rect 25053 18037 25087 18071
rect 29745 18037 29779 18071
rect 33333 18037 33367 18071
rect 38945 18037 38979 18071
rect 2145 17833 2179 17867
rect 4169 17833 4203 17867
rect 6745 17833 6779 17867
rect 19717 17833 19751 17867
rect 25973 17833 26007 17867
rect 33885 17833 33919 17867
rect 37473 17833 37507 17867
rect 40785 17833 40819 17867
rect 4905 17765 4939 17799
rect 5733 17765 5767 17799
rect 21189 17765 21223 17799
rect 31401 17765 31435 17799
rect 14105 17697 14139 17731
rect 19809 17697 19843 17731
rect 22569 17697 22603 17731
rect 24593 17697 24627 17731
rect 32321 17697 32355 17731
rect 36093 17697 36127 17731
rect 38209 17697 38243 17731
rect 41245 17697 41279 17731
rect 2329 17629 2363 17663
rect 2421 17629 2455 17663
rect 3249 17629 3283 17663
rect 4721 17629 4755 17663
rect 5549 17629 5583 17663
rect 7021 17629 7055 17663
rect 7573 17629 7607 17663
rect 10609 17629 10643 17663
rect 13047 17629 13081 17663
rect 13166 17629 13200 17663
rect 13277 17626 13311 17660
rect 13461 17629 13495 17663
rect 14361 17629 14395 17663
rect 19901 17629 19935 17663
rect 20545 17629 20579 17663
rect 23029 17629 23063 17663
rect 23305 17629 23339 17663
rect 26617 17629 26651 17663
rect 31217 17629 31251 17663
rect 31953 17629 31987 17663
rect 32781 17629 32815 17663
rect 32944 17629 32978 17663
rect 33057 17629 33091 17663
rect 33169 17629 33203 17663
rect 37933 17629 37967 17663
rect 40601 17629 40635 17663
rect 20361 17561 20395 17595
rect 20729 17561 20763 17595
rect 22302 17561 22336 17595
rect 24860 17561 24894 17595
rect 26801 17561 26835 17595
rect 32137 17561 32171 17595
rect 36360 17561 36394 17595
rect 40417 17561 40451 17595
rect 12081 17493 12115 17527
rect 12817 17493 12851 17527
rect 15485 17493 15519 17527
rect 19533 17493 19567 17527
rect 26433 17493 26467 17527
rect 33425 17493 33459 17527
rect 11529 17289 11563 17323
rect 13001 17289 13035 17323
rect 13921 17289 13955 17323
rect 16681 17289 16715 17323
rect 21833 17289 21867 17323
rect 25697 17289 25731 17323
rect 34989 17289 35023 17323
rect 36369 17289 36403 17323
rect 2697 17221 2731 17255
rect 6745 17221 6779 17255
rect 12633 17221 12667 17255
rect 14289 17221 14323 17255
rect 33149 17221 33183 17255
rect 33854 17221 33888 17255
rect 37473 17221 37507 17255
rect 37657 17221 37691 17255
rect 4445 17153 4479 17187
rect 7113 17153 7147 17187
rect 9597 17153 9631 17187
rect 9864 17153 9898 17187
rect 11713 17153 11747 17187
rect 11897 17153 11931 17187
rect 12817 17153 12851 17187
rect 14105 17153 14139 17187
rect 15209 17153 15243 17187
rect 22063 17153 22097 17187
rect 22182 17159 22216 17193
rect 22293 17156 22327 17190
rect 22477 17153 22511 17187
rect 25973 17153 26007 17187
rect 26062 17159 26096 17193
rect 26157 17153 26191 17187
rect 26341 17153 26375 17187
rect 27241 17153 27275 17187
rect 30021 17153 30055 17187
rect 30205 17153 30239 17187
rect 32505 17153 32539 17187
rect 32689 17153 32723 17187
rect 32781 17153 32815 17187
rect 32919 17153 32953 17187
rect 35725 17153 35759 17187
rect 35888 17153 35922 17187
rect 36001 17153 36035 17187
rect 36113 17153 36147 17187
rect 38761 17153 38795 17187
rect 14933 17085 14967 17119
rect 23029 17085 23063 17119
rect 23673 17085 23707 17119
rect 23949 17085 23983 17119
rect 26985 17085 27019 17119
rect 33609 17085 33643 17119
rect 37289 17085 37323 17119
rect 39037 17085 39071 17119
rect 10977 17017 11011 17051
rect 17509 17017 17543 17051
rect 58173 17017 58207 17051
rect 5181 16949 5215 16983
rect 5825 16949 5859 16983
rect 21281 16949 21315 16983
rect 25145 16949 25179 16983
rect 28365 16949 28399 16983
rect 29837 16949 29871 16983
rect 31585 16949 31619 16983
rect 3249 16745 3283 16779
rect 4997 16745 5031 16779
rect 24869 16745 24903 16779
rect 25053 16745 25087 16779
rect 26801 16745 26835 16779
rect 27445 16745 27479 16779
rect 34161 16745 34195 16779
rect 36277 16745 36311 16779
rect 39129 16745 39163 16779
rect 4353 16677 4387 16711
rect 11621 16677 11655 16711
rect 12173 16677 12207 16711
rect 20361 16677 20395 16711
rect 1869 16609 1903 16643
rect 8401 16609 8435 16643
rect 12725 16609 12759 16643
rect 14841 16609 14875 16643
rect 20821 16609 20855 16643
rect 22845 16609 22879 16643
rect 25145 16609 25179 16643
rect 27813 16609 27847 16643
rect 32781 16609 32815 16643
rect 2125 16541 2159 16575
rect 4169 16541 4203 16575
rect 10977 16541 11011 16575
rect 11070 16541 11104 16575
rect 11483 16541 11517 16575
rect 15669 16541 15703 16575
rect 15761 16541 15795 16575
rect 15853 16541 15887 16575
rect 16037 16541 16071 16575
rect 16497 16541 16531 16575
rect 16681 16541 16715 16575
rect 16773 16541 16807 16575
rect 16865 16541 16899 16575
rect 17601 16541 17635 16575
rect 17785 16541 17819 16575
rect 17877 16541 17911 16575
rect 17969 16541 18003 16575
rect 23121 16541 23155 16575
rect 25053 16541 25087 16575
rect 25329 16541 25363 16575
rect 26163 16541 26197 16575
rect 26341 16541 26375 16575
rect 26433 16541 26467 16575
rect 26525 16541 26559 16575
rect 27629 16541 27663 16575
rect 29653 16541 29687 16575
rect 31493 16541 31527 16575
rect 31769 16541 31803 16575
rect 37013 16541 37047 16575
rect 37105 16541 37139 16575
rect 37381 16541 37415 16575
rect 40049 16541 40083 16575
rect 8134 16473 8168 16507
rect 11253 16473 11287 16507
rect 11345 16473 11379 16507
rect 29898 16473 29932 16507
rect 33048 16473 33082 16507
rect 37197 16473 37231 16507
rect 39221 16473 39255 16507
rect 39865 16473 39899 16507
rect 7021 16405 7055 16439
rect 10425 16405 10459 16439
rect 13185 16405 13219 16439
rect 15393 16405 15427 16439
rect 17141 16405 17175 16439
rect 18245 16405 18279 16439
rect 19257 16405 19291 16439
rect 31033 16405 31067 16439
rect 35633 16405 35667 16439
rect 36829 16405 36863 16439
rect 40233 16405 40267 16439
rect 10057 16201 10091 16235
rect 10701 16201 10735 16235
rect 12173 16201 12207 16235
rect 12725 16201 12759 16235
rect 16773 16201 16807 16235
rect 17601 16201 17635 16235
rect 18797 16201 18831 16235
rect 20729 16201 20763 16235
rect 22477 16201 22511 16235
rect 25053 16201 25087 16235
rect 26065 16201 26099 16235
rect 28917 16201 28951 16235
rect 33793 16201 33827 16235
rect 40233 16201 40267 16235
rect 3709 16133 3743 16167
rect 11805 16133 11839 16167
rect 11897 16133 11931 16167
rect 17141 16133 17175 16167
rect 17969 16133 18003 16167
rect 18981 16133 19015 16167
rect 26249 16133 26283 16167
rect 26433 16133 26467 16167
rect 2237 16065 2271 16099
rect 3617 16065 3651 16099
rect 9965 16065 9999 16099
rect 10149 16065 10183 16099
rect 10609 16065 10643 16099
rect 10793 16065 10827 16099
rect 11529 16065 11563 16099
rect 11622 16065 11656 16099
rect 11994 16065 12028 16099
rect 12633 16065 12667 16099
rect 12817 16065 12851 16099
rect 14289 16065 14323 16099
rect 16957 16065 16991 16099
rect 17785 16065 17819 16099
rect 19165 16065 19199 16099
rect 20637 16065 20671 16099
rect 20821 16065 20855 16099
rect 22385 16065 22419 16099
rect 22569 16065 22603 16099
rect 23213 16065 23247 16099
rect 25605 16065 25639 16099
rect 29193 16065 29227 16099
rect 29285 16065 29319 16099
rect 29377 16065 29411 16099
rect 29561 16065 29595 16099
rect 31309 16065 31343 16099
rect 32505 16065 32539 16099
rect 35541 16065 35575 16099
rect 38853 16065 38887 16099
rect 39120 16065 39154 16099
rect 40969 16065 41003 16099
rect 3893 15997 3927 16031
rect 14565 15997 14599 16031
rect 23489 15997 23523 16031
rect 30021 15997 30055 16031
rect 30297 15997 30331 16031
rect 35265 15997 35299 16031
rect 40693 15997 40727 16031
rect 1777 15929 1811 15963
rect 20085 15929 20119 15963
rect 2421 15861 2455 15895
rect 3249 15861 3283 15895
rect 4537 15861 4571 15895
rect 7665 15861 7699 15895
rect 9413 15861 9447 15895
rect 13829 15861 13863 15895
rect 21833 15861 21867 15895
rect 27261 15861 27295 15895
rect 28365 15861 28399 15895
rect 31493 15861 31527 15895
rect 58173 15861 58207 15895
rect 2145 15657 2179 15691
rect 7573 15657 7607 15691
rect 8401 15657 8435 15691
rect 10241 15657 10275 15691
rect 12173 15657 12207 15691
rect 14289 15657 14323 15691
rect 19441 15657 19475 15691
rect 19901 15657 19935 15691
rect 22109 15657 22143 15691
rect 22753 15657 22787 15691
rect 27445 15657 27479 15691
rect 30941 15657 30975 15691
rect 38301 15657 38335 15691
rect 39865 15657 39899 15691
rect 20637 15589 20671 15623
rect 3801 15521 3835 15555
rect 6285 15521 6319 15555
rect 7113 15521 7147 15555
rect 7205 15521 7239 15555
rect 18705 15521 18739 15555
rect 35449 15521 35483 15555
rect 35725 15521 35759 15555
rect 2329 15453 2363 15487
rect 2421 15453 2455 15487
rect 3065 15453 3099 15487
rect 6009 15453 6043 15487
rect 6101 15453 6135 15487
rect 6837 15453 6871 15487
rect 7021 15453 7055 15487
rect 7389 15453 7423 15487
rect 8309 15453 8343 15487
rect 8401 15453 8435 15487
rect 13553 15453 13587 15487
rect 14105 15453 14139 15487
rect 14289 15453 14323 15487
rect 15117 15453 15151 15487
rect 15384 15453 15418 15487
rect 19257 15453 19291 15487
rect 19441 15453 19475 15487
rect 20453 15453 20487 15487
rect 20637 15453 20671 15487
rect 21465 15453 21499 15487
rect 22569 15453 22603 15487
rect 22753 15453 22787 15487
rect 27353 15453 27387 15487
rect 27537 15453 27571 15487
rect 29561 15453 29595 15487
rect 31585 15453 31619 15487
rect 33241 15453 33275 15487
rect 33517 15453 33551 15487
rect 37473 15453 37507 15487
rect 40141 15453 40175 15487
rect 40233 15453 40267 15487
rect 40325 15453 40359 15487
rect 40509 15453 40543 15487
rect 4046 15385 4080 15419
rect 13286 15385 13320 15419
rect 16957 15385 16991 15419
rect 23305 15385 23339 15419
rect 24409 15385 24443 15419
rect 27997 15385 28031 15419
rect 29806 15385 29840 15419
rect 31401 15385 31435 15419
rect 34713 15385 34747 15419
rect 37657 15385 37691 15419
rect 40969 15385 41003 15419
rect 3249 15317 3283 15351
rect 5181 15317 5215 15351
rect 5641 15317 5675 15351
rect 8033 15317 8067 15351
rect 10977 15317 11011 15351
rect 16497 15317 16531 15351
rect 31769 15317 31803 15351
rect 32413 15317 32447 15351
rect 37841 15317 37875 15351
rect 38853 15317 38887 15351
rect 3801 15113 3835 15147
rect 4261 15113 4295 15147
rect 7021 15113 7055 15147
rect 17233 15113 17267 15147
rect 19717 15113 19751 15147
rect 20729 15113 20763 15147
rect 21189 15113 21223 15147
rect 29653 15113 29687 15147
rect 36185 15113 36219 15147
rect 40233 15113 40267 15147
rect 9505 15045 9539 15079
rect 12909 15045 12943 15079
rect 22845 15045 22879 15079
rect 22937 15045 22971 15079
rect 38393 15045 38427 15079
rect 39098 15045 39132 15079
rect 40969 15045 41003 15079
rect 2421 14977 2455 15011
rect 2677 14977 2711 15011
rect 4445 14977 4479 15011
rect 7389 14977 7423 15011
rect 9413 14977 9447 15011
rect 9597 14977 9631 15011
rect 10425 14977 10459 15011
rect 12633 14977 12667 15011
rect 12726 14977 12760 15011
rect 13001 14977 13035 15011
rect 13139 14977 13173 15011
rect 17141 14977 17175 15011
rect 17325 14977 17359 15011
rect 18337 14977 18371 15011
rect 18593 14977 18627 15011
rect 20545 14977 20579 15011
rect 22017 14977 22051 15011
rect 22201 14977 22235 15011
rect 22661 14977 22695 15011
rect 23029 14977 23063 15011
rect 23673 14977 23707 15011
rect 23857 14977 23891 15011
rect 27169 14977 27203 15011
rect 27353 14977 27387 15011
rect 29883 14977 29917 15011
rect 30021 14977 30055 15011
rect 30134 14983 30168 15017
rect 30309 14977 30343 15011
rect 33333 14977 33367 15011
rect 33609 14977 33643 15011
rect 35081 14977 35115 15011
rect 36001 14977 36035 15011
rect 37749 14977 37783 15011
rect 37928 14977 37962 15011
rect 38028 14977 38062 15011
rect 38163 14977 38197 15011
rect 40785 14977 40819 15011
rect 4629 14909 4663 14943
rect 7297 14909 7331 14943
rect 10333 14909 10367 14943
rect 17877 14909 17911 14943
rect 20361 14909 20395 14943
rect 24317 14909 24351 14943
rect 35357 14909 35391 14943
rect 35817 14909 35851 14943
rect 36645 14909 36679 14943
rect 38853 14909 38887 14943
rect 13277 14841 13311 14875
rect 22201 14841 22235 14875
rect 7205 14773 7239 14807
rect 8861 14773 8895 14807
rect 10057 14773 10091 14807
rect 10425 14773 10459 14807
rect 13921 14773 13955 14807
rect 16037 14773 16071 14807
rect 23213 14773 23247 14807
rect 23857 14773 23891 14807
rect 26985 14773 27019 14807
rect 29101 14773 29135 14807
rect 4629 14569 4663 14603
rect 21833 14569 21867 14603
rect 36093 14569 36127 14603
rect 9045 14501 9079 14535
rect 18245 14501 18279 14535
rect 24501 14501 24535 14535
rect 25053 14501 25087 14535
rect 5089 14433 5123 14467
rect 5181 14433 5215 14467
rect 6469 14433 6503 14467
rect 7941 14433 7975 14467
rect 19901 14433 19935 14467
rect 20453 14433 20487 14467
rect 20729 14433 20763 14467
rect 33333 14433 33367 14467
rect 33793 14433 33827 14467
rect 6193 14365 6227 14399
rect 6285 14365 6319 14399
rect 7665 14365 7699 14399
rect 7849 14365 7883 14399
rect 8033 14365 8067 14399
rect 8217 14365 8251 14399
rect 14105 14365 14139 14399
rect 16865 14365 16899 14399
rect 19809 14365 19843 14399
rect 19993 14365 20027 14399
rect 21741 14365 21775 14399
rect 21925 14365 21959 14399
rect 22753 14365 22787 14399
rect 22937 14365 22971 14399
rect 23121 14365 23155 14399
rect 26433 14365 26467 14399
rect 26893 14365 26927 14399
rect 29561 14365 29595 14399
rect 33977 14365 34011 14399
rect 34713 14365 34747 14399
rect 34989 14365 35023 14399
rect 36001 14365 36035 14399
rect 36185 14365 36219 14399
rect 37289 14365 37323 14399
rect 37565 14365 37599 14399
rect 38393 14365 38427 14399
rect 39221 14365 39255 14399
rect 58173 14365 58207 14399
rect 9781 14297 9815 14331
rect 17132 14297 17166 14331
rect 23029 14297 23063 14331
rect 26188 14297 26222 14331
rect 27160 14297 27194 14331
rect 29745 14297 29779 14331
rect 38209 14297 38243 14331
rect 39037 14297 39071 14331
rect 40325 14297 40359 14331
rect 4997 14229 5031 14263
rect 5825 14229 5859 14263
rect 7481 14229 7515 14263
rect 14289 14229 14323 14263
rect 16313 14229 16347 14263
rect 19257 14229 19291 14263
rect 23305 14229 23339 14263
rect 23857 14229 23891 14263
rect 28273 14229 28307 14263
rect 29929 14229 29963 14263
rect 34161 14229 34195 14263
rect 38577 14229 38611 14263
rect 40417 14229 40451 14263
rect 8493 14025 8527 14059
rect 13185 14025 13219 14059
rect 21281 14025 21315 14059
rect 23397 14025 23431 14059
rect 25605 14025 25639 14059
rect 27169 14025 27203 14059
rect 34529 14025 34563 14059
rect 7380 13957 7414 13991
rect 18337 13957 18371 13991
rect 18889 13957 18923 13991
rect 19625 13957 19659 13991
rect 20545 13957 20579 13991
rect 22569 13957 22603 13991
rect 22661 13957 22695 13991
rect 28273 13957 28307 13991
rect 28457 13957 28491 13991
rect 28641 13957 28675 13991
rect 36553 13957 36587 13991
rect 37657 13957 37691 13991
rect 10618 13889 10652 13923
rect 10885 13889 10919 13923
rect 11989 13889 12023 13923
rect 12173 13889 12207 13923
rect 14298 13889 14332 13923
rect 14565 13889 14599 13923
rect 21833 13889 21867 13923
rect 22385 13889 22419 13923
rect 22753 13889 22787 13923
rect 23581 13889 23615 13923
rect 23857 13889 23891 13923
rect 24317 13889 24351 13923
rect 27425 13889 27459 13923
rect 27518 13889 27552 13923
rect 27629 13889 27663 13923
rect 27813 13889 27847 13923
rect 29101 13889 29135 13923
rect 29653 13889 29687 13923
rect 29837 13889 29871 13923
rect 29929 13889 29963 13923
rect 30021 13889 30055 13923
rect 35633 13889 35667 13923
rect 36737 13889 36771 13923
rect 5549 13821 5583 13855
rect 7113 13821 7147 13855
rect 20729 13821 20763 13855
rect 23765 13821 23799 13855
rect 30297 13821 30331 13855
rect 35909 13821 35943 13855
rect 9505 13685 9539 13719
rect 22937 13685 22971 13719
rect 23581 13685 23615 13719
rect 36369 13685 36403 13719
rect 38945 13685 38979 13719
rect 2329 13481 2363 13515
rect 4537 13481 4571 13515
rect 9965 13481 9999 13515
rect 10517 13481 10551 13515
rect 18613 13481 18647 13515
rect 20545 13481 20579 13515
rect 23213 13481 23247 13515
rect 24869 13481 24903 13515
rect 25973 13481 26007 13515
rect 37657 13481 37691 13515
rect 23029 13413 23063 13447
rect 24501 13413 24535 13447
rect 26985 13413 27019 13447
rect 29653 13413 29687 13447
rect 6837 13345 6871 13379
rect 9505 13345 9539 13379
rect 9597 13345 9631 13379
rect 28181 13345 28215 13379
rect 34161 13345 34195 13379
rect 35725 13345 35759 13379
rect 2513 13277 2547 13311
rect 6745 13277 6779 13311
rect 9229 13277 9263 13311
rect 9413 13277 9447 13311
rect 9781 13277 9815 13311
rect 14289 13277 14323 13311
rect 23213 13277 23247 13311
rect 23305 13277 23339 13311
rect 24685 13277 24719 13311
rect 24777 13277 24811 13311
rect 24961 13277 24995 13311
rect 27241 13277 27275 13311
rect 27350 13277 27384 13311
rect 27445 13274 27479 13308
rect 27629 13277 27663 13311
rect 31033 13277 31067 13311
rect 35081 13277 35115 13311
rect 35265 13277 35299 13311
rect 38393 13277 38427 13311
rect 38577 13277 38611 13311
rect 38669 13277 38703 13311
rect 38761 13277 38795 13311
rect 39865 13277 39899 13311
rect 58173 13277 58207 13311
rect 14105 13209 14139 13243
rect 17693 13209 17727 13243
rect 17877 13209 17911 13243
rect 19809 13209 19843 13243
rect 19993 13209 20027 13243
rect 21373 13209 21407 13243
rect 23489 13209 23523 13243
rect 30766 13209 30800 13243
rect 31953 13209 31987 13243
rect 32137 13209 32171 13243
rect 33894 13209 33928 13243
rect 35970 13209 36004 13243
rect 6377 13141 6411 13175
rect 7021 13141 7055 13175
rect 7481 13141 7515 13175
rect 14473 13141 14507 13175
rect 18061 13141 18095 13175
rect 26433 13141 26467 13175
rect 32321 13141 32355 13175
rect 32781 13141 32815 13175
rect 35265 13141 35299 13175
rect 37105 13141 37139 13175
rect 39037 13141 39071 13175
rect 4629 12937 4663 12971
rect 5089 12937 5123 12971
rect 14197 12937 14231 12971
rect 17049 12937 17083 12971
rect 25329 12937 25363 12971
rect 27813 12937 27847 12971
rect 29653 12937 29687 12971
rect 32965 12937 32999 12971
rect 34989 12937 35023 12971
rect 35633 12937 35667 12971
rect 39957 12937 39991 12971
rect 11529 12869 11563 12903
rect 15393 12869 15427 12903
rect 21005 12869 21039 12903
rect 24869 12869 24903 12903
rect 30297 12869 30331 12903
rect 30481 12869 30515 12903
rect 31493 12869 31527 12903
rect 38844 12869 38878 12903
rect 2145 12801 2179 12835
rect 3056 12801 3090 12835
rect 4997 12801 5031 12835
rect 6653 12801 6687 12835
rect 6837 12801 6871 12835
rect 6929 12801 6963 12835
rect 7205 12801 7239 12835
rect 8401 12801 8435 12835
rect 10241 12801 10275 12835
rect 10425 12801 10459 12835
rect 10793 12801 10827 12835
rect 14473 12801 14507 12835
rect 14565 12801 14599 12835
rect 14657 12801 14691 12835
rect 14841 12801 14875 12835
rect 18162 12801 18196 12835
rect 18429 12801 18463 12835
rect 19165 12801 19199 12835
rect 19257 12801 19291 12835
rect 19349 12801 19383 12835
rect 19545 12801 19579 12835
rect 20361 12801 20395 12835
rect 20821 12801 20855 12835
rect 22109 12801 22143 12835
rect 24133 12801 24167 12835
rect 24685 12801 24719 12835
rect 32309 12801 32343 12835
rect 32505 12801 32539 12835
rect 32600 12801 32634 12835
rect 32689 12801 32723 12835
rect 35909 12801 35943 12835
rect 36001 12801 36035 12835
rect 36093 12801 36127 12835
rect 36277 12801 36311 12835
rect 38577 12801 38611 12835
rect 1961 12733 1995 12767
rect 2789 12733 2823 12767
rect 5273 12733 5307 12767
rect 7021 12733 7055 12767
rect 8677 12733 8711 12767
rect 10517 12733 10551 12767
rect 10609 12733 10643 12767
rect 23857 12733 23891 12767
rect 20177 12665 20211 12699
rect 2329 12597 2363 12631
rect 4169 12597 4203 12631
rect 7389 12597 7423 12631
rect 10977 12597 11011 12631
rect 18889 12597 18923 12631
rect 21189 12597 21223 12631
rect 27077 12597 27111 12631
rect 7941 12393 7975 12427
rect 19257 12393 19291 12427
rect 22661 12393 22695 12427
rect 23673 12393 23707 12427
rect 24961 12393 24995 12427
rect 30757 12393 30791 12427
rect 12173 12325 12207 12359
rect 28181 12325 28215 12359
rect 5365 12257 5399 12291
rect 20821 12257 20855 12291
rect 21097 12257 21131 12291
rect 38209 12257 38243 12291
rect 2513 12189 2547 12223
rect 10793 12189 10827 12223
rect 11060 12189 11094 12223
rect 13553 12189 13587 12223
rect 14657 12189 14691 12223
rect 14749 12189 14783 12223
rect 14841 12189 14875 12223
rect 15025 12189 15059 12223
rect 18429 12189 18463 12223
rect 19625 12189 19659 12223
rect 21833 12189 21867 12223
rect 21922 12189 21956 12223
rect 22017 12189 22051 12223
rect 22201 12189 22235 12223
rect 25513 12189 25547 12223
rect 31309 12189 31343 12223
rect 31493 12189 31527 12223
rect 31604 12189 31638 12223
rect 31697 12189 31731 12223
rect 33793 12189 33827 12223
rect 37933 12189 37967 12223
rect 5181 12121 5215 12155
rect 6653 12121 6687 12155
rect 8953 12121 8987 12155
rect 13369 12121 13403 12155
rect 18184 12121 18218 12155
rect 19441 12121 19475 12155
rect 25758 12121 25792 12155
rect 27629 12121 27663 12155
rect 28365 12121 28399 12155
rect 31953 12121 31987 12155
rect 33526 12121 33560 12155
rect 2697 12053 2731 12087
rect 4353 12053 4387 12087
rect 4813 12053 4847 12087
rect 5273 12053 5307 12087
rect 13185 12053 13219 12087
rect 14381 12053 14415 12087
rect 15485 12053 15519 12087
rect 17049 12053 17083 12087
rect 21557 12053 21591 12087
rect 24501 12053 24535 12087
rect 26893 12053 26927 12087
rect 27537 12053 27571 12087
rect 32413 12053 32447 12087
rect 35449 12053 35483 12087
rect 4261 11849 4295 11883
rect 14013 11849 14047 11883
rect 18061 11849 18095 11883
rect 19901 11849 19935 11883
rect 25605 11849 25639 11883
rect 32505 11849 32539 11883
rect 35173 11849 35207 11883
rect 38209 11849 38243 11883
rect 3126 11781 3160 11815
rect 13645 11781 13679 11815
rect 17509 11781 17543 11815
rect 21036 11781 21070 11815
rect 35449 11781 35483 11815
rect 36277 11781 36311 11815
rect 36461 11781 36495 11815
rect 2881 11713 2915 11747
rect 4905 11713 4939 11747
rect 6653 11713 6687 11747
rect 8778 11713 8812 11747
rect 9045 11713 9079 11747
rect 11805 11713 11839 11747
rect 13829 11713 13863 11747
rect 14749 11713 14783 11747
rect 14841 11713 14875 11747
rect 14933 11716 14967 11750
rect 15117 11713 15151 11747
rect 18291 11713 18325 11747
rect 18429 11713 18463 11747
rect 18521 11713 18555 11747
rect 18705 11713 18739 11747
rect 19165 11713 19199 11747
rect 22477 11713 22511 11747
rect 22569 11713 22603 11747
rect 22661 11713 22695 11747
rect 22845 11713 22879 11747
rect 23397 11713 23431 11747
rect 25881 11713 25915 11747
rect 25973 11713 26007 11747
rect 26065 11713 26099 11747
rect 26249 11713 26283 11747
rect 28181 11713 28215 11747
rect 32137 11713 32171 11747
rect 32321 11713 32355 11747
rect 33057 11713 33091 11747
rect 33333 11713 33367 11747
rect 35357 11713 35391 11747
rect 35541 11713 35575 11747
rect 35725 11713 35759 11747
rect 38761 11713 38795 11747
rect 5089 11645 5123 11679
rect 6377 11645 6411 11679
rect 11529 11645 11563 11679
rect 21281 11645 21315 11679
rect 39037 11645 39071 11679
rect 15577 11577 15611 11611
rect 25053 11577 25087 11611
rect 58173 11577 58207 11611
rect 4721 11509 4755 11543
rect 7665 11509 7699 11543
rect 14473 11509 14507 11543
rect 19349 11509 19383 11543
rect 22201 11509 22235 11543
rect 28365 11509 28399 11543
rect 34713 11509 34747 11543
rect 3801 11305 3835 11339
rect 12449 11305 12483 11339
rect 14197 11305 14231 11339
rect 18521 11305 18555 11339
rect 21097 11305 21131 11339
rect 26157 11305 26191 11339
rect 29929 11305 29963 11339
rect 32965 11305 32999 11339
rect 34713 11305 34747 11339
rect 16037 11237 16071 11271
rect 17049 11237 17083 11271
rect 3249 11169 3283 11203
rect 5641 11169 5675 11203
rect 5733 11169 5767 11203
rect 6745 11169 6779 11203
rect 6843 11169 6877 11203
rect 7849 11169 7883 11203
rect 21649 11169 21683 11203
rect 23581 11169 23615 11203
rect 28181 11169 28215 11203
rect 28457 11169 28491 11203
rect 36369 11169 36403 11203
rect 38209 11169 38243 11203
rect 2973 11101 3007 11135
rect 3985 11101 4019 11135
rect 6561 11101 6595 11135
rect 6925 11099 6959 11133
rect 7113 11101 7147 11135
rect 7573 11101 7607 11135
rect 9137 11101 9171 11135
rect 11529 11101 11563 11135
rect 12265 11101 12299 11135
rect 15310 11101 15344 11135
rect 15577 11101 15611 11135
rect 23489 11101 23523 11135
rect 23673 11101 23707 11135
rect 25973 11101 26007 11135
rect 30665 11101 30699 11135
rect 30757 11101 30791 11135
rect 30849 11101 30883 11135
rect 31033 11101 31067 11135
rect 32045 11101 32079 11135
rect 32321 11101 32355 11135
rect 35541 11101 35575 11135
rect 35633 11101 35667 11135
rect 35725 11101 35759 11135
rect 35909 11101 35943 11135
rect 36553 11101 36587 11135
rect 38669 11101 38703 11135
rect 38853 11101 38887 11135
rect 38945 11101 38979 11135
rect 39037 11101 39071 11135
rect 39865 11101 39899 11135
rect 5273 11033 5307 11067
rect 5917 11033 5951 11067
rect 16221 11033 16255 11067
rect 16865 11033 16899 11067
rect 17785 11033 17819 11067
rect 18429 11033 18463 11067
rect 20453 11033 20487 11067
rect 21005 11033 21039 11067
rect 21916 11033 21950 11067
rect 25789 11033 25823 11067
rect 30389 11033 30423 11067
rect 36737 11033 36771 11067
rect 37841 11033 37875 11067
rect 38025 11033 38059 11067
rect 39313 11033 39347 11067
rect 6377 10965 6411 10999
rect 8953 10965 8987 10999
rect 11713 10965 11747 10999
rect 19717 10965 19751 10999
rect 23029 10965 23063 10999
rect 35265 10965 35299 10999
rect 4353 10761 4387 10795
rect 7021 10761 7055 10795
rect 7849 10761 7883 10795
rect 14013 10761 14047 10795
rect 22753 10761 22787 10795
rect 28273 10761 28307 10795
rect 31033 10761 31067 10795
rect 36461 10761 36495 10795
rect 41245 10761 41279 10795
rect 8576 10693 8610 10727
rect 15126 10693 15160 10727
rect 22569 10693 22603 10727
rect 29837 10693 29871 10727
rect 30665 10693 30699 10727
rect 37657 10693 37691 10727
rect 40132 10693 40166 10727
rect 2237 10625 2271 10659
rect 4445 10625 4479 10659
rect 7665 10625 7699 10659
rect 8309 10625 8343 10659
rect 22385 10625 22419 10659
rect 24593 10625 24627 10659
rect 25053 10625 25087 10659
rect 25320 10625 25354 10659
rect 28089 10625 28123 10659
rect 29009 10625 29043 10659
rect 29114 10628 29148 10662
rect 29214 10625 29248 10659
rect 29377 10625 29411 10659
rect 30849 10625 30883 10659
rect 35081 10625 35115 10659
rect 35348 10625 35382 10659
rect 7481 10557 7515 10591
rect 15393 10557 15427 10591
rect 24317 10557 24351 10591
rect 39865 10557 39899 10591
rect 2421 10421 2455 10455
rect 9689 10421 9723 10455
rect 10241 10421 10275 10455
rect 12449 10421 12483 10455
rect 13001 10421 13035 10455
rect 18981 10421 19015 10455
rect 19625 10421 19659 10455
rect 26433 10421 26467 10455
rect 28733 10421 28767 10455
rect 38945 10421 38979 10455
rect 58173 10421 58207 10455
rect 2053 10217 2087 10251
rect 7021 10217 7055 10251
rect 8953 10217 8987 10251
rect 21281 10217 21315 10251
rect 22201 10217 22235 10251
rect 25421 10217 25455 10251
rect 26433 10217 26467 10251
rect 27997 10217 28031 10251
rect 29561 10217 29595 10251
rect 30665 10217 30699 10251
rect 32505 10217 32539 10251
rect 36829 10217 36863 10251
rect 37473 10217 37507 10251
rect 2513 10149 2547 10183
rect 23857 10149 23891 10183
rect 29009 10149 29043 10183
rect 3157 10081 3191 10115
rect 5181 10081 5215 10115
rect 9597 10081 9631 10115
rect 10425 10081 10459 10115
rect 13185 10081 13219 10115
rect 21833 10081 21867 10115
rect 1777 10013 1811 10047
rect 1869 10013 1903 10047
rect 6929 10013 6963 10047
rect 9321 10013 9355 10047
rect 12173 10013 12207 10047
rect 22017 10013 22051 10047
rect 24777 10013 24811 10047
rect 24961 10013 24995 10047
rect 25053 10013 25087 10047
rect 25145 10013 25179 10047
rect 25881 10013 25915 10047
rect 26157 10013 26191 10047
rect 26249 10013 26283 10047
rect 27445 10013 27479 10047
rect 27629 10013 27663 10047
rect 27813 10013 27847 10047
rect 28457 10013 28491 10047
rect 28641 10013 28675 10047
rect 28825 10013 28859 10047
rect 31217 10013 31251 10047
rect 37933 10013 37967 10047
rect 38117 10013 38151 10047
rect 38209 10013 38243 10047
rect 38301 10013 38335 10047
rect 2881 9945 2915 9979
rect 4997 9945 5031 9979
rect 13001 9945 13035 9979
rect 26065 9945 26099 9979
rect 27721 9945 27755 9979
rect 28733 9945 28767 9979
rect 29745 9945 29779 9979
rect 29929 9945 29963 9979
rect 39037 9945 39071 9979
rect 2973 9877 3007 9911
rect 3893 9877 3927 9911
rect 9413 9877 9447 9911
rect 12633 9877 12667 9911
rect 13093 9877 13127 9911
rect 38577 9877 38611 9911
rect 15117 9673 15151 9707
rect 25145 9673 25179 9707
rect 29653 9673 29687 9707
rect 31585 9673 31619 9707
rect 37841 9673 37875 9707
rect 2320 9605 2354 9639
rect 10241 9605 10275 9639
rect 20729 9605 20763 9639
rect 22661 9605 22695 9639
rect 25329 9605 25363 9639
rect 33241 9605 33275 9639
rect 5549 9537 5583 9571
rect 11989 9537 12023 9571
rect 12633 9537 12667 9571
rect 12817 9537 12851 9571
rect 14933 9537 14967 9571
rect 17325 9537 17359 9571
rect 22385 9537 22419 9571
rect 22569 9537 22603 9571
rect 22753 9537 22787 9571
rect 24501 9537 24535 9571
rect 25513 9537 25547 9571
rect 28273 9537 28307 9571
rect 28540 9537 28574 9571
rect 30205 9537 30239 9571
rect 30472 9537 30506 9571
rect 32137 9537 32171 9571
rect 32321 9537 32355 9571
rect 32413 9537 32447 9571
rect 32505 9537 32539 9571
rect 35265 9537 35299 9571
rect 35449 9537 35483 9571
rect 37473 9537 37507 9571
rect 37657 9537 37691 9571
rect 39414 9537 39448 9571
rect 39681 9537 39715 9571
rect 2053 9469 2087 9503
rect 5825 9469 5859 9503
rect 10425 9469 10459 9503
rect 10517 9469 10551 9503
rect 10885 9469 10919 9503
rect 11529 9469 11563 9503
rect 11897 9469 11931 9503
rect 14473 9469 14507 9503
rect 19073 9469 19107 9503
rect 16773 9401 16807 9435
rect 22937 9401 22971 9435
rect 24685 9401 24719 9435
rect 38301 9401 38335 9435
rect 3433 9333 3467 9367
rect 6377 9333 6411 9367
rect 12173 9333 12207 9367
rect 13001 9333 13035 9367
rect 15669 9333 15703 9367
rect 32781 9333 32815 9367
rect 35633 9333 35667 9367
rect 5273 9129 5307 9163
rect 14105 9129 14139 9163
rect 20637 9129 20671 9163
rect 23397 9129 23431 9163
rect 31217 9129 31251 9163
rect 33241 9129 33275 9163
rect 36093 9129 36127 9163
rect 37933 9129 37967 9163
rect 9597 9061 9631 9095
rect 32229 9061 32263 9095
rect 4997 8993 5031 9027
rect 5825 8993 5859 9027
rect 11713 8993 11747 9027
rect 21189 8993 21223 9027
rect 22017 8993 22051 9027
rect 22293 8993 22327 9027
rect 28181 8993 28215 9027
rect 28457 8993 28491 9027
rect 39313 8993 39347 9027
rect 5089 8925 5123 8959
rect 6653 8925 6687 8959
rect 11437 8925 11471 8959
rect 11621 8925 11655 8959
rect 11805 8925 11839 8959
rect 11989 8925 12023 8959
rect 13093 8925 13127 8959
rect 15485 8925 15519 8959
rect 17325 8925 17359 8959
rect 19257 8925 19291 8959
rect 21097 8925 21131 8959
rect 21281 8925 21315 8959
rect 30849 8925 30883 8959
rect 31677 8925 31711 8959
rect 31953 8925 31987 8959
rect 32045 8925 32079 8959
rect 32689 8925 32723 8959
rect 32965 8925 32999 8959
rect 33057 8925 33091 8959
rect 34713 8925 34747 8959
rect 36829 8925 36863 8959
rect 37013 8925 37047 8959
rect 37105 8925 37139 8959
rect 37197 8925 37231 8959
rect 58173 8925 58207 8959
rect 4629 8857 4663 8891
rect 6469 8857 6503 8891
rect 9413 8857 9447 8891
rect 15218 8857 15252 8891
rect 17592 8857 17626 8891
rect 19502 8857 19536 8891
rect 31033 8857 31067 8891
rect 31861 8857 31895 8891
rect 32873 8857 32907 8891
rect 34980 8857 35014 8891
rect 37473 8857 37507 8891
rect 39046 8857 39080 8891
rect 3249 8789 3283 8823
rect 4169 8789 4203 8823
rect 7205 8789 7239 8823
rect 7757 8789 7791 8823
rect 10057 8789 10091 8823
rect 11253 8789 11287 8823
rect 13277 8789 13311 8823
rect 16313 8789 16347 8823
rect 16865 8789 16899 8823
rect 18705 8789 18739 8823
rect 8769 8585 8803 8619
rect 9689 8585 9723 8619
rect 10149 8585 10183 8619
rect 13461 8585 13495 8619
rect 14197 8585 14231 8619
rect 17509 8585 17543 8619
rect 18705 8585 18739 8619
rect 21005 8585 21039 8619
rect 29837 8585 29871 8619
rect 32689 8585 32723 8619
rect 34529 8585 34563 8619
rect 34989 8585 35023 8619
rect 37289 8585 37323 8619
rect 19349 8517 19383 8551
rect 20177 8517 20211 8551
rect 29469 8517 29503 8551
rect 29561 8517 29595 8551
rect 32321 8517 32355 8551
rect 32413 8517 32447 8551
rect 37473 8517 37507 8551
rect 6653 8449 6687 8483
rect 11713 8449 11747 8483
rect 11897 8449 11931 8483
rect 12081 8449 12115 8483
rect 12265 8449 12299 8483
rect 14013 8449 14047 8483
rect 14749 8449 14783 8483
rect 15016 8449 15050 8483
rect 16957 8449 16991 8483
rect 18061 8449 18095 8483
rect 18245 8449 18279 8483
rect 18337 8449 18371 8483
rect 18429 8449 18463 8483
rect 19533 8449 19567 8483
rect 20361 8449 20395 8483
rect 21833 8449 21867 8483
rect 22109 8449 22143 8483
rect 23673 8449 23707 8483
rect 23765 8449 23799 8483
rect 23857 8449 23891 8483
rect 24041 8449 24075 8483
rect 27997 8449 28031 8483
rect 28273 8449 28307 8483
rect 29285 8449 29319 8483
rect 29653 8449 29687 8483
rect 32137 8449 32171 8483
rect 32505 8449 32539 8483
rect 35265 8449 35299 8483
rect 35357 8449 35391 8483
rect 35449 8449 35483 8483
rect 35633 8449 35667 8483
rect 36737 8449 36771 8483
rect 37657 8449 37691 8483
rect 5825 8381 5859 8415
rect 6377 8381 6411 8415
rect 8585 8381 8619 8415
rect 8953 8381 8987 8415
rect 11989 8381 12023 8415
rect 12817 8381 12851 8415
rect 19165 8381 19199 8415
rect 1593 8313 1627 8347
rect 2145 8313 2179 8347
rect 2697 8313 2731 8347
rect 4261 8313 4295 8347
rect 7665 8313 7699 8347
rect 10701 8313 10735 8347
rect 11529 8313 11563 8347
rect 16129 8313 16163 8347
rect 19993 8313 20027 8347
rect 3433 8245 3467 8279
rect 5595 8245 5629 8279
rect 8953 8245 8987 8279
rect 23397 8245 23431 8279
rect 10793 8041 10827 8075
rect 14289 8041 14323 8075
rect 17141 8041 17175 8075
rect 17693 8041 17727 8075
rect 19441 8041 19475 8075
rect 27997 8041 28031 8075
rect 7297 7973 7331 8007
rect 13553 7973 13587 8007
rect 20637 7973 20671 8007
rect 26249 7973 26283 8007
rect 35081 7973 35115 8007
rect 3157 7905 3191 7939
rect 5089 7905 5123 7939
rect 8125 7905 8159 7939
rect 8401 7905 8435 7939
rect 9413 7905 9447 7939
rect 10609 7905 10643 7939
rect 13001 7905 13035 7939
rect 2881 7837 2915 7871
rect 4905 7837 4939 7871
rect 5181 7837 5215 7871
rect 5273 7837 5307 7871
rect 5457 7837 5491 7871
rect 5917 7837 5951 7871
rect 8217 7837 8251 7871
rect 9137 7837 9171 7871
rect 9275 7837 9309 7871
rect 9505 7837 9539 7871
rect 9689 7837 9723 7871
rect 10517 7837 10551 7871
rect 11897 7837 11931 7871
rect 14105 7837 14139 7871
rect 14841 7837 14875 7871
rect 17969 7837 18003 7871
rect 18061 7837 18095 7871
rect 18153 7837 18187 7871
rect 18337 7837 18371 7871
rect 19257 7837 19291 7871
rect 21189 7837 21223 7871
rect 21373 7837 21407 7871
rect 23049 7837 23083 7871
rect 23305 7837 23339 7871
rect 24869 7837 24903 7871
rect 27445 7837 27479 7871
rect 27721 7837 27755 7871
rect 27813 7837 27847 7871
rect 30849 7837 30883 7871
rect 35265 7837 35299 7871
rect 35449 7837 35483 7871
rect 35633 7837 35667 7871
rect 58173 7837 58207 7871
rect 2053 7769 2087 7803
rect 6162 7769 6196 7803
rect 7757 7769 7791 7803
rect 12449 7769 12483 7803
rect 25136 7769 25170 7803
rect 27629 7769 27663 7803
rect 31033 7769 31067 7803
rect 35357 7769 35391 7803
rect 1501 7701 1535 7735
rect 2513 7701 2547 7735
rect 2973 7701 3007 7735
rect 3985 7701 4019 7735
rect 4721 7701 4755 7735
rect 8953 7701 8987 7735
rect 10149 7701 10183 7735
rect 11345 7701 11379 7735
rect 15025 7701 15059 7735
rect 15577 7701 15611 7735
rect 16681 7701 16715 7735
rect 21281 7701 21315 7735
rect 21925 7701 21959 7735
rect 26893 7701 26927 7735
rect 30665 7701 30699 7735
rect 3065 7497 3099 7531
rect 3525 7497 3559 7531
rect 5181 7497 5215 7531
rect 7941 7497 7975 7531
rect 10885 7497 10919 7531
rect 14473 7497 14507 7531
rect 15025 7497 15059 7531
rect 17601 7497 17635 7531
rect 22845 7497 22879 7531
rect 23305 7497 23339 7531
rect 31585 7497 31619 7531
rect 35081 7497 35115 7531
rect 36369 7497 36403 7531
rect 38025 7497 38059 7531
rect 3433 7429 3467 7463
rect 4537 7429 4571 7463
rect 12734 7429 12768 7463
rect 16681 7429 16715 7463
rect 16865 7429 16899 7463
rect 22569 7429 22603 7463
rect 23489 7429 23523 7463
rect 23673 7429 23707 7463
rect 26157 7429 26191 7463
rect 34437 7429 34471 7463
rect 35449 7429 35483 7463
rect 2237 7361 2271 7395
rect 2421 7361 2455 7395
rect 4905 7361 4939 7395
rect 4997 7361 5031 7395
rect 6837 7361 6871 7395
rect 7849 7361 7883 7395
rect 14289 7361 14323 7395
rect 15301 7361 15335 7395
rect 15393 7361 15427 7395
rect 15485 7361 15519 7395
rect 15669 7361 15703 7395
rect 17049 7361 17083 7395
rect 18889 7361 18923 7395
rect 21097 7361 21131 7395
rect 21281 7361 21315 7395
rect 22293 7361 22327 7395
rect 22477 7361 22511 7395
rect 22661 7361 22695 7395
rect 24685 7361 24719 7395
rect 24869 7361 24903 7395
rect 24961 7361 24995 7395
rect 25053 7361 25087 7395
rect 25789 7361 25823 7395
rect 25973 7361 26007 7395
rect 27629 7361 27663 7395
rect 27718 7361 27752 7395
rect 27818 7361 27852 7395
rect 27997 7361 28031 7395
rect 28457 7361 28491 7395
rect 30472 7361 30506 7395
rect 34621 7361 34655 7395
rect 35265 7361 35299 7395
rect 35357 7361 35391 7395
rect 35633 7361 35667 7395
rect 38577 7361 38611 7395
rect 38761 7361 38795 7395
rect 3709 7293 3743 7327
rect 7021 7293 7055 7327
rect 8125 7293 8159 7327
rect 13001 7293 13035 7327
rect 20361 7293 20395 7327
rect 20913 7293 20947 7327
rect 25329 7293 25363 7327
rect 30205 7293 30239 7327
rect 1777 7225 1811 7259
rect 7481 7225 7515 7259
rect 18705 7225 18739 7259
rect 24133 7225 24167 7259
rect 34253 7225 34287 7259
rect 2605 7157 2639 7191
rect 5733 7157 5767 7191
rect 6653 7157 6687 7191
rect 8677 7157 8711 7191
rect 9229 7157 9263 7191
rect 9781 7157 9815 7191
rect 10425 7157 10459 7191
rect 11621 7157 11655 7191
rect 13829 7157 13863 7191
rect 18153 7157 18187 7191
rect 19349 7157 19383 7191
rect 27353 7157 27387 7191
rect 28641 7157 28675 7191
rect 38945 7157 38979 7191
rect 6009 6953 6043 6987
rect 3893 6817 3927 6851
rect 11897 6817 11931 6851
rect 14289 6817 14323 6851
rect 18705 6817 18739 6851
rect 25973 6817 26007 6851
rect 39865 6817 39899 6851
rect 2237 6749 2271 6783
rect 2329 6749 2363 6783
rect 3157 6749 3191 6783
rect 6193 6749 6227 6783
rect 6653 6749 6687 6783
rect 7481 6749 7515 6783
rect 7941 6749 7975 6783
rect 9137 6749 9171 6783
rect 11630 6749 11664 6783
rect 12633 6749 12667 6783
rect 15945 6749 15979 6783
rect 18429 6749 18463 6783
rect 21833 6749 21867 6783
rect 22155 6749 22189 6783
rect 23489 6749 23523 6783
rect 23581 6749 23615 6783
rect 23673 6749 23707 6783
rect 23857 6749 23891 6783
rect 24685 6749 24719 6783
rect 24777 6749 24811 6783
rect 24869 6749 24903 6783
rect 25053 6749 25087 6783
rect 26249 6749 26283 6783
rect 27261 6749 27295 6783
rect 30021 6749 30055 6783
rect 32413 6749 32447 6783
rect 32680 6749 32714 6783
rect 35357 6749 35391 6783
rect 35449 6749 35483 6783
rect 35541 6749 35575 6783
rect 35725 6749 35759 6783
rect 36645 6749 36679 6783
rect 36829 6749 36863 6783
rect 36921 6749 36955 6783
rect 37013 6749 37047 6783
rect 37749 6749 37783 6783
rect 38669 6749 38703 6783
rect 38761 6749 38795 6783
rect 38853 6749 38887 6783
rect 39037 6749 39071 6783
rect 1685 6681 1719 6715
rect 4445 6681 4479 6715
rect 10057 6681 10091 6715
rect 13553 6681 13587 6715
rect 15761 6681 15795 6715
rect 21005 6681 21039 6715
rect 27506 6681 27540 6715
rect 2513 6613 2547 6647
rect 2973 6613 3007 6647
rect 4997 6613 5031 6647
rect 5549 6613 5583 6647
rect 6837 6613 6871 6647
rect 7297 6613 7331 6647
rect 8125 6613 8159 6647
rect 8953 6613 8987 6647
rect 10517 6613 10551 6647
rect 14841 6613 14875 6647
rect 15577 6613 15611 6647
rect 16589 6613 16623 6647
rect 17417 6613 17451 6647
rect 19257 6613 19291 6647
rect 19993 6613 20027 6647
rect 20453 6613 20487 6647
rect 23213 6613 23247 6647
rect 24409 6613 24443 6647
rect 28641 6613 28675 6647
rect 31309 6613 31343 6647
rect 33793 6613 33827 6647
rect 35081 6613 35115 6647
rect 37289 6613 37323 6647
rect 38393 6613 38427 6647
rect 3709 6409 3743 6443
rect 23673 6409 23707 6443
rect 28273 6409 28307 6443
rect 29653 6409 29687 6443
rect 30205 6409 30239 6443
rect 32229 6409 32263 6443
rect 36001 6409 36035 6443
rect 37289 6409 37323 6443
rect 39681 6409 39715 6443
rect 2596 6341 2630 6375
rect 13921 6341 13955 6375
rect 14381 6341 14415 6375
rect 18797 6341 18831 6375
rect 19257 6341 19291 6375
rect 19441 6341 19475 6375
rect 23397 6341 23431 6375
rect 25973 6341 26007 6375
rect 34345 6341 34379 6375
rect 37473 6341 37507 6375
rect 37657 6341 37691 6375
rect 38546 6341 38580 6375
rect 4905 6273 4939 6307
rect 5089 6273 5123 6307
rect 5825 6273 5859 6307
rect 6653 6273 6687 6307
rect 7665 6273 7699 6307
rect 8953 6273 8987 6307
rect 9209 6273 9243 6307
rect 16957 6273 16991 6307
rect 18613 6273 18647 6307
rect 23121 6273 23155 6307
rect 23305 6273 23339 6307
rect 23489 6273 23523 6307
rect 27261 6273 27295 6307
rect 28457 6273 28491 6307
rect 28641 6273 28675 6307
rect 30435 6273 30469 6307
rect 30573 6273 30607 6307
rect 30665 6273 30699 6307
rect 30849 6273 30883 6307
rect 35173 6273 35207 6307
rect 35262 6273 35296 6307
rect 35357 6273 35391 6307
rect 35541 6273 35575 6307
rect 36185 6273 36219 6307
rect 36369 6273 36403 6307
rect 2329 6205 2363 6239
rect 4445 6205 4479 6239
rect 6929 6205 6963 6239
rect 16037 6205 16071 6239
rect 16681 6205 16715 6239
rect 21833 6205 21867 6239
rect 22155 6205 22189 6239
rect 26985 6205 27019 6239
rect 38301 6205 38335 6239
rect 6745 6137 6779 6171
rect 7849 6137 7883 6171
rect 10333 6137 10367 6171
rect 11805 6137 11839 6171
rect 58173 6137 58207 6171
rect 1869 6069 1903 6103
rect 5089 6069 5123 6103
rect 5641 6069 5675 6103
rect 6653 6069 6687 6103
rect 8493 6069 8527 6103
rect 10793 6069 10827 6103
rect 12265 6069 12299 6103
rect 13277 6069 13311 6103
rect 18429 6069 18463 6103
rect 19625 6069 19659 6103
rect 20177 6069 20211 6103
rect 20637 6069 20671 6103
rect 21189 6069 21223 6103
rect 24685 6069 24719 6103
rect 33793 6069 33827 6103
rect 34897 6069 34931 6103
rect 4629 5865 4663 5899
rect 7757 5865 7791 5899
rect 15669 5865 15703 5899
rect 20637 5865 20671 5899
rect 24961 5865 24995 5899
rect 26157 5865 26191 5899
rect 26893 5865 26927 5899
rect 31401 5865 31435 5899
rect 36553 5865 36587 5899
rect 13461 5797 13495 5831
rect 23121 5797 23155 5831
rect 24501 5797 24535 5831
rect 32597 5797 32631 5831
rect 34713 5797 34747 5831
rect 9137 5729 9171 5763
rect 17417 5729 17451 5763
rect 19257 5729 19291 5763
rect 2237 5661 2271 5695
rect 5917 5661 5951 5695
rect 6929 5661 6963 5695
rect 7021 5661 7055 5695
rect 7573 5661 7607 5695
rect 9781 5661 9815 5695
rect 10425 5661 10459 5695
rect 11069 5661 11103 5695
rect 11713 5661 11747 5695
rect 12357 5661 12391 5695
rect 12817 5661 12851 5695
rect 14289 5661 14323 5695
rect 16405 5661 16439 5695
rect 16497 5661 16531 5695
rect 16589 5661 16623 5695
rect 16773 5661 16807 5695
rect 17969 5661 18003 5695
rect 18153 5661 18187 5695
rect 18245 5661 18279 5695
rect 18337 5661 18371 5695
rect 22569 5661 22603 5695
rect 22753 5661 22787 5695
rect 22937 5661 22971 5695
rect 25145 5661 25179 5695
rect 25329 5661 25363 5695
rect 28181 5661 28215 5695
rect 30297 5661 30331 5695
rect 30481 5661 30515 5695
rect 30573 5661 30607 5695
rect 30685 5661 30719 5695
rect 31585 5661 31619 5695
rect 32413 5661 32447 5695
rect 35826 5661 35860 5695
rect 36093 5661 36127 5695
rect 3249 5593 3283 5627
rect 8401 5593 8435 5627
rect 14556 5593 14590 5627
rect 18613 5593 18647 5627
rect 19502 5593 19536 5627
rect 22845 5593 22879 5627
rect 28365 5593 28399 5627
rect 31769 5593 31803 5627
rect 32229 5593 32263 5627
rect 37105 5593 37139 5627
rect 1777 5525 1811 5559
rect 2421 5525 2455 5559
rect 6745 5525 6779 5559
rect 16129 5525 16163 5559
rect 21373 5525 21407 5559
rect 21925 5525 21959 5559
rect 23673 5525 23707 5559
rect 27997 5525 28031 5559
rect 29745 5525 29779 5559
rect 30941 5525 30975 5559
rect 38393 5525 38427 5559
rect 3617 5321 3651 5355
rect 6561 5321 6595 5355
rect 9229 5321 9263 5355
rect 12265 5321 12299 5355
rect 14565 5321 14599 5355
rect 16773 5321 16807 5355
rect 24777 5321 24811 5355
rect 38761 5321 38795 5355
rect 1777 5253 1811 5287
rect 6377 5253 6411 5287
rect 7113 5253 7147 5287
rect 8769 5253 8803 5287
rect 17141 5253 17175 5287
rect 24593 5253 24627 5287
rect 37626 5253 37660 5287
rect 2237 5185 2271 5219
rect 2504 5185 2538 5219
rect 4169 5185 4203 5219
rect 4813 5185 4847 5219
rect 5549 5185 5583 5219
rect 7665 5185 7699 5219
rect 8125 5185 8159 5219
rect 9045 5185 9079 5219
rect 11713 5185 11747 5219
rect 12081 5185 12115 5219
rect 14841 5185 14875 5219
rect 14933 5185 14967 5219
rect 15025 5185 15059 5219
rect 15209 5185 15243 5219
rect 16957 5185 16991 5219
rect 18245 5185 18279 5219
rect 18429 5185 18463 5219
rect 18521 5185 18555 5219
rect 18659 5185 18693 5219
rect 24409 5185 24443 5219
rect 27537 5185 27571 5219
rect 27629 5185 27663 5219
rect 27721 5185 27755 5219
rect 27905 5185 27939 5219
rect 30205 5185 30239 5219
rect 30389 5185 30423 5219
rect 30481 5185 30515 5219
rect 30573 5185 30607 5219
rect 37381 5185 37415 5219
rect 6653 5117 6687 5151
rect 7941 5117 7975 5151
rect 8861 5117 8895 5151
rect 11621 5117 11655 5151
rect 23029 5117 23063 5151
rect 29653 5117 29687 5151
rect 54401 5117 54435 5151
rect 7113 5049 7147 5083
rect 8309 5049 8343 5083
rect 10333 5049 10367 5083
rect 23581 5049 23615 5083
rect 55045 5049 55079 5083
rect 4353 4981 4387 5015
rect 4997 4981 5031 5015
rect 5733 4981 5767 5015
rect 8033 4981 8067 5015
rect 8769 4981 8803 5015
rect 10977 4981 11011 5015
rect 12081 4981 12115 5015
rect 13461 4981 13495 5015
rect 14105 4981 14139 5015
rect 15669 4981 15703 5015
rect 17601 4981 17635 5015
rect 18889 4981 18923 5015
rect 19349 4981 19383 5015
rect 20177 4981 20211 5015
rect 21005 4981 21039 5015
rect 21833 4981 21867 5015
rect 22385 4981 22419 5015
rect 26341 4981 26375 5015
rect 27261 4981 27295 5015
rect 30849 4981 30883 5015
rect 53757 4981 53791 5015
rect 58173 4981 58207 5015
rect 1961 4777 1995 4811
rect 6469 4777 6503 4811
rect 7941 4777 7975 4811
rect 8309 4777 8343 4811
rect 9965 4777 9999 4811
rect 10333 4777 10367 4811
rect 10977 4777 11011 4811
rect 12725 4777 12759 4811
rect 20913 4777 20947 4811
rect 25789 4777 25823 4811
rect 28549 4777 28583 4811
rect 32597 4777 32631 4811
rect 4537 4709 4571 4743
rect 5365 4709 5399 4743
rect 11345 4709 11379 4743
rect 11437 4709 11471 4743
rect 15761 4709 15795 4743
rect 18705 4709 18739 4743
rect 52837 4709 52871 4743
rect 55321 4709 55355 4743
rect 8033 4641 8067 4675
rect 9836 4641 9870 4675
rect 10057 4641 10091 4675
rect 11253 4641 11287 4675
rect 19533 4641 19567 4675
rect 27169 4641 27203 4675
rect 31217 4641 31251 4675
rect 54125 4641 54159 4675
rect 55965 4641 55999 4675
rect 2421 4573 2455 4607
rect 3065 4573 3099 4607
rect 3893 4573 3927 4607
rect 5549 4573 5583 4607
rect 6009 4573 6043 4607
rect 6377 4573 6411 4607
rect 6653 4573 6687 4607
rect 7481 4573 7515 4607
rect 7573 4573 7607 4607
rect 9229 4573 9263 4607
rect 11805 4573 11839 4607
rect 12725 4573 12759 4607
rect 12909 4573 12943 4607
rect 13553 4573 13587 4607
rect 14289 4573 14323 4607
rect 15117 4573 15151 4607
rect 16405 4573 16439 4607
rect 16865 4573 16899 4607
rect 18061 4573 18095 4607
rect 19789 4573 19823 4607
rect 21741 4573 21775 4607
rect 22385 4573 22419 4607
rect 23029 4573 23063 4607
rect 23489 4573 23523 4607
rect 24409 4573 24443 4607
rect 27425 4573 27459 4607
rect 31473 4573 31507 4607
rect 52193 4573 52227 4607
rect 53481 4573 53515 4607
rect 4721 4505 4755 4539
rect 9689 4505 9723 4539
rect 24676 4505 24710 4539
rect 2605 4437 2639 4471
rect 3157 4437 3191 4471
rect 4077 4437 4111 4471
rect 6193 4437 6227 4471
rect 9045 4437 9079 4471
rect 14473 4437 14507 4471
rect 3065 4233 3099 4267
rect 5825 4233 5859 4267
rect 6577 4233 6611 4267
rect 6377 4165 6411 4199
rect 25145 4165 25179 4199
rect 1777 4097 1811 4131
rect 2421 4097 2455 4131
rect 3249 4097 3283 4131
rect 4353 4097 4387 4131
rect 4997 4097 5031 4131
rect 5641 4097 5675 4131
rect 7573 4097 7607 4131
rect 9689 4097 9723 4131
rect 10977 4097 11011 4131
rect 14565 4097 14599 4131
rect 15669 4097 15703 4131
rect 17325 4097 17359 4131
rect 22928 4097 22962 4131
rect 35173 4097 35207 4131
rect 35440 4097 35474 4131
rect 54677 4097 54711 4131
rect 4813 4029 4847 4063
rect 5181 4029 5215 4063
rect 7481 4029 7515 4063
rect 8033 4029 8067 4063
rect 8585 4029 8619 4063
rect 8677 4029 8711 4063
rect 10241 4029 10275 4063
rect 11529 4029 11563 4063
rect 12081 4029 12115 4063
rect 12357 4029 12391 4063
rect 13277 4029 13311 4063
rect 22661 4029 22695 4063
rect 24501 4029 24535 4063
rect 52745 4029 52779 4063
rect 55965 4029 55999 4063
rect 2605 3961 2639 3995
rect 7205 3961 7239 3995
rect 8401 3961 8435 3995
rect 9505 3961 9539 3995
rect 11989 3961 12023 3995
rect 13921 3961 13955 3995
rect 15853 3961 15887 3995
rect 18705 3961 18739 3995
rect 20637 3961 20671 3995
rect 36553 3961 36587 3995
rect 1961 3893 1995 3927
rect 4169 3893 4203 3927
rect 6561 3893 6595 3927
rect 6745 3893 6779 3927
rect 7573 3893 7607 3927
rect 8493 3893 8527 3927
rect 10793 3893 10827 3927
rect 11897 3893 11931 3927
rect 15209 3893 15243 3927
rect 16865 3893 16899 3927
rect 17509 3893 17543 3927
rect 19349 3893 19383 3927
rect 19993 3893 20027 3927
rect 21281 3893 21315 3927
rect 22201 3893 22235 3927
rect 24041 3893 24075 3927
rect 25697 3893 25731 3927
rect 26249 3893 26283 3927
rect 51181 3893 51215 3927
rect 51825 3893 51859 3927
rect 53389 3893 53423 3927
rect 54033 3893 54067 3927
rect 55321 3893 55355 3927
rect 58173 3893 58207 3927
rect 17417 3689 17451 3723
rect 20269 3689 20303 3723
rect 21005 3689 21039 3723
rect 32137 3689 32171 3723
rect 3249 3621 3283 3655
rect 8217 3621 8251 3655
rect 9413 3621 9447 3655
rect 11529 3621 11563 3655
rect 12265 3621 12299 3655
rect 14841 3621 14875 3655
rect 18705 3621 18739 3655
rect 46949 3621 46983 3655
rect 52837 3621 52871 3655
rect 55321 3621 55355 3655
rect 6561 3553 6595 3587
rect 6837 3553 6871 3587
rect 14289 3553 14323 3587
rect 16037 3553 16071 3587
rect 19625 3553 19659 3587
rect 21741 3553 21775 3587
rect 51549 3553 51583 3587
rect 53481 3553 53515 3587
rect 56609 3553 56643 3587
rect 1869 3485 1903 3519
rect 4261 3485 4295 3519
rect 8401 3485 8435 3519
rect 9689 3485 9723 3519
rect 10885 3485 10919 3519
rect 11345 3485 11379 3519
rect 12081 3485 12115 3519
rect 12909 3485 12943 3519
rect 13369 3485 13403 3519
rect 15577 3485 15611 3519
rect 16293 3485 16327 3519
rect 18521 3485 18555 3519
rect 20177 3485 20211 3519
rect 21925 3485 21959 3519
rect 23213 3485 23247 3519
rect 23857 3485 23891 3519
rect 24869 3485 24903 3519
rect 25697 3485 25731 3519
rect 26801 3485 26835 3519
rect 27629 3485 27663 3519
rect 28733 3485 28767 3519
rect 30757 3485 30791 3519
rect 34805 3485 34839 3519
rect 35449 3485 35483 3519
rect 36093 3485 36127 3519
rect 36737 3485 36771 3519
rect 37565 3485 37599 3519
rect 38669 3485 38703 3519
rect 40049 3485 40083 3519
rect 40693 3485 40727 3519
rect 41337 3485 41371 3519
rect 42533 3485 42567 3519
rect 43177 3485 43211 3519
rect 45017 3485 45051 3519
rect 45661 3485 45695 3519
rect 46305 3485 46339 3519
rect 47777 3485 47811 3519
rect 48421 3485 48455 3519
rect 50261 3485 50295 3519
rect 50905 3485 50939 3519
rect 52193 3485 52227 3519
rect 54125 3485 54159 3519
rect 55965 3485 55999 3519
rect 57529 3485 57563 3519
rect 58173 3485 58207 3519
rect 2136 3417 2170 3451
rect 4528 3417 4562 3451
rect 14381 3417 14415 3451
rect 14841 3417 14875 3451
rect 17969 3417 18003 3451
rect 21097 3417 21131 3451
rect 31002 3417 31036 3451
rect 5641 3349 5675 3383
rect 10701 3349 10735 3383
rect 13553 3349 13587 3383
rect 14105 3349 14139 3383
rect 22569 3349 22603 3383
rect 1869 3145 1903 3179
rect 3801 3145 3835 3179
rect 5667 3145 5701 3179
rect 13553 3145 13587 3179
rect 14565 3145 14599 3179
rect 15209 3145 15243 3179
rect 15945 3145 15979 3179
rect 17417 3145 17451 3179
rect 23029 3145 23063 3179
rect 2666 3077 2700 3111
rect 5457 3077 5491 3111
rect 10425 3077 10459 3111
rect 18061 3077 18095 3111
rect 18797 3077 18831 3111
rect 18981 3077 19015 3111
rect 20453 3077 20487 3111
rect 21005 3077 21039 3111
rect 21189 3077 21223 3111
rect 22201 3077 22235 3111
rect 22385 3077 22419 3111
rect 1777 3009 1811 3043
rect 2421 3009 2455 3043
rect 4997 3009 5031 3043
rect 6745 3009 6779 3043
rect 7021 3009 7055 3043
rect 8033 3009 8067 3043
rect 8953 3009 8987 3043
rect 9505 3009 9539 3043
rect 9873 3009 9907 3043
rect 10793 3009 10827 3043
rect 11529 3009 11563 3043
rect 12909 3009 12943 3043
rect 13369 3009 13403 3043
rect 14381 3009 14415 3043
rect 15393 3009 15427 3043
rect 16129 3009 16163 3043
rect 17601 3009 17635 3043
rect 18245 3009 18279 3043
rect 19809 3009 19843 3043
rect 22845 3009 22879 3043
rect 54033 3009 54067 3043
rect 54677 3009 54711 3043
rect 55321 3009 55355 3043
rect 8585 2941 8619 2975
rect 20269 2941 20303 2975
rect 23857 2941 23891 2975
rect 33425 2941 33459 2975
rect 39221 2941 39255 2975
rect 43085 2941 43119 2975
rect 55965 2941 55999 2975
rect 56609 2941 56643 2975
rect 5825 2873 5859 2907
rect 11713 2873 11747 2907
rect 34713 2873 34747 2907
rect 37933 2873 37967 2907
rect 39865 2873 39899 2907
rect 41153 2873 41187 2907
rect 43729 2873 43763 2907
rect 45017 2873 45051 2907
rect 45661 2873 45695 2907
rect 48237 2873 48271 2907
rect 49525 2873 49559 2907
rect 50813 2873 50847 2907
rect 52745 2873 52779 2907
rect 57897 2873 57931 2907
rect 4813 2805 4847 2839
rect 5641 2805 5675 2839
rect 8401 2805 8435 2839
rect 8493 2805 8527 2839
rect 16865 2805 16899 2839
rect 19625 2805 19659 2839
rect 24501 2805 24535 2839
rect 25145 2805 25179 2839
rect 25789 2805 25823 2839
rect 26433 2805 26467 2839
rect 27629 2805 27663 2839
rect 28089 2805 28123 2839
rect 28917 2805 28951 2839
rect 29561 2805 29595 2839
rect 30021 2805 30055 2839
rect 30665 2805 30699 2839
rect 32137 2805 32171 2839
rect 32781 2805 32815 2839
rect 34069 2805 34103 2839
rect 35357 2805 35391 2839
rect 36001 2805 36035 2839
rect 37289 2805 37323 2839
rect 38577 2805 38611 2839
rect 40509 2805 40543 2839
rect 42441 2805 42475 2839
rect 44373 2805 44407 2839
rect 46305 2805 46339 2839
rect 47593 2805 47627 2839
rect 48881 2805 48915 2839
rect 50169 2805 50203 2839
rect 51457 2805 51491 2839
rect 53389 2805 53423 2839
rect 1777 2601 1811 2635
rect 6653 2601 6687 2635
rect 10425 2601 10459 2635
rect 11713 2601 11747 2635
rect 13461 2601 13495 2635
rect 14565 2601 14599 2635
rect 20361 2601 20395 2635
rect 22753 2601 22787 2635
rect 26985 2601 27019 2635
rect 55321 2601 55355 2635
rect 2237 2533 2271 2567
rect 3065 2533 3099 2567
rect 12449 2533 12483 2567
rect 16129 2533 16163 2567
rect 16865 2533 16899 2567
rect 17693 2533 17727 2567
rect 18705 2533 18739 2567
rect 21281 2533 21315 2567
rect 25789 2533 25823 2567
rect 27721 2533 27755 2567
rect 36001 2533 36035 2567
rect 39865 2533 39899 2567
rect 43729 2533 43763 2567
rect 47593 2533 47627 2567
rect 51457 2533 51491 2567
rect 54033 2533 54067 2567
rect 7573 2465 7607 2499
rect 32781 2465 32815 2499
rect 34713 2465 34747 2499
rect 37289 2465 37323 2499
rect 40509 2465 40543 2499
rect 42441 2465 42475 2499
rect 45017 2465 45051 2499
rect 48237 2465 48271 2499
rect 50169 2465 50203 2499
rect 52745 2465 52779 2499
rect 57897 2465 57931 2499
rect 1593 2397 1627 2431
rect 2421 2397 2455 2431
rect 3249 2397 3283 2431
rect 4261 2397 4295 2431
rect 5549 2397 5583 2431
rect 5825 2397 5859 2431
rect 7297 2397 7331 2431
rect 9229 2397 9263 2431
rect 10149 2397 10183 2431
rect 11529 2397 11563 2431
rect 12265 2397 12299 2431
rect 13277 2397 13311 2431
rect 14381 2397 14415 2431
rect 15117 2397 15151 2431
rect 16681 2397 16715 2431
rect 17877 2397 17911 2431
rect 19533 2397 19567 2431
rect 22201 2397 22235 2431
rect 22937 2397 22971 2431
rect 23397 2397 23431 2431
rect 24409 2397 24443 2431
rect 25145 2397 25179 2431
rect 26433 2397 26467 2431
rect 28365 2397 28399 2431
rect 29009 2397 29043 2431
rect 30113 2397 30147 2431
rect 30757 2397 30791 2431
rect 31217 2397 31251 2431
rect 32137 2397 32171 2431
rect 33425 2397 33459 2431
rect 35357 2397 35391 2431
rect 37933 2397 37967 2431
rect 38577 2397 38611 2431
rect 41153 2397 41187 2431
rect 43085 2397 43119 2431
rect 45661 2397 45695 2431
rect 46305 2397 46339 2431
rect 48881 2397 48915 2431
rect 50813 2397 50847 2431
rect 53389 2397 53423 2431
rect 55965 2397 55999 2431
rect 56609 2397 56643 2431
rect 6745 2329 6779 2363
rect 15945 2329 15979 2363
rect 18521 2329 18555 2363
rect 20453 2329 20487 2363
rect 21097 2329 21131 2363
rect 4445 2261 4479 2295
rect 9045 2261 9079 2295
rect 15301 2261 15335 2295
rect 19349 2261 19383 2295
rect 22017 2261 22051 2295
rect 23581 2261 23615 2295
<< metal1 >>
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 1762 57536 1768 57588
rect 1820 57576 1826 57588
rect 1949 57579 2007 57585
rect 1949 57576 1961 57579
rect 1820 57548 1961 57576
rect 1820 57536 1826 57548
rect 1949 57545 1961 57548
rect 1995 57545 2007 57579
rect 1949 57539 2007 57545
rect 3326 57536 3332 57588
rect 3384 57576 3390 57588
rect 3881 57579 3939 57585
rect 3881 57576 3893 57579
rect 3384 57548 3893 57576
rect 3384 57536 3390 57548
rect 3881 57545 3893 57548
rect 3927 57545 3939 57579
rect 3881 57539 3939 57545
rect 4890 57536 4896 57588
rect 4948 57576 4954 57588
rect 5077 57579 5135 57585
rect 5077 57576 5089 57579
rect 4948 57548 5089 57576
rect 4948 57536 4954 57548
rect 5077 57545 5089 57548
rect 5123 57545 5135 57579
rect 5077 57539 5135 57545
rect 6454 57536 6460 57588
rect 6512 57576 6518 57588
rect 6641 57579 6699 57585
rect 6641 57576 6653 57579
rect 6512 57548 6653 57576
rect 6512 57536 6518 57548
rect 6641 57545 6653 57548
rect 6687 57545 6699 57579
rect 6641 57539 6699 57545
rect 8018 57536 8024 57588
rect 8076 57576 8082 57588
rect 8205 57579 8263 57585
rect 8205 57576 8217 57579
rect 8076 57548 8217 57576
rect 8076 57536 8082 57548
rect 8205 57545 8217 57548
rect 8251 57545 8263 57579
rect 8205 57539 8263 57545
rect 9674 57536 9680 57588
rect 9732 57576 9738 57588
rect 9769 57579 9827 57585
rect 9769 57576 9781 57579
rect 9732 57548 9781 57576
rect 9732 57536 9738 57548
rect 9769 57545 9781 57548
rect 9815 57545 9827 57579
rect 9769 57539 9827 57545
rect 11146 57536 11152 57588
rect 11204 57576 11210 57588
rect 11609 57579 11667 57585
rect 11609 57576 11621 57579
rect 11204 57548 11621 57576
rect 11204 57536 11210 57548
rect 11609 57545 11621 57548
rect 11655 57545 11667 57579
rect 11609 57539 11667 57545
rect 12710 57536 12716 57588
rect 12768 57576 12774 57588
rect 12897 57579 12955 57585
rect 12897 57576 12909 57579
rect 12768 57548 12909 57576
rect 12768 57536 12774 57548
rect 12897 57545 12909 57548
rect 12943 57545 12955 57579
rect 12897 57539 12955 57545
rect 14274 57536 14280 57588
rect 14332 57576 14338 57588
rect 14461 57579 14519 57585
rect 14461 57576 14473 57579
rect 14332 57548 14473 57576
rect 14332 57536 14338 57548
rect 14461 57545 14473 57548
rect 14507 57545 14519 57579
rect 14461 57539 14519 57545
rect 15838 57536 15844 57588
rect 15896 57576 15902 57588
rect 16761 57579 16819 57585
rect 16761 57576 16773 57579
rect 15896 57548 16773 57576
rect 15896 57536 15902 57548
rect 16761 57545 16773 57548
rect 16807 57545 16819 57579
rect 16761 57539 16819 57545
rect 17402 57536 17408 57588
rect 17460 57576 17466 57588
rect 17681 57579 17739 57585
rect 17681 57576 17693 57579
rect 17460 57548 17693 57576
rect 17460 57536 17466 57548
rect 17681 57545 17693 57548
rect 17727 57545 17739 57579
rect 17681 57539 17739 57545
rect 19334 57536 19340 57588
rect 19392 57576 19398 57588
rect 19429 57579 19487 57585
rect 19429 57576 19441 57579
rect 19392 57548 19441 57576
rect 19392 57536 19398 57548
rect 19429 57545 19441 57548
rect 19475 57545 19487 57579
rect 19429 57539 19487 57545
rect 20714 57536 20720 57588
rect 20772 57576 20778 57588
rect 20809 57579 20867 57585
rect 20809 57576 20821 57579
rect 20772 57548 20821 57576
rect 20772 57536 20778 57548
rect 20809 57545 20821 57548
rect 20855 57545 20867 57579
rect 20809 57539 20867 57545
rect 22094 57536 22100 57588
rect 22152 57576 22158 57588
rect 22373 57579 22431 57585
rect 22373 57576 22385 57579
rect 22152 57548 22385 57576
rect 22152 57536 22158 57548
rect 22373 57545 22385 57548
rect 22419 57545 22431 57579
rect 22373 57539 22431 57545
rect 23658 57536 23664 57588
rect 23716 57576 23722 57588
rect 24581 57579 24639 57585
rect 24581 57576 24593 57579
rect 23716 57548 24593 57576
rect 23716 57536 23722 57548
rect 24581 57545 24593 57548
rect 24627 57545 24639 57579
rect 24581 57539 24639 57545
rect 25222 57536 25228 57588
rect 25280 57576 25286 57588
rect 25501 57579 25559 57585
rect 25501 57576 25513 57579
rect 25280 57548 25513 57576
rect 25280 57536 25286 57548
rect 25501 57545 25513 57548
rect 25547 57545 25559 57579
rect 25501 57539 25559 57545
rect 26786 57536 26792 57588
rect 26844 57576 26850 57588
rect 27157 57579 27215 57585
rect 27157 57576 27169 57579
rect 26844 57548 27169 57576
rect 26844 57536 26850 57548
rect 27157 57545 27169 57548
rect 27203 57545 27215 57579
rect 27157 57539 27215 57545
rect 28350 57536 28356 57588
rect 28408 57576 28414 57588
rect 28629 57579 28687 57585
rect 28629 57576 28641 57579
rect 28408 57548 28641 57576
rect 28408 57536 28414 57548
rect 28629 57545 28641 57548
rect 28675 57545 28687 57579
rect 28629 57539 28687 57545
rect 29914 57536 29920 57588
rect 29972 57576 29978 57588
rect 30193 57579 30251 57585
rect 30193 57576 30205 57579
rect 29972 57548 30205 57576
rect 29972 57536 29978 57548
rect 30193 57545 30205 57548
rect 30239 57545 30251 57579
rect 30193 57539 30251 57545
rect 31478 57536 31484 57588
rect 31536 57576 31542 57588
rect 32309 57579 32367 57585
rect 32309 57576 32321 57579
rect 31536 57548 32321 57576
rect 31536 57536 31542 57548
rect 32309 57545 32321 57548
rect 32355 57545 32367 57579
rect 32309 57539 32367 57545
rect 33134 57536 33140 57588
rect 33192 57576 33198 57588
rect 33321 57579 33379 57585
rect 33321 57576 33333 57579
rect 33192 57548 33333 57576
rect 33192 57536 33198 57548
rect 33321 57545 33333 57548
rect 33367 57545 33379 57579
rect 33321 57539 33379 57545
rect 34606 57536 34612 57588
rect 34664 57576 34670 57588
rect 34885 57579 34943 57585
rect 34885 57576 34897 57579
rect 34664 57548 34897 57576
rect 34664 57536 34670 57548
rect 34885 57545 34897 57548
rect 34931 57545 34943 57579
rect 34885 57539 34943 57545
rect 36170 57536 36176 57588
rect 36228 57576 36234 57588
rect 36449 57579 36507 57585
rect 36449 57576 36461 57579
rect 36228 57548 36461 57576
rect 36228 57536 36234 57548
rect 36449 57545 36461 57548
rect 36495 57545 36507 57579
rect 36449 57539 36507 57545
rect 37734 57536 37740 57588
rect 37792 57576 37798 57588
rect 38013 57579 38071 57585
rect 38013 57576 38025 57579
rect 37792 57548 38025 57576
rect 37792 57536 37798 57548
rect 38013 57545 38025 57548
rect 38059 57545 38071 57579
rect 38013 57539 38071 57545
rect 39298 57536 39304 57588
rect 39356 57576 39362 57588
rect 40037 57579 40095 57585
rect 40037 57576 40049 57579
rect 39356 57548 40049 57576
rect 39356 57536 39362 57548
rect 40037 57545 40049 57548
rect 40083 57545 40095 57579
rect 40037 57539 40095 57545
rect 40862 57536 40868 57588
rect 40920 57576 40926 57588
rect 41141 57579 41199 57585
rect 41141 57576 41153 57579
rect 40920 57548 41153 57576
rect 40920 57536 40926 57548
rect 41141 57545 41153 57548
rect 41187 57545 41199 57579
rect 41141 57539 41199 57545
rect 42426 57536 42432 57588
rect 42484 57576 42490 57588
rect 42705 57579 42763 57585
rect 42705 57576 42717 57579
rect 42484 57548 42717 57576
rect 42484 57536 42490 57548
rect 42705 57545 42717 57548
rect 42751 57545 42763 57579
rect 42705 57539 42763 57545
rect 44174 57536 44180 57588
rect 44232 57576 44238 57588
rect 44269 57579 44327 57585
rect 44269 57576 44281 57579
rect 44232 57548 44281 57576
rect 44232 57536 44238 57548
rect 44269 57545 44281 57548
rect 44315 57545 44327 57579
rect 44269 57539 44327 57545
rect 45554 57536 45560 57588
rect 45612 57576 45618 57588
rect 45833 57579 45891 57585
rect 45833 57576 45845 57579
rect 45612 57548 45845 57576
rect 45612 57536 45618 57548
rect 45833 57545 45845 57548
rect 45879 57545 45891 57579
rect 45833 57539 45891 57545
rect 47118 57536 47124 57588
rect 47176 57576 47182 57588
rect 47765 57579 47823 57585
rect 47765 57576 47777 57579
rect 47176 57548 47777 57576
rect 47176 57536 47182 57548
rect 47765 57545 47777 57548
rect 47811 57545 47823 57579
rect 47765 57539 47823 57545
rect 26326 57468 26332 57520
rect 26384 57508 26390 57520
rect 26384 57480 30052 57508
rect 26384 57468 26390 57480
rect 2133 57443 2191 57449
rect 2133 57409 2145 57443
rect 2179 57440 2191 57443
rect 2682 57440 2688 57452
rect 2179 57412 2688 57440
rect 2179 57409 2191 57412
rect 2133 57403 2191 57409
rect 2682 57400 2688 57412
rect 2740 57400 2746 57452
rect 4062 57440 4068 57452
rect 4023 57412 4068 57440
rect 4062 57400 4068 57412
rect 4120 57400 4126 57452
rect 5258 57440 5264 57452
rect 5219 57412 5264 57440
rect 5258 57400 5264 57412
rect 5316 57400 5322 57452
rect 6822 57440 6828 57452
rect 6783 57412 6828 57440
rect 6822 57400 6828 57412
rect 6880 57400 6886 57452
rect 8389 57443 8447 57449
rect 8389 57409 8401 57443
rect 8435 57409 8447 57443
rect 8389 57403 8447 57409
rect 9953 57443 10011 57449
rect 9953 57409 9965 57443
rect 9999 57409 10011 57443
rect 11790 57440 11796 57452
rect 11751 57412 11796 57440
rect 9953 57403 10011 57409
rect 8404 57304 8432 57403
rect 9968 57372 9996 57403
rect 11790 57400 11796 57412
rect 11848 57400 11854 57452
rect 13078 57440 13084 57452
rect 13039 57412 13084 57440
rect 13078 57400 13084 57412
rect 13136 57400 13142 57452
rect 14645 57443 14703 57449
rect 14645 57409 14657 57443
rect 14691 57440 14703 57443
rect 15746 57440 15752 57452
rect 14691 57412 15752 57440
rect 14691 57409 14703 57412
rect 14645 57403 14703 57409
rect 15746 57400 15752 57412
rect 15804 57400 15810 57452
rect 16942 57440 16948 57452
rect 16903 57412 16948 57440
rect 16942 57400 16948 57412
rect 17000 57400 17006 57452
rect 17494 57440 17500 57452
rect 17455 57412 17500 57440
rect 17494 57400 17500 57412
rect 17552 57400 17558 57452
rect 18690 57400 18696 57452
rect 18748 57440 18754 57452
rect 19245 57443 19303 57449
rect 19245 57440 19257 57443
rect 18748 57412 19257 57440
rect 18748 57400 18754 57412
rect 19245 57409 19257 57412
rect 19291 57409 19303 57443
rect 19245 57403 19303 57409
rect 19518 57400 19524 57452
rect 19576 57440 19582 57452
rect 20625 57443 20683 57449
rect 20625 57440 20637 57443
rect 19576 57412 20637 57440
rect 19576 57400 19582 57412
rect 20625 57409 20637 57412
rect 20671 57409 20683 57443
rect 22186 57440 22192 57452
rect 22147 57412 22192 57440
rect 20625 57403 20683 57409
rect 22186 57400 22192 57412
rect 22244 57400 22250 57452
rect 24394 57440 24400 57452
rect 24355 57412 24400 57440
rect 24394 57400 24400 57412
rect 24452 57400 24458 57452
rect 25314 57440 25320 57452
rect 25275 57412 25320 57440
rect 25314 57400 25320 57412
rect 25372 57400 25378 57452
rect 26970 57440 26976 57452
rect 26931 57412 26976 57440
rect 26970 57400 26976 57412
rect 27028 57400 27034 57452
rect 28442 57440 28448 57452
rect 28403 57412 28448 57440
rect 28442 57400 28448 57412
rect 28500 57400 28506 57452
rect 30024 57449 30052 57480
rect 30374 57468 30380 57520
rect 30432 57508 30438 57520
rect 30432 57480 35894 57508
rect 30432 57468 30438 57480
rect 30009 57443 30067 57449
rect 30009 57409 30021 57443
rect 30055 57409 30067 57443
rect 30009 57403 30067 57409
rect 30098 57400 30104 57452
rect 30156 57440 30162 57452
rect 32125 57443 32183 57449
rect 32125 57440 32137 57443
rect 30156 57412 32137 57440
rect 30156 57400 30162 57412
rect 32125 57409 32137 57412
rect 32171 57409 32183 57443
rect 32125 57403 32183 57409
rect 32214 57400 32220 57452
rect 32272 57440 32278 57452
rect 33137 57443 33195 57449
rect 33137 57440 33149 57443
rect 32272 57412 33149 57440
rect 32272 57400 32278 57412
rect 33137 57409 33149 57412
rect 33183 57409 33195 57443
rect 33137 57403 33195 57409
rect 33226 57400 33232 57452
rect 33284 57440 33290 57452
rect 34701 57443 34759 57449
rect 34701 57440 34713 57443
rect 33284 57412 34713 57440
rect 33284 57400 33290 57412
rect 34701 57409 34713 57412
rect 34747 57409 34759 57443
rect 35866 57440 35894 57480
rect 36265 57443 36323 57449
rect 36265 57440 36277 57443
rect 35866 57412 36277 57440
rect 34701 57403 34759 57409
rect 36265 57409 36277 57412
rect 36311 57409 36323 57443
rect 36265 57403 36323 57409
rect 37829 57443 37887 57449
rect 37829 57409 37841 57443
rect 37875 57409 37887 57443
rect 37829 57403 37887 57409
rect 39853 57443 39911 57449
rect 39853 57409 39865 57443
rect 39899 57409 39911 57443
rect 39853 57403 39911 57409
rect 19978 57372 19984 57384
rect 9968 57344 19984 57372
rect 19978 57332 19984 57344
rect 20036 57332 20042 57384
rect 37844 57372 37872 57403
rect 26206 57344 37872 57372
rect 18506 57304 18512 57316
rect 8404 57276 18512 57304
rect 18506 57264 18512 57276
rect 18564 57264 18570 57316
rect 24670 57264 24676 57316
rect 24728 57304 24734 57316
rect 26206 57304 26234 57344
rect 24728 57276 26234 57304
rect 24728 57264 24734 57276
rect 37182 57264 37188 57316
rect 37240 57304 37246 57316
rect 39868 57304 39896 57403
rect 40770 57400 40776 57452
rect 40828 57440 40834 57452
rect 40957 57443 41015 57449
rect 40957 57440 40969 57443
rect 40828 57412 40969 57440
rect 40828 57400 40834 57412
rect 40957 57409 40969 57412
rect 41003 57409 41015 57443
rect 42518 57440 42524 57452
rect 42479 57412 42524 57440
rect 40957 57403 41015 57409
rect 42518 57400 42524 57412
rect 42576 57400 42582 57452
rect 44082 57440 44088 57452
rect 44043 57412 44088 57440
rect 44082 57400 44088 57412
rect 44140 57400 44146 57452
rect 44174 57400 44180 57452
rect 44232 57440 44238 57452
rect 45649 57443 45707 57449
rect 45649 57440 45661 57443
rect 44232 57412 45661 57440
rect 44232 57400 44238 57412
rect 45649 57409 45661 57412
rect 45695 57409 45707 57443
rect 47578 57440 47584 57452
rect 47539 57412 47584 57440
rect 45649 57403 45707 57409
rect 47578 57400 47584 57412
rect 47636 57400 47642 57452
rect 48682 57400 48688 57452
rect 48740 57440 48746 57452
rect 48777 57443 48835 57449
rect 48777 57440 48789 57443
rect 48740 57412 48789 57440
rect 48740 57400 48746 57412
rect 48777 57409 48789 57412
rect 48823 57409 48835 57443
rect 48777 57403 48835 57409
rect 50154 57400 50160 57452
rect 50212 57440 50218 57452
rect 50341 57443 50399 57449
rect 50341 57440 50353 57443
rect 50212 57412 50353 57440
rect 50212 57400 50218 57412
rect 50341 57409 50353 57412
rect 50387 57409 50399 57443
rect 50341 57403 50399 57409
rect 51810 57400 51816 57452
rect 51868 57440 51874 57452
rect 51905 57443 51963 57449
rect 51905 57440 51917 57443
rect 51868 57412 51917 57440
rect 51868 57400 51874 57412
rect 51905 57409 51917 57412
rect 51951 57409 51963 57443
rect 51905 57403 51963 57409
rect 53374 57400 53380 57452
rect 53432 57440 53438 57452
rect 53469 57443 53527 57449
rect 53469 57440 53481 57443
rect 53432 57412 53481 57440
rect 53432 57400 53438 57412
rect 53469 57409 53481 57412
rect 53515 57409 53527 57443
rect 56594 57440 56600 57452
rect 56555 57412 56600 57440
rect 53469 57403 53527 57409
rect 56594 57400 56600 57412
rect 56652 57400 56658 57452
rect 57977 57443 58035 57449
rect 57977 57409 57989 57443
rect 58023 57440 58035 57443
rect 58066 57440 58072 57452
rect 58023 57412 58072 57440
rect 58023 57409 58035 57412
rect 57977 57403 58035 57409
rect 58066 57400 58072 57412
rect 58124 57400 58130 57452
rect 54938 57332 54944 57384
rect 54996 57372 55002 57384
rect 55309 57375 55367 57381
rect 55309 57372 55321 57375
rect 54996 57344 55321 57372
rect 54996 57332 55002 57344
rect 55309 57341 55321 57344
rect 55355 57341 55367 57375
rect 55309 57335 55367 57341
rect 37240 57276 39896 57304
rect 37240 57264 37246 57276
rect 2682 57236 2688 57248
rect 2643 57208 2688 57236
rect 2682 57196 2688 57208
rect 2740 57196 2746 57248
rect 18693 57239 18751 57245
rect 18693 57205 18705 57239
rect 18739 57236 18751 57239
rect 18966 57236 18972 57248
rect 18739 57208 18972 57236
rect 18739 57205 18751 57208
rect 18693 57199 18751 57205
rect 18966 57196 18972 57208
rect 19024 57196 19030 57248
rect 20073 57239 20131 57245
rect 20073 57205 20085 57239
rect 20119 57236 20131 57239
rect 20162 57236 20168 57248
rect 20119 57208 20168 57236
rect 20119 57205 20131 57208
rect 20073 57199 20131 57205
rect 20162 57196 20168 57208
rect 20220 57196 20226 57248
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 18690 57032 18696 57044
rect 18651 57004 18696 57032
rect 18690 56992 18696 57004
rect 18748 56992 18754 57044
rect 19518 57032 19524 57044
rect 19479 57004 19524 57032
rect 19518 56992 19524 57004
rect 19576 56992 19582 57044
rect 19978 57032 19984 57044
rect 19939 57004 19984 57032
rect 19978 56992 19984 57004
rect 20036 56992 20042 57044
rect 57514 57032 57520 57044
rect 57475 57004 57520 57032
rect 57514 56992 57520 57004
rect 57572 56992 57578 57044
rect 6822 56924 6828 56976
rect 6880 56964 6886 56976
rect 18782 56964 18788 56976
rect 6880 56936 18788 56964
rect 6880 56924 6886 56936
rect 18782 56924 18788 56936
rect 18840 56924 18846 56976
rect 19334 56924 19340 56976
rect 19392 56924 19398 56976
rect 11790 56856 11796 56908
rect 11848 56896 11854 56908
rect 19352 56896 19380 56924
rect 11848 56868 19380 56896
rect 11848 56856 11854 56868
rect 1394 56828 1400 56840
rect 1355 56800 1400 56828
rect 1394 56788 1400 56800
rect 1452 56788 1458 56840
rect 17497 56831 17555 56837
rect 17497 56797 17509 56831
rect 17543 56828 17555 56831
rect 18138 56828 18144 56840
rect 17543 56800 18144 56828
rect 17543 56797 17555 56800
rect 17497 56791 17555 56797
rect 18138 56788 18144 56800
rect 18196 56828 18202 56840
rect 18509 56831 18567 56837
rect 18509 56828 18521 56831
rect 18196 56800 18521 56828
rect 18196 56788 18202 56800
rect 18509 56797 18521 56800
rect 18555 56797 18567 56831
rect 18509 56791 18567 56797
rect 19337 56831 19395 56837
rect 19337 56797 19349 56831
rect 19383 56797 19395 56831
rect 20162 56828 20168 56840
rect 20123 56800 20168 56828
rect 19337 56791 19395 56797
rect 18049 56763 18107 56769
rect 18049 56729 18061 56763
rect 18095 56760 18107 56763
rect 19058 56760 19064 56772
rect 18095 56732 19064 56760
rect 18095 56729 18107 56732
rect 18049 56723 18107 56729
rect 19058 56720 19064 56732
rect 19116 56760 19122 56772
rect 19352 56760 19380 56791
rect 20162 56788 20168 56800
rect 20220 56788 20226 56840
rect 57882 56788 57888 56840
rect 57940 56828 57946 56840
rect 58161 56831 58219 56837
rect 58161 56828 58173 56831
rect 57940 56800 58173 56828
rect 57940 56788 57946 56800
rect 58161 56797 58173 56800
rect 58207 56797 58219 56831
rect 58161 56791 58219 56797
rect 42337 56763 42395 56769
rect 42337 56760 42349 56763
rect 19116 56732 19380 56760
rect 26206 56732 42349 56760
rect 19116 56720 19122 56732
rect 20714 56692 20720 56704
rect 20675 56664 20720 56692
rect 20714 56652 20720 56664
rect 20772 56652 20778 56704
rect 23382 56652 23388 56704
rect 23440 56692 23446 56704
rect 26206 56692 26234 56732
rect 42337 56729 42349 56732
rect 42383 56760 42395 56763
rect 42518 56760 42524 56772
rect 42383 56732 42524 56760
rect 42383 56729 42395 56732
rect 42337 56723 42395 56729
rect 42518 56720 42524 56732
rect 42576 56720 42582 56772
rect 40770 56692 40776 56704
rect 23440 56664 26234 56692
rect 40731 56664 40776 56692
rect 23440 56652 23446 56664
rect 40770 56652 40776 56664
rect 40828 56652 40834 56704
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 13078 56448 13084 56500
rect 13136 56488 13142 56500
rect 13541 56491 13599 56497
rect 13541 56488 13553 56491
rect 13136 56460 13553 56488
rect 13136 56448 13142 56460
rect 13541 56457 13553 56460
rect 13587 56457 13599 56491
rect 15746 56488 15752 56500
rect 15707 56460 15752 56488
rect 13541 56451 13599 56457
rect 15746 56448 15752 56460
rect 15804 56448 15810 56500
rect 17494 56488 17500 56500
rect 17455 56460 17500 56488
rect 17494 56448 17500 56460
rect 17552 56448 17558 56500
rect 18782 56488 18788 56500
rect 18743 56460 18788 56488
rect 18782 56448 18788 56460
rect 18840 56448 18846 56500
rect 21269 56491 21327 56497
rect 21269 56457 21281 56491
rect 21315 56488 21327 56491
rect 22186 56488 22192 56500
rect 21315 56460 22192 56488
rect 21315 56457 21327 56460
rect 21269 56451 21327 56457
rect 22186 56448 22192 56460
rect 22244 56448 22250 56500
rect 22741 56491 22799 56497
rect 22741 56457 22753 56491
rect 22787 56488 22799 56491
rect 24394 56488 24400 56500
rect 22787 56460 24400 56488
rect 22787 56457 22799 56460
rect 22741 56451 22799 56457
rect 24394 56448 24400 56460
rect 24452 56448 24458 56500
rect 24670 56488 24676 56500
rect 24631 56460 24676 56488
rect 24670 56448 24676 56460
rect 24728 56448 24734 56500
rect 25317 56491 25375 56497
rect 25317 56457 25329 56491
rect 25363 56488 25375 56491
rect 26326 56488 26332 56500
rect 25363 56460 26332 56488
rect 25363 56457 25375 56460
rect 25317 56451 25375 56457
rect 26326 56448 26332 56460
rect 26384 56448 26390 56500
rect 26421 56491 26479 56497
rect 26421 56457 26433 56491
rect 26467 56488 26479 56491
rect 26970 56488 26976 56500
rect 26467 56460 26976 56488
rect 26467 56457 26479 56460
rect 26421 56451 26479 56457
rect 26970 56448 26976 56460
rect 27028 56448 27034 56500
rect 27157 56491 27215 56497
rect 27157 56457 27169 56491
rect 27203 56488 27215 56491
rect 28442 56488 28448 56500
rect 27203 56460 28448 56488
rect 27203 56457 27215 56460
rect 27157 56451 27215 56457
rect 28442 56448 28448 56460
rect 28500 56448 28506 56500
rect 28721 56491 28779 56497
rect 28721 56457 28733 56491
rect 28767 56488 28779 56491
rect 30098 56488 30104 56500
rect 28767 56460 30104 56488
rect 28767 56457 28779 56460
rect 28721 56451 28779 56457
rect 30098 56448 30104 56460
rect 30156 56448 30162 56500
rect 31297 56491 31355 56497
rect 31297 56457 31309 56491
rect 31343 56488 31355 56491
rect 32214 56488 32220 56500
rect 31343 56460 32220 56488
rect 31343 56457 31355 56460
rect 31297 56451 31355 56457
rect 32214 56448 32220 56460
rect 32272 56448 32278 56500
rect 32309 56491 32367 56497
rect 32309 56457 32321 56491
rect 32355 56488 32367 56491
rect 33226 56488 33232 56500
rect 32355 56460 33232 56488
rect 32355 56457 32367 56460
rect 32309 56451 32367 56457
rect 33226 56448 33232 56460
rect 33284 56448 33290 56500
rect 35713 56491 35771 56497
rect 35713 56457 35725 56491
rect 35759 56488 35771 56491
rect 37182 56488 37188 56500
rect 35759 56460 37188 56488
rect 35759 56457 35771 56460
rect 35713 56451 35771 56457
rect 37182 56448 37188 56460
rect 37240 56448 37246 56500
rect 43993 56491 44051 56497
rect 43993 56457 44005 56491
rect 44039 56488 44051 56491
rect 44174 56488 44180 56500
rect 44039 56460 44180 56488
rect 44039 56457 44051 56460
rect 43993 56451 44051 56457
rect 44174 56448 44180 56460
rect 44232 56448 44238 56500
rect 46293 56491 46351 56497
rect 46293 56457 46305 56491
rect 46339 56488 46351 56491
rect 47578 56488 47584 56500
rect 46339 56460 47584 56488
rect 46339 56457 46351 56460
rect 46293 56451 46351 56457
rect 47578 56448 47584 56460
rect 47636 56448 47642 56500
rect 17037 56423 17095 56429
rect 17037 56389 17049 56423
rect 17083 56420 17095 56423
rect 17083 56392 18368 56420
rect 17083 56389 17095 56392
rect 17037 56383 17095 56389
rect 13725 56355 13783 56361
rect 13725 56321 13737 56355
rect 13771 56352 13783 56355
rect 14182 56352 14188 56364
rect 13771 56324 14188 56352
rect 13771 56321 13783 56324
rect 13725 56315 13783 56321
rect 14182 56312 14188 56324
rect 14240 56312 14246 56364
rect 15930 56352 15936 56364
rect 15891 56324 15936 56352
rect 15930 56312 15936 56324
rect 15988 56312 15994 56364
rect 17678 56352 17684 56364
rect 17639 56324 17684 56352
rect 17678 56312 17684 56324
rect 17736 56312 17742 56364
rect 18340 56361 18368 56392
rect 19426 56380 19432 56432
rect 19484 56420 19490 56432
rect 20714 56420 20720 56432
rect 19484 56392 20720 56420
rect 19484 56380 19490 56392
rect 18325 56355 18383 56361
rect 18325 56321 18337 56355
rect 18371 56352 18383 56355
rect 18874 56352 18880 56364
rect 18371 56324 18880 56352
rect 18371 56321 18383 56324
rect 18325 56315 18383 56321
rect 18874 56312 18880 56324
rect 18932 56312 18938 56364
rect 18966 56312 18972 56364
rect 19024 56352 19030 56364
rect 19613 56355 19671 56361
rect 19024 56324 19117 56352
rect 19024 56312 19030 56324
rect 19613 56321 19625 56355
rect 19659 56352 19671 56355
rect 19978 56352 19984 56364
rect 19659 56324 19984 56352
rect 19659 56321 19671 56324
rect 19613 56315 19671 56321
rect 19978 56312 19984 56324
rect 20036 56312 20042 56364
rect 20272 56361 20300 56392
rect 20714 56380 20720 56392
rect 20772 56380 20778 56432
rect 20257 56355 20315 56361
rect 20257 56321 20269 56355
rect 20303 56321 20315 56355
rect 20257 56315 20315 56321
rect 20898 56312 20904 56364
rect 20956 56352 20962 56364
rect 21085 56355 21143 56361
rect 21085 56352 21097 56355
rect 20956 56324 21097 56352
rect 20956 56312 20962 56324
rect 21085 56321 21097 56324
rect 21131 56321 21143 56355
rect 21085 56315 21143 56321
rect 21726 56312 21732 56364
rect 21784 56352 21790 56364
rect 21913 56355 21971 56361
rect 21913 56352 21925 56355
rect 21784 56324 21925 56352
rect 21784 56312 21790 56324
rect 21913 56321 21925 56324
rect 21959 56321 21971 56355
rect 22554 56352 22560 56364
rect 22515 56324 22560 56352
rect 21913 56315 21971 56321
rect 22554 56312 22560 56324
rect 22612 56312 22618 56364
rect 23014 56312 23020 56364
rect 23072 56352 23078 56364
rect 23201 56355 23259 56361
rect 23201 56352 23213 56355
rect 23072 56324 23213 56352
rect 23072 56312 23078 56324
rect 23201 56321 23213 56324
rect 23247 56321 23259 56355
rect 23201 56315 23259 56321
rect 23750 56312 23756 56364
rect 23808 56352 23814 56364
rect 23845 56355 23903 56361
rect 23845 56352 23857 56355
rect 23808 56324 23857 56352
rect 23808 56312 23814 56324
rect 23845 56321 23857 56324
rect 23891 56321 23903 56355
rect 23845 56315 23903 56321
rect 24394 56312 24400 56364
rect 24452 56352 24458 56364
rect 24489 56355 24547 56361
rect 24489 56352 24501 56355
rect 24452 56324 24501 56352
rect 24452 56312 24458 56324
rect 24489 56321 24501 56324
rect 24535 56321 24547 56355
rect 25130 56352 25136 56364
rect 25091 56324 25136 56352
rect 24489 56315 24547 56321
rect 25130 56312 25136 56324
rect 25188 56312 25194 56364
rect 26050 56312 26056 56364
rect 26108 56352 26114 56364
rect 26237 56355 26295 56361
rect 26237 56352 26249 56355
rect 26108 56324 26249 56352
rect 26108 56312 26114 56324
rect 26237 56321 26249 56324
rect 26283 56321 26295 56355
rect 26237 56315 26295 56321
rect 26786 56312 26792 56364
rect 26844 56352 26850 56364
rect 26973 56355 27031 56361
rect 26973 56352 26985 56355
rect 26844 56324 26985 56352
rect 26844 56312 26850 56324
rect 26973 56321 26985 56324
rect 27019 56321 27031 56355
rect 26973 56315 27031 56321
rect 27982 56312 27988 56364
rect 28040 56352 28046 56364
rect 28537 56355 28595 56361
rect 28537 56352 28549 56355
rect 28040 56324 28549 56352
rect 28040 56312 28046 56324
rect 28537 56321 28549 56324
rect 28583 56321 28595 56355
rect 29178 56352 29184 56364
rect 29139 56324 29184 56352
rect 28537 56315 28595 56321
rect 29178 56312 29184 56324
rect 29236 56312 29242 56364
rect 29914 56312 29920 56364
rect 29972 56352 29978 56364
rect 30469 56355 30527 56361
rect 30469 56352 30481 56355
rect 29972 56324 30481 56352
rect 29972 56312 29978 56324
rect 30469 56321 30481 56324
rect 30515 56321 30527 56355
rect 30469 56315 30527 56321
rect 30926 56312 30932 56364
rect 30984 56352 30990 56364
rect 31113 56355 31171 56361
rect 31113 56352 31125 56355
rect 30984 56324 31125 56352
rect 30984 56312 30990 56324
rect 31113 56321 31125 56324
rect 31159 56321 31171 56355
rect 32122 56352 32128 56364
rect 32083 56324 32128 56352
rect 31113 56315 31171 56321
rect 32122 56312 32128 56324
rect 32180 56352 32186 56364
rect 32769 56355 32827 56361
rect 32769 56352 32781 56355
rect 32180 56324 32781 56352
rect 32180 56312 32186 56324
rect 32769 56321 32781 56324
rect 32815 56321 32827 56355
rect 32769 56315 32827 56321
rect 35529 56355 35587 56361
rect 35529 56321 35541 56355
rect 35575 56352 35587 56355
rect 35710 56352 35716 56364
rect 35575 56324 35716 56352
rect 35575 56321 35587 56324
rect 35529 56315 35587 56321
rect 35710 56312 35716 56324
rect 35768 56352 35774 56364
rect 36173 56355 36231 56361
rect 36173 56352 36185 56355
rect 35768 56324 36185 56352
rect 35768 56312 35774 56324
rect 36173 56321 36185 56324
rect 36219 56321 36231 56355
rect 43806 56352 43812 56364
rect 43767 56324 43812 56352
rect 36173 56315 36231 56321
rect 43806 56312 43812 56324
rect 43864 56352 43870 56364
rect 44453 56355 44511 56361
rect 44453 56352 44465 56355
rect 43864 56324 44465 56352
rect 43864 56312 43870 56324
rect 44453 56321 44465 56324
rect 44499 56321 44511 56355
rect 44453 56315 44511 56321
rect 46109 56355 46167 56361
rect 46109 56321 46121 56355
rect 46155 56352 46167 56355
rect 46750 56352 46756 56364
rect 46155 56324 46756 56352
rect 46155 56321 46167 56324
rect 46109 56315 46167 56321
rect 46750 56312 46756 56324
rect 46808 56312 46814 56364
rect 58161 56355 58219 56361
rect 58161 56321 58173 56355
rect 58207 56352 58219 56355
rect 58434 56352 58440 56364
rect 58207 56324 58440 56352
rect 58207 56321 58219 56324
rect 58161 56315 58219 56321
rect 58434 56312 58440 56324
rect 58492 56312 58498 56364
rect 5258 56244 5264 56296
rect 5316 56284 5322 56296
rect 18984 56284 19012 56312
rect 20162 56284 20168 56296
rect 5316 56256 18184 56284
rect 18984 56256 20168 56284
rect 5316 56244 5322 56256
rect 4062 56176 4068 56228
rect 4120 56216 4126 56228
rect 18156 56225 18184 56256
rect 20162 56244 20168 56256
rect 20220 56244 20226 56296
rect 40770 56284 40776 56296
rect 26206 56256 40776 56284
rect 18141 56219 18199 56225
rect 4120 56188 18000 56216
rect 4120 56176 4126 56188
rect 14182 56148 14188 56160
rect 14143 56120 14188 56148
rect 14182 56108 14188 56120
rect 14240 56108 14246 56160
rect 17972 56148 18000 56188
rect 18141 56185 18153 56219
rect 18187 56185 18199 56219
rect 19429 56219 19487 56225
rect 19429 56216 19441 56219
rect 18141 56179 18199 56185
rect 18248 56188 19441 56216
rect 18248 56148 18276 56188
rect 19429 56185 19441 56188
rect 19475 56185 19487 56219
rect 19429 56179 19487 56185
rect 22097 56219 22155 56225
rect 22097 56185 22109 56219
rect 22143 56216 22155 56219
rect 26206 56216 26234 56256
rect 40770 56244 40776 56256
rect 40828 56244 40834 56296
rect 29914 56216 29920 56228
rect 22143 56188 26234 56216
rect 29875 56188 29920 56216
rect 22143 56185 22155 56188
rect 22097 56179 22155 56185
rect 29914 56176 29920 56188
rect 29972 56176 29978 56228
rect 30653 56219 30711 56225
rect 30653 56185 30665 56219
rect 30699 56216 30711 56219
rect 44082 56216 44088 56228
rect 30699 56188 44088 56216
rect 30699 56185 30711 56188
rect 30653 56179 30711 56185
rect 44082 56176 44088 56188
rect 44140 56176 44146 56228
rect 20070 56148 20076 56160
rect 17972 56120 18276 56148
rect 20031 56120 20076 56148
rect 20070 56108 20076 56120
rect 20128 56108 20134 56160
rect 23382 56148 23388 56160
rect 23343 56120 23388 56148
rect 23382 56108 23388 56120
rect 23440 56108 23446 56160
rect 24029 56151 24087 56157
rect 24029 56117 24041 56151
rect 24075 56148 24087 56151
rect 25314 56148 25320 56160
rect 24075 56120 25320 56148
rect 24075 56117 24087 56120
rect 24029 56111 24087 56117
rect 25314 56108 25320 56120
rect 25372 56108 25378 56160
rect 27982 56148 27988 56160
rect 27943 56120 27988 56148
rect 27982 56108 27988 56120
rect 28040 56108 28046 56160
rect 29365 56151 29423 56157
rect 29365 56117 29377 56151
rect 29411 56148 29423 56151
rect 30374 56148 30380 56160
rect 29411 56120 30380 56148
rect 29411 56117 29423 56120
rect 29365 56111 29423 56117
rect 30374 56108 30380 56120
rect 30432 56108 30438 56160
rect 46750 56148 46756 56160
rect 46711 56120 46756 56148
rect 46750 56108 46756 56120
rect 46808 56108 46814 56160
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 2682 55904 2688 55956
rect 2740 55944 2746 55956
rect 20070 55944 20076 55956
rect 2740 55916 20076 55944
rect 2740 55904 2746 55916
rect 20070 55904 20076 55916
rect 20128 55904 20134 55956
rect 16942 55836 16948 55888
rect 17000 55876 17006 55888
rect 17497 55879 17555 55885
rect 17497 55876 17509 55879
rect 17000 55848 17509 55876
rect 17000 55836 17006 55848
rect 17497 55845 17509 55848
rect 17543 55845 17555 55879
rect 18506 55876 18512 55888
rect 18467 55848 18512 55876
rect 17497 55839 17555 55845
rect 18506 55836 18512 55848
rect 18564 55836 18570 55888
rect 19334 55836 19340 55888
rect 19392 55876 19398 55888
rect 19613 55879 19671 55885
rect 19613 55876 19625 55879
rect 19392 55848 19625 55876
rect 19392 55836 19398 55848
rect 19613 55845 19625 55848
rect 19659 55845 19671 55879
rect 19613 55839 19671 55845
rect 20070 55768 20076 55820
rect 20128 55808 20134 55820
rect 22373 55811 22431 55817
rect 22373 55808 22385 55811
rect 20128 55780 22385 55808
rect 20128 55768 20134 55780
rect 22373 55777 22385 55780
rect 22419 55808 22431 55811
rect 22554 55808 22560 55820
rect 22419 55780 22560 55808
rect 22419 55777 22431 55780
rect 22373 55771 22431 55777
rect 22554 55768 22560 55780
rect 22612 55768 22618 55820
rect 1394 55740 1400 55752
rect 1355 55712 1400 55740
rect 1394 55700 1400 55712
rect 1452 55700 1458 55752
rect 17681 55743 17739 55749
rect 17681 55709 17693 55743
rect 17727 55740 17739 55743
rect 17770 55740 17776 55752
rect 17727 55712 17776 55740
rect 17727 55709 17739 55712
rect 17681 55703 17739 55709
rect 17770 55700 17776 55712
rect 17828 55700 17834 55752
rect 18693 55743 18751 55749
rect 18693 55709 18705 55743
rect 18739 55740 18751 55743
rect 18782 55740 18788 55752
rect 18739 55712 18788 55740
rect 18739 55709 18751 55712
rect 18693 55703 18751 55709
rect 18782 55700 18788 55712
rect 18840 55700 18846 55752
rect 19797 55743 19855 55749
rect 19797 55709 19809 55743
rect 19843 55740 19855 55743
rect 19843 55712 20300 55740
rect 19843 55709 19855 55712
rect 19797 55703 19855 55709
rect 20272 55616 20300 55712
rect 15930 55564 15936 55616
rect 15988 55604 15994 55616
rect 16117 55607 16175 55613
rect 16117 55604 16129 55607
rect 15988 55576 16129 55604
rect 15988 55564 15994 55576
rect 16117 55573 16129 55576
rect 16163 55604 16175 55607
rect 16482 55604 16488 55616
rect 16163 55576 16488 55604
rect 16163 55573 16175 55576
rect 16117 55567 16175 55573
rect 16482 55564 16488 55576
rect 16540 55564 16546 55616
rect 17034 55604 17040 55616
rect 16995 55576 17040 55604
rect 17034 55564 17040 55576
rect 17092 55564 17098 55616
rect 20254 55604 20260 55616
rect 20215 55576 20260 55604
rect 20254 55564 20260 55576
rect 20312 55564 20318 55616
rect 20898 55604 20904 55616
rect 20859 55576 20904 55604
rect 20898 55564 20904 55576
rect 20956 55564 20962 55616
rect 21726 55604 21732 55616
rect 21687 55576 21732 55604
rect 21726 55564 21732 55576
rect 21784 55564 21790 55616
rect 23014 55604 23020 55616
rect 22975 55576 23020 55604
rect 23014 55564 23020 55576
rect 23072 55564 23078 55616
rect 23750 55604 23756 55616
rect 23711 55576 23756 55604
rect 23750 55564 23756 55576
rect 23808 55564 23814 55616
rect 24394 55604 24400 55616
rect 24355 55576 24400 55604
rect 24394 55564 24400 55576
rect 24452 55564 24458 55616
rect 25041 55607 25099 55613
rect 25041 55573 25053 55607
rect 25087 55604 25099 55607
rect 25130 55604 25136 55616
rect 25087 55576 25136 55604
rect 25087 55573 25099 55576
rect 25041 55567 25099 55573
rect 25130 55564 25136 55576
rect 25188 55564 25194 55616
rect 26050 55604 26056 55616
rect 26011 55576 26056 55604
rect 26050 55564 26056 55576
rect 26108 55564 26114 55616
rect 26786 55604 26792 55616
rect 26747 55576 26792 55604
rect 26786 55564 26792 55576
rect 26844 55564 26850 55616
rect 29178 55564 29184 55616
rect 29236 55604 29242 55616
rect 29549 55607 29607 55613
rect 29549 55604 29561 55607
rect 29236 55576 29561 55604
rect 29236 55564 29242 55576
rect 29549 55573 29561 55576
rect 29595 55573 29607 55607
rect 30926 55604 30932 55616
rect 30887 55576 30932 55604
rect 29549 55567 29607 55573
rect 30926 55564 30932 55576
rect 30984 55564 30990 55616
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 17770 55332 17776 55344
rect 17731 55304 17776 55332
rect 17770 55292 17776 55304
rect 17828 55292 17834 55344
rect 18782 55332 18788 55344
rect 18743 55304 18788 55332
rect 18782 55292 18788 55304
rect 18840 55292 18846 55344
rect 19794 55332 19800 55344
rect 19755 55304 19800 55332
rect 19794 55292 19800 55304
rect 19852 55332 19858 55344
rect 19978 55332 19984 55344
rect 19852 55304 19984 55332
rect 19852 55292 19858 55304
rect 19978 55292 19984 55304
rect 20036 55292 20042 55344
rect 58158 55128 58164 55140
rect 58119 55100 58164 55128
rect 58158 55088 58164 55100
rect 58216 55088 58222 55140
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 1394 54652 1400 54664
rect 1355 54624 1400 54652
rect 1394 54612 1400 54624
rect 1452 54612 1458 54664
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 57882 53932 57888 53984
rect 57940 53972 57946 53984
rect 58161 53975 58219 53981
rect 58161 53972 58173 53975
rect 57940 53944 58173 53972
rect 57940 53932 57946 53944
rect 58161 53941 58173 53944
rect 58207 53941 58219 53975
rect 58161 53935 58219 53941
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 1394 53564 1400 53576
rect 1355 53536 1400 53564
rect 1394 53524 1400 53536
rect 1452 53524 1458 53576
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 1394 52476 1400 52488
rect 1355 52448 1400 52476
rect 1394 52436 1400 52448
rect 1452 52436 1458 52488
rect 57882 52436 57888 52488
rect 57940 52476 57946 52488
rect 58161 52479 58219 52485
rect 58161 52476 58173 52479
rect 57940 52448 58173 52476
rect 57940 52436 57946 52448
rect 58161 52445 58173 52448
rect 58207 52445 58219 52479
rect 58161 52439 58219 52445
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 1394 51388 1400 51400
rect 1355 51360 1400 51388
rect 1394 51348 1400 51360
rect 1452 51348 1458 51400
rect 58158 51388 58164 51400
rect 58119 51360 58164 51388
rect 58158 51348 58164 51360
rect 58216 51348 58222 51400
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 16206 50328 16212 50380
rect 16264 50368 16270 50380
rect 20898 50368 20904 50380
rect 16264 50340 20904 50368
rect 16264 50328 16270 50340
rect 20898 50328 20904 50340
rect 20956 50328 20962 50380
rect 1394 50300 1400 50312
rect 1355 50272 1400 50300
rect 1394 50260 1400 50272
rect 1452 50260 1458 50312
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 58158 49756 58164 49768
rect 58119 49728 58164 49756
rect 58158 49716 58164 49728
rect 58216 49716 58222 49768
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 1394 49212 1400 49224
rect 1355 49184 1400 49212
rect 1394 49172 1400 49184
rect 1452 49172 1458 49224
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 58158 48532 58164 48544
rect 58119 48504 58164 48532
rect 58158 48492 58164 48504
rect 58216 48492 58222 48544
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 1394 48124 1400 48136
rect 1355 48096 1400 48124
rect 1394 48084 1400 48096
rect 1452 48084 1458 48136
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 58158 47036 58164 47048
rect 58119 47008 58164 47036
rect 58158 46996 58164 47008
rect 58216 46996 58222 47048
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 58158 45948 58164 45960
rect 58119 45920 58164 45948
rect 58158 45908 58164 45920
rect 58216 45908 58222 45960
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 13630 44820 13636 44872
rect 13688 44860 13694 44872
rect 24394 44860 24400 44872
rect 13688 44832 24400 44860
rect 13688 44820 13694 44832
rect 24394 44820 24400 44832
rect 24452 44820 24458 44872
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 58158 44248 58164 44260
rect 58119 44220 58164 44248
rect 58158 44208 58164 44220
rect 58216 44208 58222 44260
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 58158 43092 58164 43104
rect 58119 43064 58164 43092
rect 58158 43052 58164 43064
rect 58216 43052 58222 43104
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 16574 42548 16580 42560
rect 16535 42520 16580 42548
rect 16574 42508 16580 42520
rect 16632 42508 16638 42560
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 16666 42208 16672 42220
rect 16627 42180 16672 42208
rect 16666 42168 16672 42180
rect 16724 42168 16730 42220
rect 16853 42211 16911 42217
rect 16853 42177 16865 42211
rect 16899 42208 16911 42211
rect 16942 42208 16948 42220
rect 16899 42180 16948 42208
rect 16899 42177 16911 42180
rect 16853 42171 16911 42177
rect 16942 42168 16948 42180
rect 17000 42168 17006 42220
rect 16022 41964 16028 42016
rect 16080 42004 16086 42016
rect 17037 42007 17095 42013
rect 17037 42004 17049 42007
rect 16080 41976 17049 42004
rect 16080 41964 16086 41976
rect 17037 41973 17049 41976
rect 17083 41973 17095 42007
rect 17037 41967 17095 41973
rect 17310 41964 17316 42016
rect 17368 42004 17374 42016
rect 17773 42007 17831 42013
rect 17773 42004 17785 42007
rect 17368 41976 17785 42004
rect 17368 41964 17374 41976
rect 17773 41973 17785 41976
rect 17819 42004 17831 42007
rect 18598 42004 18604 42016
rect 17819 41976 18604 42004
rect 17819 41973 17831 41976
rect 17773 41967 17831 41973
rect 18598 41964 18604 41976
rect 18656 41964 18662 42016
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 14734 41692 14740 41744
rect 14792 41732 14798 41744
rect 18598 41732 18604 41744
rect 14792 41704 15884 41732
rect 18511 41704 18604 41732
rect 14792 41692 14798 41704
rect 13906 41624 13912 41676
rect 13964 41664 13970 41676
rect 15856 41664 15884 41704
rect 18598 41692 18604 41704
rect 18656 41732 18662 41744
rect 24302 41732 24308 41744
rect 18656 41704 24308 41732
rect 18656 41692 18662 41704
rect 24302 41692 24308 41704
rect 24360 41692 24366 41744
rect 13964 41636 15424 41664
rect 13964 41624 13970 41636
rect 14476 41605 14504 41636
rect 14369 41599 14427 41605
rect 14369 41565 14381 41599
rect 14415 41565 14427 41599
rect 14369 41559 14427 41565
rect 14461 41599 14519 41605
rect 14461 41565 14473 41599
rect 14507 41565 14519 41599
rect 14461 41559 14519 41565
rect 12434 41488 12440 41540
rect 12492 41528 12498 41540
rect 12805 41531 12863 41537
rect 12805 41528 12817 41531
rect 12492 41500 12817 41528
rect 12492 41488 12498 41500
rect 12805 41497 12817 41500
rect 12851 41497 12863 41531
rect 12986 41528 12992 41540
rect 12947 41500 12992 41528
rect 12805 41491 12863 41497
rect 12986 41488 12992 41500
rect 13044 41488 13050 41540
rect 14384 41528 14412 41559
rect 14550 41556 14556 41608
rect 14608 41596 14614 41608
rect 14608 41568 14653 41596
rect 14608 41556 14614 41568
rect 14734 41556 14740 41608
rect 14792 41596 14798 41608
rect 14792 41568 14837 41596
rect 14792 41556 14798 41568
rect 15396 41528 15424 41636
rect 15856 41636 16988 41664
rect 15856 41605 15884 41636
rect 15841 41599 15899 41605
rect 15841 41565 15853 41599
rect 15887 41565 15899 41599
rect 16022 41596 16028 41608
rect 15983 41568 16028 41596
rect 15841 41559 15899 41565
rect 16022 41556 16028 41568
rect 16080 41556 16086 41608
rect 16117 41599 16175 41605
rect 16117 41565 16129 41599
rect 16163 41565 16175 41599
rect 16117 41559 16175 41565
rect 16209 41599 16267 41605
rect 16209 41565 16221 41599
rect 16255 41596 16267 41599
rect 16574 41596 16580 41608
rect 16255 41568 16580 41596
rect 16255 41565 16267 41568
rect 16209 41559 16267 41565
rect 16132 41528 16160 41559
rect 16574 41556 16580 41568
rect 16632 41556 16638 41608
rect 16960 41605 16988 41636
rect 18690 41624 18696 41676
rect 18748 41664 18754 41676
rect 26050 41664 26056 41676
rect 18748 41636 26056 41664
rect 18748 41624 18754 41636
rect 26050 41624 26056 41636
rect 26108 41624 26114 41676
rect 16945 41599 17003 41605
rect 16945 41565 16957 41599
rect 16991 41565 17003 41599
rect 17126 41596 17132 41608
rect 17087 41568 17132 41596
rect 16945 41559 17003 41565
rect 17126 41556 17132 41568
rect 17184 41556 17190 41608
rect 17221 41599 17279 41605
rect 17221 41565 17233 41599
rect 17267 41565 17279 41599
rect 17221 41559 17279 41565
rect 17236 41528 17264 41559
rect 17310 41556 17316 41608
rect 17368 41596 17374 41608
rect 19429 41599 19487 41605
rect 17368 41568 17413 41596
rect 17368 41556 17374 41568
rect 19429 41565 19441 41599
rect 19475 41596 19487 41599
rect 19978 41596 19984 41608
rect 19475 41568 19984 41596
rect 19475 41565 19487 41568
rect 19429 41559 19487 41565
rect 19978 41556 19984 41568
rect 20036 41556 20042 41608
rect 58158 41596 58164 41608
rect 58119 41568 58164 41596
rect 58158 41556 58164 41568
rect 58216 41556 58222 41608
rect 14384 41500 15332 41528
rect 15396 41500 17264 41528
rect 15304 41472 15332 41500
rect 17954 41488 17960 41540
rect 18012 41528 18018 41540
rect 19245 41531 19303 41537
rect 19245 41528 19257 41531
rect 18012 41500 19257 41528
rect 18012 41488 18018 41500
rect 19245 41497 19257 41500
rect 19291 41497 19303 41531
rect 19245 41491 19303 41497
rect 19613 41531 19671 41537
rect 19613 41497 19625 41531
rect 19659 41528 19671 41531
rect 20254 41528 20260 41540
rect 19659 41500 20260 41528
rect 19659 41497 19671 41500
rect 19613 41491 19671 41497
rect 20254 41488 20260 41500
rect 20312 41488 20318 41540
rect 9858 41420 9864 41472
rect 9916 41460 9922 41472
rect 10321 41463 10379 41469
rect 10321 41460 10333 41463
rect 9916 41432 10333 41460
rect 9916 41420 9922 41432
rect 10321 41429 10333 41432
rect 10367 41429 10379 41463
rect 10321 41423 10379 41429
rect 12621 41463 12679 41469
rect 12621 41429 12633 41463
rect 12667 41460 12679 41463
rect 13078 41460 13084 41472
rect 12667 41432 13084 41460
rect 12667 41429 12679 41432
rect 12621 41423 12679 41429
rect 13078 41420 13084 41432
rect 13136 41420 13142 41472
rect 13538 41460 13544 41472
rect 13499 41432 13544 41460
rect 13538 41420 13544 41432
rect 13596 41420 13602 41472
rect 14090 41460 14096 41472
rect 14051 41432 14096 41460
rect 14090 41420 14096 41432
rect 14148 41420 14154 41472
rect 15286 41460 15292 41472
rect 15247 41432 15292 41460
rect 15286 41420 15292 41432
rect 15344 41420 15350 41472
rect 16390 41420 16396 41472
rect 16448 41460 16454 41472
rect 16485 41463 16543 41469
rect 16485 41460 16497 41463
rect 16448 41432 16497 41460
rect 16448 41420 16454 41432
rect 16485 41429 16497 41432
rect 16531 41429 16543 41463
rect 16485 41423 16543 41429
rect 17589 41463 17647 41469
rect 17589 41429 17601 41463
rect 17635 41460 17647 41463
rect 17770 41460 17776 41472
rect 17635 41432 17776 41460
rect 17635 41429 17647 41432
rect 17589 41423 17647 41429
rect 17770 41420 17776 41432
rect 17828 41420 17834 41472
rect 19426 41420 19432 41472
rect 19484 41460 19490 41472
rect 20073 41463 20131 41469
rect 20073 41460 20085 41463
rect 19484 41432 20085 41460
rect 19484 41420 19490 41432
rect 20073 41429 20085 41432
rect 20119 41429 20131 41463
rect 20073 41423 20131 41429
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 12986 41216 12992 41268
rect 13044 41256 13050 41268
rect 13044 41228 15240 41256
rect 13044 41216 13050 41228
rect 6546 41148 6552 41200
rect 6604 41188 6610 41200
rect 10229 41191 10287 41197
rect 6604 41160 6773 41188
rect 6604 41148 6610 41160
rect 6745 41132 6773 41160
rect 10229 41157 10241 41191
rect 10275 41188 10287 41191
rect 11054 41188 11060 41200
rect 10275 41160 11060 41188
rect 10275 41157 10287 41160
rect 10229 41151 10287 41157
rect 11054 41148 11060 41160
rect 11112 41148 11118 41200
rect 15212 41197 15240 41228
rect 16574 41216 16580 41268
rect 16632 41256 16638 41268
rect 17037 41259 17095 41265
rect 16632 41228 16988 41256
rect 16632 41216 16638 41228
rect 15197 41191 15255 41197
rect 13280 41160 14412 41188
rect 6641 41123 6699 41129
rect 6641 41089 6653 41123
rect 6687 41089 6699 41123
rect 6641 41083 6699 41089
rect 6730 41126 6788 41132
rect 6730 41092 6742 41126
rect 6776 41092 6788 41126
rect 6730 41086 6788 41092
rect 6846 41123 6904 41129
rect 6846 41089 6858 41123
rect 6892 41120 6904 41123
rect 7009 41123 7067 41129
rect 6892 41092 6960 41120
rect 6892 41089 6904 41092
rect 6846 41083 6904 41089
rect 6656 40984 6684 41083
rect 6932 41052 6960 41092
rect 7009 41089 7021 41123
rect 7055 41120 7067 41123
rect 7650 41120 7656 41132
rect 7055 41092 7656 41120
rect 7055 41089 7067 41092
rect 7009 41083 7067 41089
rect 7650 41080 7656 41092
rect 7708 41080 7714 41132
rect 10413 41123 10471 41129
rect 10413 41089 10425 41123
rect 10459 41120 10471 41123
rect 10594 41120 10600 41132
rect 10459 41092 10600 41120
rect 10459 41089 10471 41092
rect 10413 41083 10471 41089
rect 10594 41080 10600 41092
rect 10652 41080 10658 41132
rect 12897 41123 12955 41129
rect 12897 41089 12909 41123
rect 12943 41089 12955 41123
rect 12897 41083 12955 41089
rect 12989 41123 13047 41129
rect 12989 41089 13001 41123
rect 13035 41089 13047 41123
rect 12989 41083 13047 41089
rect 7098 41052 7104 41064
rect 6932 41024 7104 41052
rect 7098 41012 7104 41024
rect 7156 41012 7162 41064
rect 12912 40984 12940 41083
rect 13004 41052 13032 41083
rect 13078 41080 13084 41132
rect 13136 41120 13142 41132
rect 13280 41129 13308 41160
rect 14384 41132 14412 41160
rect 15197 41157 15209 41191
rect 15243 41188 15255 41191
rect 16666 41188 16672 41200
rect 15243 41160 16672 41188
rect 15243 41157 15255 41160
rect 15197 41151 15255 41157
rect 16666 41148 16672 41160
rect 16724 41148 16730 41200
rect 16960 41188 16988 41228
rect 17037 41225 17049 41259
rect 17083 41256 17095 41259
rect 17126 41256 17132 41268
rect 17083 41228 17132 41256
rect 17083 41225 17095 41228
rect 17037 41219 17095 41225
rect 17126 41216 17132 41228
rect 17184 41216 17190 41268
rect 20809 41259 20867 41265
rect 20809 41256 20821 41259
rect 17880 41228 20821 41256
rect 17880 41188 17908 41228
rect 16960 41160 17908 41188
rect 18708 41160 19196 41188
rect 13265 41123 13323 41129
rect 13136 41092 13181 41120
rect 13136 41080 13142 41092
rect 13265 41089 13277 41123
rect 13311 41089 13323 41123
rect 13265 41083 13323 41089
rect 14001 41123 14059 41129
rect 14001 41089 14013 41123
rect 14047 41089 14059 41123
rect 14001 41083 14059 41089
rect 14093 41123 14151 41129
rect 14093 41089 14105 41123
rect 14139 41089 14151 41123
rect 14093 41083 14151 41089
rect 14185 41123 14243 41129
rect 14185 41089 14197 41123
rect 14231 41089 14243 41123
rect 14185 41083 14243 41089
rect 13906 41052 13912 41064
rect 13004 41024 13912 41052
rect 13906 41012 13912 41024
rect 13964 41012 13970 41064
rect 13538 40984 13544 40996
rect 6656 40956 7604 40984
rect 12912 40956 13544 40984
rect 7576 40928 7604 40956
rect 13538 40944 13544 40956
rect 13596 40944 13602 40996
rect 6362 40916 6368 40928
rect 6323 40888 6368 40916
rect 6362 40876 6368 40888
rect 6420 40876 6426 40928
rect 7558 40916 7564 40928
rect 7519 40888 7564 40916
rect 7558 40876 7564 40888
rect 7616 40876 7622 40928
rect 10410 40876 10416 40928
rect 10468 40916 10474 40928
rect 10597 40919 10655 40925
rect 10597 40916 10609 40919
rect 10468 40888 10609 40916
rect 10468 40876 10474 40888
rect 10597 40885 10609 40888
rect 10643 40885 10655 40919
rect 12618 40916 12624 40928
rect 12579 40888 12624 40916
rect 10597 40879 10655 40885
rect 12618 40876 12624 40888
rect 12676 40876 12682 40928
rect 13722 40916 13728 40928
rect 13683 40888 13728 40916
rect 13722 40876 13728 40888
rect 13780 40876 13786 40928
rect 14016 40916 14044 41083
rect 14108 40984 14136 41083
rect 14200 41052 14228 41083
rect 14366 41080 14372 41132
rect 14424 41120 14430 41132
rect 14734 41120 14740 41132
rect 14424 41092 14740 41120
rect 14424 41080 14430 41092
rect 14734 41080 14740 41092
rect 14792 41080 14798 41132
rect 15010 41120 15016 41132
rect 14971 41092 15016 41120
rect 15010 41080 15016 41092
rect 15068 41080 15074 41132
rect 16853 41123 16911 41129
rect 16853 41089 16865 41123
rect 16899 41120 16911 41123
rect 17034 41120 17040 41132
rect 16899 41092 17040 41120
rect 16899 41089 16911 41092
rect 16853 41083 16911 41089
rect 17034 41080 17040 41092
rect 17092 41080 17098 41132
rect 17773 41123 17831 41129
rect 17773 41089 17785 41123
rect 17819 41089 17831 41123
rect 17954 41120 17960 41132
rect 17915 41092 17960 41120
rect 17773 41083 17831 41089
rect 14829 41055 14887 41061
rect 14829 41052 14841 41055
rect 14200 41024 14841 41052
rect 14829 41021 14841 41024
rect 14875 41021 14887 41055
rect 14829 41015 14887 41021
rect 14182 40984 14188 40996
rect 14108 40956 14188 40984
rect 14182 40944 14188 40956
rect 14240 40944 14246 40996
rect 17788 40984 17816 41083
rect 17954 41080 17960 41092
rect 18012 41080 18018 41132
rect 18049 41123 18107 41129
rect 18049 41089 18061 41123
rect 18095 41089 18107 41123
rect 18049 41083 18107 41089
rect 18141 41123 18199 41129
rect 18141 41089 18153 41123
rect 18187 41120 18199 41123
rect 18598 41120 18604 41132
rect 18187 41092 18604 41120
rect 18187 41089 18199 41092
rect 18141 41083 18199 41089
rect 18064 41052 18092 41083
rect 18598 41080 18604 41092
rect 18656 41080 18662 41132
rect 18708 41064 18736 41160
rect 19168 41132 19196 41160
rect 18877 41123 18935 41129
rect 18877 41089 18889 41123
rect 18923 41089 18935 41123
rect 19061 41123 19119 41129
rect 19061 41120 19073 41123
rect 18877 41083 18935 41089
rect 18984 41092 19073 41120
rect 18690 41052 18696 41064
rect 18064 41024 18696 41052
rect 18690 41012 18696 41024
rect 18748 41012 18754 41064
rect 18598 40984 18604 40996
rect 17788 40956 18604 40984
rect 18598 40944 18604 40956
rect 18656 40984 18662 40996
rect 18892 40984 18920 41083
rect 18656 40956 18920 40984
rect 18656 40944 18662 40956
rect 15657 40919 15715 40925
rect 15657 40916 15669 40919
rect 14016 40888 15669 40916
rect 15657 40885 15669 40888
rect 15703 40916 15715 40919
rect 17678 40916 17684 40928
rect 15703 40888 17684 40916
rect 15703 40885 15715 40888
rect 15657 40879 15715 40885
rect 17678 40876 17684 40888
rect 17736 40876 17742 40928
rect 18414 40916 18420 40928
rect 18375 40888 18420 40916
rect 18414 40876 18420 40888
rect 18472 40876 18478 40928
rect 18984 40916 19012 41092
rect 19061 41089 19073 41092
rect 19107 41089 19119 41123
rect 19061 41083 19119 41089
rect 19153 41126 19211 41132
rect 19260 41129 19288 41228
rect 20809 41225 20821 41228
rect 20855 41256 20867 41259
rect 24118 41256 24124 41268
rect 20855 41228 24124 41256
rect 20855 41225 20867 41228
rect 20809 41219 20867 41225
rect 24118 41216 24124 41228
rect 24176 41216 24182 41268
rect 20165 41191 20223 41197
rect 20165 41157 20177 41191
rect 20211 41188 20223 41191
rect 20622 41188 20628 41200
rect 20211 41160 20628 41188
rect 20211 41157 20223 41160
rect 20165 41151 20223 41157
rect 20622 41148 20628 41160
rect 20680 41148 20686 41200
rect 19153 41092 19165 41126
rect 19199 41092 19211 41126
rect 19153 41086 19211 41092
rect 19245 41123 19303 41129
rect 19245 41089 19257 41123
rect 19291 41089 19303 41123
rect 19245 41083 19303 41089
rect 20070 41080 20076 41132
rect 20128 41120 20134 41132
rect 20254 41120 20260 41132
rect 20128 41092 20260 41120
rect 20128 41080 20134 41092
rect 20254 41080 20260 41092
rect 20312 41120 20318 41132
rect 20349 41123 20407 41129
rect 20349 41120 20361 41123
rect 20312 41092 20361 41120
rect 20312 41080 20318 41092
rect 20349 41089 20361 41092
rect 20395 41089 20407 41123
rect 20349 41083 20407 41089
rect 19981 41055 20039 41061
rect 19981 41052 19993 41055
rect 19260 41024 19993 41052
rect 19260 40916 19288 41024
rect 19981 41021 19993 41024
rect 20027 41021 20039 41055
rect 19981 41015 20039 41021
rect 22649 40987 22707 40993
rect 22649 40953 22661 40987
rect 22695 40984 22707 40987
rect 23750 40984 23756 40996
rect 22695 40956 23756 40984
rect 22695 40953 22707 40956
rect 22649 40947 22707 40953
rect 19518 40916 19524 40928
rect 18984 40888 19288 40916
rect 19479 40888 19524 40916
rect 19518 40876 19524 40888
rect 19576 40876 19582 40928
rect 22094 40876 22100 40928
rect 22152 40916 22158 40928
rect 22664 40916 22692 40947
rect 23750 40944 23756 40956
rect 23808 40944 23814 40996
rect 22152 40888 22692 40916
rect 22152 40876 22158 40888
rect 23014 40876 23020 40928
rect 23072 40916 23078 40928
rect 23201 40919 23259 40925
rect 23201 40916 23213 40919
rect 23072 40888 23213 40916
rect 23072 40876 23078 40888
rect 23201 40885 23213 40888
rect 23247 40885 23259 40919
rect 23201 40879 23259 40885
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 9858 40672 9864 40724
rect 9916 40712 9922 40724
rect 13541 40715 13599 40721
rect 9916 40684 13492 40712
rect 9916 40672 9922 40684
rect 13464 40644 13492 40684
rect 13541 40681 13553 40715
rect 13587 40712 13599 40715
rect 14550 40712 14556 40724
rect 13587 40684 14556 40712
rect 13587 40681 13599 40684
rect 13541 40675 13599 40681
rect 14550 40672 14556 40684
rect 14608 40672 14614 40724
rect 18598 40712 18604 40724
rect 18559 40684 18604 40712
rect 18598 40672 18604 40684
rect 18656 40672 18662 40724
rect 15194 40644 15200 40656
rect 13464 40616 15200 40644
rect 15194 40604 15200 40616
rect 15252 40604 15258 40656
rect 9214 40536 9220 40588
rect 9272 40576 9278 40588
rect 10689 40579 10747 40585
rect 10689 40576 10701 40579
rect 9272 40548 10701 40576
rect 9272 40536 9278 40548
rect 10689 40545 10701 40548
rect 10735 40545 10747 40579
rect 10689 40539 10747 40545
rect 13906 40536 13912 40588
rect 13964 40576 13970 40588
rect 14182 40576 14188 40588
rect 13964 40548 14188 40576
rect 13964 40536 13970 40548
rect 14182 40536 14188 40548
rect 14240 40536 14246 40588
rect 14366 40576 14372 40588
rect 14327 40548 14372 40576
rect 14366 40536 14372 40548
rect 14424 40536 14430 40588
rect 3789 40511 3847 40517
rect 3789 40477 3801 40511
rect 3835 40508 3847 40511
rect 6086 40508 6092 40520
rect 3835 40480 5396 40508
rect 6047 40480 6092 40508
rect 3835 40477 3847 40480
rect 3789 40471 3847 40477
rect 3970 40440 3976 40452
rect 3931 40412 3976 40440
rect 3970 40400 3976 40412
rect 4028 40400 4034 40452
rect 5368 40440 5396 40480
rect 6086 40468 6092 40480
rect 6144 40468 6150 40520
rect 6362 40517 6368 40520
rect 6356 40508 6368 40517
rect 6323 40480 6368 40508
rect 6356 40471 6368 40480
rect 6362 40468 6368 40471
rect 6420 40468 6426 40520
rect 9858 40508 9864 40520
rect 9819 40480 9864 40508
rect 9858 40468 9864 40480
rect 9916 40468 9922 40520
rect 9950 40508 10008 40514
rect 9950 40474 9962 40508
rect 9996 40474 10008 40508
rect 9950 40468 10008 40474
rect 10042 40468 10048 40520
rect 10100 40508 10106 40520
rect 10229 40511 10287 40517
rect 10100 40480 10145 40508
rect 10100 40468 10106 40480
rect 10229 40477 10241 40511
rect 10275 40508 10287 40511
rect 10502 40508 10508 40520
rect 10275 40480 10508 40508
rect 10275 40477 10287 40480
rect 10229 40471 10287 40477
rect 10502 40468 10508 40480
rect 10560 40468 10566 40520
rect 10956 40511 11014 40517
rect 10956 40477 10968 40511
rect 11002 40508 11014 40511
rect 12618 40508 12624 40520
rect 11002 40480 12624 40508
rect 11002 40477 11014 40480
rect 10956 40471 11014 40477
rect 12618 40468 12624 40480
rect 12676 40468 12682 40520
rect 12802 40468 12808 40520
rect 12860 40508 12866 40520
rect 13357 40511 13415 40517
rect 13357 40508 13369 40511
rect 12860 40480 13369 40508
rect 12860 40468 12866 40480
rect 13357 40477 13369 40480
rect 13403 40477 13415 40511
rect 13357 40471 13415 40477
rect 13814 40468 13820 40520
rect 13872 40508 13878 40520
rect 14093 40511 14151 40517
rect 14093 40508 14105 40511
rect 13872 40480 14105 40508
rect 13872 40468 13878 40480
rect 14093 40477 14105 40480
rect 14139 40477 14151 40511
rect 14093 40471 14151 40477
rect 15378 40468 15384 40520
rect 15436 40508 15442 40520
rect 16390 40517 16396 40520
rect 16117 40511 16175 40517
rect 16117 40508 16129 40511
rect 15436 40480 16129 40508
rect 15436 40468 15442 40480
rect 16117 40477 16129 40480
rect 16163 40477 16175 40511
rect 16117 40471 16175 40477
rect 16384 40471 16396 40517
rect 16448 40508 16454 40520
rect 16448 40480 16484 40508
rect 16390 40468 16396 40471
rect 16448 40468 16454 40480
rect 18322 40468 18328 40520
rect 18380 40508 18386 40520
rect 19518 40517 19524 40520
rect 19245 40511 19303 40517
rect 19245 40508 19257 40511
rect 18380 40480 19257 40508
rect 18380 40468 18386 40480
rect 19245 40477 19257 40480
rect 19291 40477 19303 40511
rect 19512 40508 19524 40517
rect 19479 40480 19524 40508
rect 19245 40471 19303 40477
rect 19512 40471 19524 40480
rect 19518 40468 19524 40471
rect 19576 40468 19582 40520
rect 22094 40508 22100 40520
rect 22055 40480 22100 40508
rect 22094 40468 22100 40480
rect 22152 40468 22158 40520
rect 22189 40511 22247 40517
rect 22189 40477 22201 40511
rect 22235 40477 22247 40511
rect 22189 40471 22247 40477
rect 9965 40440 9993 40468
rect 10134 40440 10140 40452
rect 5368 40412 6408 40440
rect 9965 40412 10140 40440
rect 6380 40384 6408 40412
rect 10134 40400 10140 40412
rect 10192 40400 10198 40452
rect 13078 40400 13084 40452
rect 13136 40440 13142 40452
rect 13173 40443 13231 40449
rect 13173 40440 13185 40443
rect 13136 40412 13185 40440
rect 13136 40400 13142 40412
rect 13173 40409 13185 40412
rect 13219 40409 13231 40443
rect 22112 40440 22140 40468
rect 13173 40403 13231 40409
rect 15304 40412 22140 40440
rect 22204 40440 22232 40471
rect 22278 40468 22284 40520
rect 22336 40508 22342 40520
rect 22336 40480 22381 40508
rect 22336 40468 22342 40480
rect 22462 40468 22468 40520
rect 22520 40508 22526 40520
rect 23201 40511 23259 40517
rect 22520 40480 22565 40508
rect 22520 40468 22526 40480
rect 23201 40477 23213 40511
rect 23247 40508 23259 40511
rect 23382 40508 23388 40520
rect 23247 40480 23388 40508
rect 23247 40477 23259 40480
rect 23201 40471 23259 40477
rect 23382 40468 23388 40480
rect 23440 40468 23446 40520
rect 27338 40508 27344 40520
rect 27299 40480 27344 40508
rect 27338 40468 27344 40480
rect 27396 40468 27402 40520
rect 31202 40508 31208 40520
rect 31163 40480 31208 40508
rect 31202 40468 31208 40480
rect 31260 40468 31266 40520
rect 58158 40508 58164 40520
rect 58119 40480 58164 40508
rect 58158 40468 58164 40480
rect 58216 40468 58222 40520
rect 22738 40440 22744 40452
rect 22204 40412 22744 40440
rect 4157 40375 4215 40381
rect 4157 40341 4169 40375
rect 4203 40372 4215 40375
rect 4614 40372 4620 40384
rect 4203 40344 4620 40372
rect 4203 40341 4215 40344
rect 4157 40335 4215 40341
rect 4614 40332 4620 40344
rect 4672 40332 4678 40384
rect 6362 40332 6368 40384
rect 6420 40332 6426 40384
rect 7469 40375 7527 40381
rect 7469 40341 7481 40375
rect 7515 40372 7527 40375
rect 7742 40372 7748 40384
rect 7515 40344 7748 40372
rect 7515 40341 7527 40344
rect 7469 40335 7527 40341
rect 7742 40332 7748 40344
rect 7800 40332 7806 40384
rect 9582 40372 9588 40384
rect 9543 40344 9588 40372
rect 9582 40332 9588 40344
rect 9640 40332 9646 40384
rect 12069 40375 12127 40381
rect 12069 40341 12081 40375
rect 12115 40372 12127 40375
rect 12434 40372 12440 40384
rect 12115 40344 12440 40372
rect 12115 40341 12127 40344
rect 12069 40335 12127 40341
rect 12434 40332 12440 40344
rect 12492 40332 12498 40384
rect 12618 40332 12624 40384
rect 12676 40372 12682 40384
rect 15102 40372 15108 40384
rect 12676 40344 15108 40372
rect 12676 40332 12682 40344
rect 15102 40332 15108 40344
rect 15160 40372 15166 40384
rect 15304 40372 15332 40412
rect 22738 40400 22744 40412
rect 22796 40400 22802 40452
rect 23017 40443 23075 40449
rect 23017 40409 23029 40443
rect 23063 40440 23075 40443
rect 23106 40440 23112 40452
rect 23063 40412 23112 40440
rect 23063 40409 23075 40412
rect 23017 40403 23075 40409
rect 23106 40400 23112 40412
rect 23164 40400 23170 40452
rect 27614 40449 27620 40452
rect 27608 40403 27620 40449
rect 27672 40440 27678 40452
rect 31478 40449 31484 40452
rect 27672 40412 27708 40440
rect 27614 40400 27620 40403
rect 27672 40400 27678 40412
rect 31472 40403 31484 40449
rect 31536 40440 31542 40452
rect 31536 40412 31572 40440
rect 31478 40400 31484 40403
rect 31536 40400 31542 40412
rect 15160 40344 15332 40372
rect 15160 40332 15166 40344
rect 16942 40332 16948 40384
rect 17000 40372 17006 40384
rect 17494 40372 17500 40384
rect 17000 40344 17500 40372
rect 17000 40332 17006 40344
rect 17494 40332 17500 40344
rect 17552 40332 17558 40384
rect 18598 40332 18604 40384
rect 18656 40372 18662 40384
rect 19426 40372 19432 40384
rect 18656 40344 19432 40372
rect 18656 40332 18662 40344
rect 19426 40332 19432 40344
rect 19484 40372 19490 40384
rect 20346 40372 20352 40384
rect 19484 40344 20352 40372
rect 19484 40332 19490 40344
rect 20346 40332 20352 40344
rect 20404 40332 20410 40384
rect 20622 40372 20628 40384
rect 20583 40344 20628 40372
rect 20622 40332 20628 40344
rect 20680 40332 20686 40384
rect 21821 40375 21879 40381
rect 21821 40341 21833 40375
rect 21867 40372 21879 40375
rect 22094 40372 22100 40384
rect 21867 40344 22100 40372
rect 21867 40341 21879 40344
rect 21821 40335 21879 40341
rect 22094 40332 22100 40344
rect 22152 40332 22158 40384
rect 23290 40332 23296 40384
rect 23348 40372 23354 40384
rect 23385 40375 23443 40381
rect 23385 40372 23397 40375
rect 23348 40344 23397 40372
rect 23348 40332 23354 40344
rect 23385 40341 23397 40344
rect 23431 40341 23443 40375
rect 28718 40372 28724 40384
rect 28679 40344 28724 40372
rect 23385 40335 23443 40341
rect 28718 40332 28724 40344
rect 28776 40332 28782 40384
rect 32030 40332 32036 40384
rect 32088 40372 32094 40384
rect 32585 40375 32643 40381
rect 32585 40372 32597 40375
rect 32088 40344 32597 40372
rect 32088 40332 32094 40344
rect 32585 40341 32597 40344
rect 32631 40341 32643 40375
rect 32585 40335 32643 40341
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 3510 40128 3516 40180
rect 3568 40168 3574 40180
rect 3970 40168 3976 40180
rect 3568 40140 3976 40168
rect 3568 40128 3574 40140
rect 3970 40128 3976 40140
rect 4028 40128 4034 40180
rect 7742 40168 7748 40180
rect 6748 40140 7748 40168
rect 6086 40060 6092 40112
rect 6144 40100 6150 40112
rect 6144 40072 6684 40100
rect 6144 40060 6150 40072
rect 2860 40035 2918 40041
rect 2860 40001 2872 40035
rect 2906 40032 2918 40035
rect 3786 40032 3792 40044
rect 2906 40004 3792 40032
rect 2906 40001 2918 40004
rect 2860 39995 2918 40001
rect 3786 39992 3792 40004
rect 3844 39992 3850 40044
rect 6362 39992 6368 40044
rect 6420 40032 6426 40044
rect 6549 40035 6607 40041
rect 6549 40032 6561 40035
rect 6420 40004 6561 40032
rect 6420 39992 6426 40004
rect 6549 40001 6561 40004
rect 6595 40001 6607 40035
rect 6549 39995 6607 40001
rect 2590 39964 2596 39976
rect 2551 39936 2596 39964
rect 2590 39924 2596 39936
rect 2648 39924 2654 39976
rect 6656 39964 6684 40072
rect 6748 40041 6776 40140
rect 7742 40128 7748 40140
rect 7800 40128 7806 40180
rect 8757 40171 8815 40177
rect 8757 40137 8769 40171
rect 8803 40168 8815 40171
rect 11238 40168 11244 40180
rect 8803 40140 11244 40168
rect 8803 40137 8815 40140
rect 8757 40131 8815 40137
rect 11238 40128 11244 40140
rect 11296 40128 11302 40180
rect 12161 40171 12219 40177
rect 12161 40168 12173 40171
rect 11348 40140 12173 40168
rect 6917 40103 6975 40109
rect 6917 40069 6929 40103
rect 6963 40100 6975 40103
rect 7098 40100 7104 40112
rect 6963 40072 7104 40100
rect 6963 40069 6975 40072
rect 6917 40063 6975 40069
rect 7098 40060 7104 40072
rect 7156 40060 7162 40112
rect 9214 40100 9220 40112
rect 7392 40072 9220 40100
rect 7392 40041 7420 40072
rect 9214 40060 9220 40072
rect 9272 40060 9278 40112
rect 9484 40103 9542 40109
rect 9484 40069 9496 40103
rect 9530 40100 9542 40103
rect 9582 40100 9588 40112
rect 9530 40072 9588 40100
rect 9530 40069 9542 40072
rect 9484 40063 9542 40069
rect 9582 40060 9588 40072
rect 9640 40060 9646 40112
rect 11348 40100 11376 40140
rect 12161 40137 12173 40140
rect 12207 40137 12219 40171
rect 12802 40168 12808 40180
rect 12763 40140 12808 40168
rect 12161 40131 12219 40137
rect 12802 40128 12808 40140
rect 12860 40128 12866 40180
rect 16669 40171 16727 40177
rect 16669 40137 16681 40171
rect 16715 40168 16727 40171
rect 17034 40168 17040 40180
rect 16715 40140 17040 40168
rect 16715 40137 16727 40140
rect 16669 40131 16727 40137
rect 17034 40128 17040 40140
rect 17092 40128 17098 40180
rect 19889 40171 19947 40177
rect 19889 40137 19901 40171
rect 19935 40168 19947 40171
rect 19978 40168 19984 40180
rect 19935 40140 19984 40168
rect 19935 40137 19947 40140
rect 19889 40131 19947 40137
rect 19978 40128 19984 40140
rect 20036 40128 20042 40180
rect 27614 40168 27620 40180
rect 27575 40140 27620 40168
rect 27614 40128 27620 40140
rect 27672 40128 27678 40180
rect 12618 40100 12624 40112
rect 10428 40072 11376 40100
rect 11900 40072 12624 40100
rect 6733 40035 6791 40041
rect 6733 40001 6745 40035
rect 6779 40001 6791 40035
rect 6733 39995 6791 40001
rect 7377 40035 7435 40041
rect 7377 40001 7389 40035
rect 7423 40001 7435 40035
rect 7377 39995 7435 40001
rect 7644 40035 7702 40041
rect 7644 40001 7656 40035
rect 7690 40032 7702 40035
rect 10428 40032 10456 40072
rect 7690 40004 10456 40032
rect 7690 40001 7702 40004
rect 7644 39995 7702 40001
rect 7392 39964 7420 39995
rect 10502 39992 10508 40044
rect 10560 40032 10566 40044
rect 10686 40032 10692 40044
rect 10560 40004 10692 40032
rect 10560 39992 10566 40004
rect 10686 39992 10692 40004
rect 10744 40032 10750 40044
rect 11517 40035 11575 40041
rect 11517 40032 11529 40035
rect 10744 40004 11529 40032
rect 10744 39992 10750 40004
rect 11517 40001 11529 40004
rect 11563 40001 11575 40035
rect 11698 40032 11704 40044
rect 11659 40004 11704 40032
rect 11517 39995 11575 40001
rect 11698 39992 11704 40004
rect 11756 39992 11762 40044
rect 11900 40041 11928 40072
rect 12618 40060 12624 40072
rect 12676 40060 12682 40112
rect 18414 40060 18420 40112
rect 18472 40100 18478 40112
rect 18754 40103 18812 40109
rect 18754 40100 18766 40103
rect 18472 40072 18766 40100
rect 18472 40060 18478 40072
rect 18754 40069 18766 40072
rect 18800 40069 18812 40103
rect 18754 40063 18812 40069
rect 20901 40103 20959 40109
rect 20901 40069 20913 40103
rect 20947 40100 20959 40103
rect 21450 40100 21456 40112
rect 20947 40072 21456 40100
rect 20947 40069 20959 40072
rect 20901 40063 20959 40069
rect 21450 40060 21456 40072
rect 21508 40060 21514 40112
rect 28718 40060 28724 40112
rect 28776 40100 28782 40112
rect 28905 40103 28963 40109
rect 28905 40100 28917 40103
rect 28776 40072 28917 40100
rect 28776 40060 28782 40072
rect 28905 40069 28917 40072
rect 28951 40069 28963 40103
rect 29086 40100 29092 40112
rect 29047 40072 29092 40100
rect 28905 40063 28963 40069
rect 29086 40060 29092 40072
rect 29144 40060 29150 40112
rect 11796 40035 11854 40041
rect 11796 40001 11808 40035
rect 11842 40001 11854 40035
rect 11796 39995 11854 40001
rect 11885 40035 11943 40041
rect 11885 40001 11897 40035
rect 11931 40001 11943 40035
rect 11885 39995 11943 40001
rect 13929 40035 13987 40041
rect 13929 40001 13941 40035
rect 13975 40032 13987 40035
rect 14090 40032 14096 40044
rect 13975 40004 14096 40032
rect 13975 40001 13987 40004
rect 13929 39995 13987 40001
rect 9214 39964 9220 39976
rect 6656 39936 7420 39964
rect 9175 39936 9220 39964
rect 9214 39924 9220 39936
rect 9272 39924 9278 39976
rect 11808 39896 11836 39995
rect 14090 39992 14096 40004
rect 14148 39992 14154 40044
rect 17770 39992 17776 40044
rect 17828 40041 17834 40044
rect 17828 40032 17840 40041
rect 17828 40004 17873 40032
rect 17828 39995 17840 40004
rect 17828 39992 17834 39995
rect 20990 39992 20996 40044
rect 21048 40032 21054 40044
rect 21085 40035 21143 40041
rect 21085 40032 21097 40035
rect 21048 40004 21097 40032
rect 21048 39992 21054 40004
rect 21085 40001 21097 40004
rect 21131 40001 21143 40035
rect 21085 39995 21143 40001
rect 21269 40035 21327 40041
rect 21269 40001 21281 40035
rect 21315 40032 21327 40035
rect 22278 40032 22284 40044
rect 21315 40004 22284 40032
rect 21315 40001 21327 40004
rect 21269 39995 21327 40001
rect 22278 39992 22284 40004
rect 22336 39992 22342 40044
rect 22462 40032 22468 40044
rect 22423 40004 22468 40032
rect 22462 39992 22468 40004
rect 22520 39992 22526 40044
rect 22646 40032 22652 40044
rect 22607 40004 22652 40032
rect 22646 39992 22652 40004
rect 22704 39992 22710 40044
rect 22738 39992 22744 40044
rect 22796 40032 22802 40044
rect 22879 40035 22937 40041
rect 22796 40004 22841 40032
rect 22796 39992 22802 40004
rect 22879 40001 22891 40035
rect 22925 40032 22937 40035
rect 23014 40032 23020 40044
rect 22925 40004 23020 40032
rect 22925 40001 22937 40004
rect 22879 39995 22937 40001
rect 23014 39992 23020 40004
rect 23072 39992 23078 40044
rect 24682 40035 24740 40041
rect 24682 40032 24694 40035
rect 23124 40004 24694 40032
rect 14185 39967 14243 39973
rect 14185 39933 14197 39967
rect 14231 39964 14243 39967
rect 15378 39964 15384 39976
rect 14231 39936 15384 39964
rect 14231 39933 14243 39936
rect 14185 39927 14243 39933
rect 15378 39924 15384 39936
rect 15436 39924 15442 39976
rect 18049 39967 18107 39973
rect 18049 39933 18061 39967
rect 18095 39964 18107 39967
rect 18322 39964 18328 39976
rect 18095 39936 18328 39964
rect 18095 39933 18107 39936
rect 18049 39927 18107 39933
rect 10152 39868 11836 39896
rect 10152 39840 10180 39868
rect 10134 39788 10140 39840
rect 10192 39788 10198 39840
rect 10502 39788 10508 39840
rect 10560 39828 10566 39840
rect 10597 39831 10655 39837
rect 10597 39828 10609 39831
rect 10560 39800 10609 39828
rect 10560 39788 10566 39800
rect 10597 39797 10609 39800
rect 10643 39797 10655 39831
rect 10597 39791 10655 39797
rect 13814 39788 13820 39840
rect 13872 39828 13878 39840
rect 14645 39831 14703 39837
rect 14645 39828 14657 39831
rect 13872 39800 14657 39828
rect 13872 39788 13878 39800
rect 14645 39797 14657 39800
rect 14691 39797 14703 39831
rect 14645 39791 14703 39797
rect 15378 39788 15384 39840
rect 15436 39828 15442 39840
rect 18064 39828 18092 39927
rect 18322 39924 18328 39936
rect 18380 39964 18386 39976
rect 23124 39973 23152 40004
rect 24682 40001 24694 40004
rect 24728 40001 24740 40035
rect 24682 39995 24740 40001
rect 27062 39992 27068 40044
rect 27120 40032 27126 40044
rect 27847 40035 27905 40041
rect 27847 40032 27859 40035
rect 27120 40004 27859 40032
rect 27120 39992 27126 40004
rect 27847 40001 27859 40004
rect 27893 40001 27905 40035
rect 27982 40032 27988 40044
rect 27943 40004 27988 40032
rect 27847 39995 27905 40001
rect 27982 39992 27988 40004
rect 28040 39992 28046 40044
rect 28098 40035 28156 40041
rect 28098 40032 28110 40035
rect 28097 40001 28110 40032
rect 28144 40001 28156 40035
rect 28258 40032 28264 40044
rect 28219 40004 28264 40032
rect 28097 39995 28156 40001
rect 18509 39967 18567 39973
rect 18509 39964 18521 39967
rect 18380 39936 18521 39964
rect 18380 39924 18386 39936
rect 18509 39933 18521 39936
rect 18555 39933 18567 39967
rect 18509 39927 18567 39933
rect 23109 39967 23167 39973
rect 23109 39933 23121 39967
rect 23155 39933 23167 39967
rect 23109 39927 23167 39933
rect 24949 39967 25007 39973
rect 24949 39933 24961 39967
rect 24995 39933 25007 39967
rect 28097 39964 28125 39995
rect 28258 39992 28264 40004
rect 28316 39992 28322 40044
rect 28721 39967 28779 39973
rect 28721 39964 28733 39967
rect 28097 39936 28733 39964
rect 24949 39927 25007 39933
rect 28721 39933 28733 39936
rect 28767 39933 28779 39967
rect 28721 39927 28779 39933
rect 23566 39828 23572 39840
rect 15436 39800 18092 39828
rect 23527 39800 23572 39828
rect 15436 39788 15442 39800
rect 23566 39788 23572 39800
rect 23624 39788 23630 39840
rect 24762 39788 24768 39840
rect 24820 39828 24826 39840
rect 24964 39828 24992 39927
rect 27062 39828 27068 39840
rect 24820 39800 24992 39828
rect 27023 39800 27068 39828
rect 24820 39788 24826 39800
rect 27062 39788 27068 39800
rect 27120 39788 27126 39840
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 3786 39624 3792 39636
rect 3747 39596 3792 39624
rect 3786 39584 3792 39596
rect 3844 39584 3850 39636
rect 11425 39627 11483 39633
rect 3988 39596 5580 39624
rect 2590 39448 2596 39500
rect 2648 39488 2654 39500
rect 3988 39488 4016 39596
rect 4893 39559 4951 39565
rect 4893 39556 4905 39559
rect 2648 39460 4016 39488
rect 4080 39528 4905 39556
rect 2648 39448 2654 39460
rect 4080 39429 4108 39528
rect 4893 39525 4905 39528
rect 4939 39556 4951 39559
rect 5258 39556 5264 39568
rect 4939 39528 5264 39556
rect 4939 39525 4951 39528
rect 4893 39519 4951 39525
rect 5258 39516 5264 39528
rect 5316 39516 5322 39568
rect 4614 39488 4620 39500
rect 4264 39460 4620 39488
rect 4264 39429 4292 39460
rect 4614 39448 4620 39460
rect 4672 39448 4678 39500
rect 5552 39497 5580 39596
rect 11425 39593 11437 39627
rect 11471 39624 11483 39627
rect 11698 39624 11704 39636
rect 11471 39596 11704 39624
rect 11471 39593 11483 39596
rect 11425 39587 11483 39593
rect 11698 39584 11704 39596
rect 11756 39584 11762 39636
rect 12161 39627 12219 39633
rect 12161 39593 12173 39627
rect 12207 39624 12219 39627
rect 14090 39624 14096 39636
rect 12207 39596 14096 39624
rect 12207 39593 12219 39596
rect 12161 39587 12219 39593
rect 14090 39584 14096 39596
rect 14148 39624 14154 39636
rect 15010 39624 15016 39636
rect 14148 39596 15016 39624
rect 14148 39584 14154 39596
rect 15010 39584 15016 39596
rect 15068 39584 15074 39636
rect 15194 39584 15200 39636
rect 15252 39624 15258 39636
rect 16298 39624 16304 39636
rect 15252 39596 16304 39624
rect 15252 39584 15258 39596
rect 16298 39584 16304 39596
rect 16356 39624 16362 39636
rect 23014 39624 23020 39636
rect 16356 39596 23020 39624
rect 16356 39584 16362 39596
rect 23014 39584 23020 39596
rect 23072 39624 23078 39636
rect 23474 39624 23480 39636
rect 23072 39596 23480 39624
rect 23072 39584 23078 39596
rect 23474 39584 23480 39596
rect 23532 39584 23538 39636
rect 31478 39624 31484 39636
rect 31439 39596 31484 39624
rect 31478 39584 31484 39596
rect 31536 39584 31542 39636
rect 32309 39559 32367 39565
rect 32309 39556 32321 39559
rect 30944 39528 32321 39556
rect 5537 39491 5595 39497
rect 5537 39457 5549 39491
rect 5583 39457 5595 39491
rect 5537 39451 5595 39457
rect 13541 39491 13599 39497
rect 13541 39457 13553 39491
rect 13587 39488 13599 39491
rect 15378 39488 15384 39500
rect 13587 39460 15384 39488
rect 13587 39457 13599 39460
rect 13541 39451 13599 39457
rect 15378 39448 15384 39460
rect 15436 39448 15442 39500
rect 22373 39491 22431 39497
rect 22373 39457 22385 39491
rect 22419 39488 22431 39491
rect 30944 39488 30972 39528
rect 32309 39525 32321 39528
rect 32355 39525 32367 39559
rect 32309 39519 32367 39525
rect 22419 39460 24440 39488
rect 30944 39460 31064 39488
rect 22419 39457 22431 39460
rect 22373 39451 22431 39457
rect 4065 39423 4123 39429
rect 4065 39389 4077 39423
rect 4111 39389 4123 39423
rect 4065 39383 4123 39389
rect 4157 39423 4215 39429
rect 4157 39389 4169 39423
rect 4203 39389 4215 39423
rect 4157 39383 4215 39389
rect 4249 39423 4307 39429
rect 4249 39389 4261 39423
rect 4295 39389 4307 39423
rect 4249 39383 4307 39389
rect 4433 39423 4491 39429
rect 4433 39389 4445 39423
rect 4479 39420 4491 39423
rect 4890 39420 4896 39432
rect 4479 39392 4896 39420
rect 4479 39389 4491 39392
rect 4433 39383 4491 39389
rect 4172 39352 4200 39383
rect 4890 39380 4896 39392
rect 4948 39380 4954 39432
rect 7282 39380 7288 39432
rect 7340 39420 7346 39432
rect 7377 39423 7435 39429
rect 7377 39420 7389 39423
rect 7340 39392 7389 39420
rect 7340 39380 7346 39392
rect 7377 39389 7389 39392
rect 7423 39389 7435 39423
rect 7650 39420 7656 39432
rect 7611 39392 7656 39420
rect 7377 39383 7435 39389
rect 7650 39380 7656 39392
rect 7708 39380 7714 39432
rect 9214 39420 9220 39432
rect 9175 39392 9220 39420
rect 9214 39380 9220 39392
rect 9272 39380 9278 39432
rect 11054 39420 11060 39432
rect 11015 39392 11060 39420
rect 11054 39380 11060 39392
rect 11112 39380 11118 39432
rect 11238 39420 11244 39432
rect 11199 39392 11244 39420
rect 11238 39380 11244 39392
rect 11296 39380 11302 39432
rect 14093 39423 14151 39429
rect 14093 39420 14105 39423
rect 12406 39392 14105 39420
rect 4614 39352 4620 39364
rect 4172 39324 4620 39352
rect 4614 39312 4620 39324
rect 4672 39312 4678 39364
rect 5804 39355 5862 39361
rect 5804 39321 5816 39355
rect 5850 39352 5862 39355
rect 6086 39352 6092 39364
rect 5850 39324 6092 39352
rect 5850 39321 5862 39324
rect 5804 39315 5862 39321
rect 6086 39312 6092 39324
rect 6144 39312 6150 39364
rect 9484 39355 9542 39361
rect 9484 39321 9496 39355
rect 9530 39352 9542 39355
rect 9950 39352 9956 39364
rect 9530 39324 9956 39352
rect 9530 39321 9542 39324
rect 9484 39315 9542 39321
rect 9950 39312 9956 39324
rect 10008 39312 10014 39364
rect 12406 39352 12434 39392
rect 14093 39389 14105 39392
rect 14139 39389 14151 39423
rect 14093 39383 14151 39389
rect 14182 39380 14188 39432
rect 14240 39420 14246 39432
rect 14369 39423 14427 39429
rect 14369 39420 14381 39423
rect 14240 39392 14381 39420
rect 14240 39380 14246 39392
rect 14369 39389 14381 39392
rect 14415 39389 14427 39423
rect 22388 39420 22416 39451
rect 14369 39383 14427 39389
rect 22020 39392 22416 39420
rect 22020 39364 22048 39392
rect 22554 39380 22560 39432
rect 22612 39420 22618 39432
rect 23017 39423 23075 39429
rect 23017 39420 23029 39423
rect 22612 39392 23029 39420
rect 22612 39380 22618 39392
rect 23017 39389 23029 39392
rect 23063 39389 23075 39423
rect 23198 39420 23204 39432
rect 23159 39392 23204 39420
rect 23017 39383 23075 39389
rect 23198 39380 23204 39392
rect 23256 39380 23262 39432
rect 23293 39423 23351 39429
rect 23293 39389 23305 39423
rect 23339 39389 23351 39423
rect 23293 39383 23351 39389
rect 23385 39423 23443 39429
rect 23385 39389 23397 39423
rect 23431 39420 23443 39423
rect 23842 39420 23848 39432
rect 23431 39392 23848 39420
rect 23431 39389 23443 39392
rect 23385 39383 23443 39389
rect 10428 39324 12434 39352
rect 13296 39355 13354 39361
rect 6822 39244 6828 39296
rect 6880 39284 6886 39296
rect 6917 39287 6975 39293
rect 6917 39284 6929 39287
rect 6880 39256 6929 39284
rect 6880 39244 6886 39256
rect 6917 39253 6929 39256
rect 6963 39253 6975 39287
rect 6917 39247 6975 39253
rect 8202 39244 8208 39296
rect 8260 39284 8266 39296
rect 10428 39284 10456 39324
rect 13296 39321 13308 39355
rect 13342 39352 13354 39355
rect 13722 39352 13728 39364
rect 13342 39324 13728 39352
rect 13342 39321 13354 39324
rect 13296 39315 13354 39321
rect 13722 39312 13728 39324
rect 13780 39312 13786 39364
rect 22002 39312 22008 39364
rect 22060 39312 22066 39364
rect 22094 39312 22100 39364
rect 22152 39361 22158 39364
rect 22152 39352 22164 39361
rect 22152 39324 22197 39352
rect 22152 39315 22164 39324
rect 22152 39312 22158 39315
rect 22462 39312 22468 39364
rect 22520 39352 22526 39364
rect 22738 39352 22744 39364
rect 22520 39324 22744 39352
rect 22520 39312 22526 39324
rect 22738 39312 22744 39324
rect 22796 39352 22802 39364
rect 23308 39352 23336 39383
rect 23842 39380 23848 39392
rect 23900 39380 23906 39432
rect 24412 39429 24440 39460
rect 24397 39423 24455 39429
rect 24397 39389 24409 39423
rect 24443 39420 24455 39423
rect 27249 39423 27307 39429
rect 24443 39392 24808 39420
rect 24443 39389 24455 39392
rect 24397 39383 24455 39389
rect 24780 39364 24808 39392
rect 27249 39389 27261 39423
rect 27295 39420 27307 39423
rect 27338 39420 27344 39432
rect 27295 39392 27344 39420
rect 27295 39389 27307 39392
rect 27249 39383 27307 39389
rect 27338 39380 27344 39392
rect 27396 39380 27402 39432
rect 28258 39380 28264 39432
rect 28316 39420 28322 39432
rect 30282 39420 30288 39432
rect 28316 39392 30288 39420
rect 28316 39380 28322 39392
rect 30282 39380 30288 39392
rect 30340 39420 30346 39432
rect 30837 39423 30895 39429
rect 31036 39426 31064 39460
rect 30837 39420 30849 39423
rect 30340 39392 30849 39420
rect 30340 39380 30346 39392
rect 30837 39389 30849 39392
rect 30883 39389 30895 39423
rect 30837 39383 30895 39389
rect 31016 39420 31074 39426
rect 31016 39386 31028 39420
rect 31062 39386 31074 39420
rect 31016 39380 31074 39386
rect 31110 39380 31116 39432
rect 31168 39420 31174 39432
rect 31294 39429 31300 39432
rect 31251 39423 31300 39429
rect 31168 39392 31213 39420
rect 31168 39380 31174 39392
rect 31251 39389 31263 39423
rect 31297 39389 31300 39423
rect 31251 39383 31300 39389
rect 31294 39380 31300 39383
rect 31352 39380 31358 39432
rect 22796 39324 23336 39352
rect 23661 39355 23719 39361
rect 22796 39312 22802 39324
rect 23661 39321 23673 39355
rect 23707 39352 23719 39355
rect 24642 39355 24700 39361
rect 24642 39352 24654 39355
rect 23707 39324 24654 39352
rect 23707 39321 23719 39324
rect 23661 39315 23719 39321
rect 24642 39321 24654 39324
rect 24688 39321 24700 39355
rect 24642 39315 24700 39321
rect 24762 39312 24768 39364
rect 24820 39312 24826 39364
rect 27522 39361 27528 39364
rect 27516 39315 27528 39361
rect 27580 39352 27586 39364
rect 27580 39324 27616 39352
rect 27522 39312 27528 39315
rect 27580 39312 27586 39324
rect 31754 39312 31760 39364
rect 31812 39352 31818 39364
rect 31941 39355 31999 39361
rect 31941 39352 31953 39355
rect 31812 39324 31953 39352
rect 31812 39312 31818 39324
rect 31941 39321 31953 39324
rect 31987 39321 31999 39355
rect 31941 39315 31999 39321
rect 32030 39312 32036 39364
rect 32088 39352 32094 39364
rect 32125 39355 32183 39361
rect 32125 39352 32137 39355
rect 32088 39324 32137 39352
rect 32088 39312 32094 39324
rect 32125 39321 32137 39324
rect 32171 39321 32183 39355
rect 32125 39315 32183 39321
rect 10594 39284 10600 39296
rect 8260 39256 10456 39284
rect 10555 39256 10600 39284
rect 8260 39244 8266 39256
rect 10594 39244 10600 39256
rect 10652 39244 10658 39296
rect 16850 39284 16856 39296
rect 16811 39256 16856 39284
rect 16850 39244 16856 39256
rect 16908 39244 16914 39296
rect 20990 39284 20996 39296
rect 20951 39256 20996 39284
rect 20990 39244 20996 39256
rect 21048 39244 21054 39296
rect 23382 39244 23388 39296
rect 23440 39284 23446 39296
rect 25777 39287 25835 39293
rect 25777 39284 25789 39287
rect 23440 39256 25789 39284
rect 23440 39244 23446 39256
rect 25777 39253 25789 39256
rect 25823 39253 25835 39287
rect 28626 39284 28632 39296
rect 28587 39256 28632 39284
rect 25777 39247 25835 39253
rect 28626 39244 28632 39256
rect 28684 39244 28690 39296
rect 30377 39287 30435 39293
rect 30377 39253 30389 39287
rect 30423 39284 30435 39287
rect 30558 39284 30564 39296
rect 30423 39256 30564 39284
rect 30423 39253 30435 39256
rect 30377 39247 30435 39253
rect 30558 39244 30564 39256
rect 30616 39284 30622 39296
rect 31294 39284 31300 39296
rect 30616 39256 31300 39284
rect 30616 39244 30622 39256
rect 31294 39244 31300 39256
rect 31352 39244 31358 39296
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 9950 39080 9956 39092
rect 4356 39052 5120 39080
rect 9911 39052 9956 39080
rect 2676 39015 2734 39021
rect 2676 38981 2688 39015
rect 2722 39012 2734 39015
rect 4249 39015 4307 39021
rect 4249 39012 4261 39015
rect 2722 38984 4261 39012
rect 2722 38981 2734 38984
rect 2676 38975 2734 38981
rect 4249 38981 4261 38984
rect 4295 38981 4307 39015
rect 4249 38975 4307 38981
rect 2409 38947 2467 38953
rect 2409 38913 2421 38947
rect 2455 38944 2467 38947
rect 2498 38944 2504 38956
rect 2455 38916 2504 38944
rect 2455 38913 2467 38916
rect 2409 38907 2467 38913
rect 2498 38904 2504 38916
rect 2556 38904 2562 38956
rect 4356 38944 4384 39052
rect 5092 39024 5120 39052
rect 9950 39040 9956 39052
rect 10008 39040 10014 39092
rect 13078 39080 13084 39092
rect 10060 39052 12434 39080
rect 13039 39052 13084 39080
rect 5074 38972 5080 39024
rect 5132 39012 5138 39024
rect 5445 39015 5503 39021
rect 5445 39012 5457 39015
rect 5132 38984 5457 39012
rect 5132 38972 5138 38984
rect 5445 38981 5457 38984
rect 5491 39012 5503 39015
rect 10060 39012 10088 39052
rect 11517 39015 11575 39021
rect 11517 39012 11529 39015
rect 5491 38984 10088 39012
rect 10244 38984 11529 39012
rect 5491 38981 5503 38984
rect 5445 38975 5503 38981
rect 4479 38947 4537 38953
rect 4479 38944 4491 38947
rect 4356 38916 4491 38944
rect 4479 38913 4491 38916
rect 4525 38913 4537 38947
rect 4614 38944 4620 38956
rect 4575 38916 4620 38944
rect 4479 38907 4537 38913
rect 4614 38904 4620 38916
rect 4672 38904 4678 38956
rect 4730 38947 4788 38953
rect 4730 38913 4742 38947
rect 4776 38944 4788 38947
rect 4776 38916 4844 38944
rect 4776 38913 4788 38916
rect 4730 38907 4788 38913
rect 4816 38876 4844 38916
rect 4890 38904 4896 38956
rect 4948 38944 4954 38956
rect 6362 38944 6368 38956
rect 4948 38916 4993 38944
rect 6323 38916 6368 38944
rect 4948 38904 4954 38916
rect 6362 38904 6368 38916
rect 6420 38904 6426 38956
rect 6549 38947 6607 38953
rect 6549 38913 6561 38947
rect 6595 38944 6607 38947
rect 6822 38944 6828 38956
rect 6595 38916 6828 38944
rect 6595 38913 6607 38916
rect 6549 38907 6607 38913
rect 6822 38904 6828 38916
rect 6880 38904 6886 38956
rect 10244 38953 10272 38984
rect 11517 38981 11529 38984
rect 11563 38981 11575 39015
rect 12406 39012 12434 39052
rect 13078 39040 13084 39052
rect 13136 39040 13142 39092
rect 18322 39080 18328 39092
rect 18283 39052 18328 39080
rect 18322 39040 18328 39052
rect 18380 39040 18386 39092
rect 22646 39040 22652 39092
rect 22704 39080 22710 39092
rect 22833 39083 22891 39089
rect 22833 39080 22845 39083
rect 22704 39052 22845 39080
rect 22704 39040 22710 39052
rect 22833 39049 22845 39052
rect 22879 39049 22891 39083
rect 27522 39080 27528 39092
rect 27483 39052 27528 39080
rect 22833 39043 22891 39049
rect 27522 39040 27528 39052
rect 27580 39040 27586 39092
rect 27982 39040 27988 39092
rect 28040 39040 28046 39092
rect 12406 38984 19334 39012
rect 11517 38975 11575 38981
rect 10209 38947 10272 38953
rect 10209 38913 10221 38947
rect 10255 38916 10272 38947
rect 10334 38950 10392 38956
rect 10334 38916 10346 38950
rect 10380 38916 10392 38950
rect 10434 38947 10492 38953
rect 10434 38944 10446 38947
rect 10255 38913 10267 38916
rect 10209 38907 10267 38913
rect 10334 38910 10392 38916
rect 10428 38913 10446 38944
rect 10480 38913 10492 38947
rect 7837 38879 7895 38885
rect 7837 38876 7849 38879
rect 4724 38848 4844 38876
rect 6564 38848 7849 38876
rect 4724 38820 4752 38848
rect 4706 38768 4712 38820
rect 4764 38768 4770 38820
rect 6564 38752 6592 38848
rect 7837 38845 7849 38848
rect 7883 38845 7895 38879
rect 7837 38839 7895 38845
rect 8113 38879 8171 38885
rect 8113 38845 8125 38879
rect 8159 38876 8171 38879
rect 8202 38876 8208 38888
rect 8159 38848 8208 38876
rect 8159 38845 8171 38848
rect 8113 38839 8171 38845
rect 8202 38836 8208 38848
rect 8260 38836 8266 38888
rect 10336 38876 10364 38910
rect 10152 38848 10364 38876
rect 10428 38907 10492 38913
rect 10597 38947 10655 38953
rect 10597 38913 10609 38947
rect 10643 38944 10655 38947
rect 10686 38944 10692 38956
rect 10643 38916 10692 38944
rect 10643 38913 10655 38916
rect 10597 38907 10655 38913
rect 10152 38820 10180 38848
rect 10428 38820 10456 38907
rect 10686 38904 10692 38916
rect 10744 38904 10750 38956
rect 11532 38876 11560 38975
rect 12894 38944 12900 38956
rect 12855 38916 12900 38944
rect 12894 38904 12900 38916
rect 12952 38904 12958 38956
rect 16850 38904 16856 38956
rect 16908 38944 16914 38956
rect 17037 38947 17095 38953
rect 17037 38944 17049 38947
rect 16908 38916 17049 38944
rect 16908 38904 16914 38916
rect 17037 38913 17049 38916
rect 17083 38913 17095 38947
rect 17037 38907 17095 38913
rect 19306 38876 19334 38984
rect 21450 38972 21456 39024
rect 21508 39012 21514 39024
rect 23106 39012 23112 39024
rect 21508 38984 23112 39012
rect 21508 38972 21514 38984
rect 23106 38972 23112 38984
rect 23164 39012 23170 39024
rect 23201 39015 23259 39021
rect 23201 39012 23213 39015
rect 23164 38984 23213 39012
rect 23164 38972 23170 38984
rect 23201 38981 23213 38984
rect 23247 38981 23259 39015
rect 28000 39012 28028 39040
rect 31110 39012 31116 39024
rect 23201 38975 23259 38981
rect 27908 38984 31116 39012
rect 23017 38947 23075 38953
rect 23017 38913 23029 38947
rect 23063 38944 23075 38947
rect 23566 38944 23572 38956
rect 23063 38916 23572 38944
rect 23063 38913 23075 38916
rect 23017 38907 23075 38913
rect 23566 38904 23572 38916
rect 23624 38904 23630 38956
rect 26970 38944 26976 38956
rect 26883 38916 26976 38944
rect 26970 38904 26976 38916
rect 27028 38944 27034 38956
rect 27908 38953 27936 38984
rect 31110 38972 31116 38984
rect 31168 38972 31174 39024
rect 27781 38947 27839 38953
rect 27781 38944 27793 38947
rect 27028 38916 27793 38944
rect 27028 38904 27034 38916
rect 27781 38913 27793 38916
rect 27827 38913 27839 38947
rect 27781 38907 27839 38913
rect 27893 38947 27951 38953
rect 27893 38913 27905 38947
rect 27939 38913 27951 38947
rect 27893 38907 27951 38913
rect 27985 38947 28043 38953
rect 27985 38913 27997 38947
rect 28031 38944 28043 38947
rect 28169 38947 28227 38953
rect 28031 38916 28120 38944
rect 28031 38913 28043 38916
rect 27985 38907 28043 38913
rect 28092 38888 28120 38916
rect 28169 38913 28181 38947
rect 28215 38944 28227 38947
rect 28258 38944 28264 38956
rect 28215 38916 28264 38944
rect 28215 38913 28227 38916
rect 28169 38907 28227 38913
rect 28258 38904 28264 38916
rect 28316 38904 28322 38956
rect 27062 38876 27068 38888
rect 11532 38848 16574 38876
rect 19306 38848 27068 38876
rect 10134 38768 10140 38820
rect 10192 38768 10198 38820
rect 10410 38768 10416 38820
rect 10468 38768 10474 38820
rect 3789 38743 3847 38749
rect 3789 38709 3801 38743
rect 3835 38740 3847 38743
rect 3970 38740 3976 38752
rect 3835 38712 3976 38740
rect 3835 38709 3847 38712
rect 3789 38703 3847 38709
rect 3970 38700 3976 38712
rect 4028 38700 4034 38752
rect 4614 38700 4620 38752
rect 4672 38740 4678 38752
rect 6546 38740 6552 38752
rect 4672 38712 6552 38740
rect 4672 38700 4678 38712
rect 6546 38700 6552 38712
rect 6604 38700 6610 38752
rect 6638 38700 6644 38752
rect 6696 38740 6702 38752
rect 6733 38743 6791 38749
rect 6733 38740 6745 38743
rect 6696 38712 6745 38740
rect 6696 38700 6702 38712
rect 6733 38709 6745 38712
rect 6779 38709 6791 38743
rect 6733 38703 6791 38709
rect 7282 38700 7288 38752
rect 7340 38740 7346 38752
rect 8573 38743 8631 38749
rect 8573 38740 8585 38743
rect 7340 38712 8585 38740
rect 7340 38700 7346 38712
rect 8573 38709 8585 38712
rect 8619 38740 8631 38743
rect 13814 38740 13820 38752
rect 8619 38712 13820 38740
rect 8619 38709 8631 38712
rect 8573 38703 8631 38709
rect 13814 38700 13820 38712
rect 13872 38700 13878 38752
rect 16546 38740 16574 38848
rect 27062 38836 27068 38848
rect 27120 38836 27126 38888
rect 28074 38836 28080 38888
rect 28132 38836 28138 38888
rect 58158 38808 58164 38820
rect 58119 38780 58164 38808
rect 58158 38768 58164 38780
rect 58216 38768 58222 38820
rect 18966 38740 18972 38752
rect 16546 38712 18972 38740
rect 18966 38700 18972 38712
rect 19024 38740 19030 38752
rect 23842 38740 23848 38752
rect 19024 38712 23848 38740
rect 19024 38700 19030 38712
rect 23842 38700 23848 38712
rect 23900 38740 23906 38752
rect 26786 38740 26792 38752
rect 23900 38712 26792 38740
rect 23900 38700 23906 38712
rect 26786 38700 26792 38712
rect 26844 38700 26850 38752
rect 28810 38700 28816 38752
rect 28868 38740 28874 38752
rect 29641 38743 29699 38749
rect 29641 38740 29653 38743
rect 28868 38712 29653 38740
rect 28868 38700 28874 38712
rect 29641 38709 29653 38712
rect 29687 38709 29699 38743
rect 29641 38703 29699 38709
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 4157 38539 4215 38545
rect 4157 38505 4169 38539
rect 4203 38536 4215 38539
rect 4706 38536 4712 38548
rect 4203 38508 4712 38536
rect 4203 38505 4215 38508
rect 4157 38499 4215 38505
rect 4706 38496 4712 38508
rect 4764 38496 4770 38548
rect 6086 38536 6092 38548
rect 6047 38508 6092 38536
rect 6086 38496 6092 38508
rect 6144 38496 6150 38548
rect 17494 38536 17500 38548
rect 16040 38508 17500 38536
rect 6454 38468 6460 38480
rect 6196 38440 6460 38468
rect 4614 38400 4620 38412
rect 2976 38372 4620 38400
rect 2866 38332 2872 38344
rect 2827 38304 2872 38332
rect 2866 38292 2872 38304
rect 2924 38292 2930 38344
rect 2976 38341 3004 38372
rect 4614 38360 4620 38372
rect 4672 38360 4678 38412
rect 2961 38335 3019 38341
rect 2961 38301 2973 38335
rect 3007 38301 3019 38335
rect 2961 38295 3019 38301
rect 3050 38292 3056 38344
rect 3108 38332 3114 38344
rect 3237 38335 3295 38341
rect 3108 38304 3153 38332
rect 3108 38292 3114 38304
rect 3237 38301 3249 38335
rect 3283 38332 3295 38335
rect 4890 38332 4896 38344
rect 3283 38304 4896 38332
rect 3283 38301 3295 38304
rect 3237 38295 3295 38301
rect 4890 38292 4896 38304
rect 4948 38292 4954 38344
rect 6196 38326 6224 38440
rect 6454 38428 6460 38440
rect 6512 38428 6518 38480
rect 6638 38360 6644 38412
rect 6696 38360 6702 38412
rect 6345 38335 6403 38341
rect 6345 38326 6357 38335
rect 6196 38301 6357 38326
rect 6391 38301 6403 38335
rect 6196 38298 6403 38301
rect 6345 38295 6403 38298
rect 6454 38335 6512 38341
rect 6454 38301 6466 38335
rect 6500 38332 6512 38335
rect 6549 38335 6607 38341
rect 6500 38301 6513 38332
rect 6454 38295 6513 38301
rect 6549 38301 6561 38335
rect 6595 38332 6607 38335
rect 6656 38332 6684 38360
rect 6595 38304 6684 38332
rect 6595 38301 6607 38304
rect 6549 38295 6607 38301
rect 3789 38267 3847 38273
rect 3789 38233 3801 38267
rect 3835 38233 3847 38267
rect 3970 38264 3976 38276
rect 3931 38236 3976 38264
rect 3789 38227 3847 38233
rect 2130 38156 2136 38208
rect 2188 38196 2194 38208
rect 2593 38199 2651 38205
rect 2593 38196 2605 38199
rect 2188 38168 2605 38196
rect 2188 38156 2194 38168
rect 2593 38165 2605 38168
rect 2639 38165 2651 38199
rect 2593 38159 2651 38165
rect 3418 38156 3424 38208
rect 3476 38196 3482 38208
rect 3804 38196 3832 38227
rect 3970 38224 3976 38236
rect 4028 38224 4034 38276
rect 6485 38264 6513 38295
rect 6730 38292 6736 38344
rect 6788 38332 6794 38344
rect 7650 38332 7656 38344
rect 6788 38304 7656 38332
rect 6788 38292 6794 38304
rect 7650 38292 7656 38304
rect 7708 38292 7714 38344
rect 10594 38292 10600 38344
rect 10652 38332 10658 38344
rect 16040 38341 16068 38508
rect 17494 38496 17500 38508
rect 17552 38496 17558 38548
rect 23474 38496 23480 38548
rect 23532 38536 23538 38548
rect 25498 38536 25504 38548
rect 23532 38508 25504 38536
rect 23532 38496 23538 38508
rect 25498 38496 25504 38508
rect 25556 38496 25562 38548
rect 28074 38536 28080 38548
rect 28035 38508 28080 38536
rect 28074 38496 28080 38508
rect 28132 38496 28138 38548
rect 16301 38471 16359 38477
rect 16301 38437 16313 38471
rect 16347 38437 16359 38471
rect 16301 38431 16359 38437
rect 16316 38400 16344 38431
rect 30929 38403 30987 38409
rect 16316 38372 19380 38400
rect 15749 38335 15807 38341
rect 15749 38332 15761 38335
rect 10652 38304 15761 38332
rect 10652 38292 10658 38304
rect 15749 38301 15761 38304
rect 15795 38301 15807 38335
rect 15749 38295 15807 38301
rect 16025 38335 16083 38341
rect 16025 38301 16037 38335
rect 16071 38301 16083 38335
rect 16025 38295 16083 38301
rect 16114 38292 16120 38344
rect 16172 38332 16178 38344
rect 16758 38332 16764 38344
rect 16172 38304 16217 38332
rect 16719 38304 16764 38332
rect 16172 38292 16178 38304
rect 16758 38292 16764 38304
rect 16816 38292 16822 38344
rect 17034 38332 17040 38344
rect 16995 38304 17040 38332
rect 17034 38292 17040 38304
rect 17092 38292 17098 38344
rect 17126 38292 17132 38344
rect 17184 38332 17190 38344
rect 19352 38341 19380 38372
rect 30929 38369 30941 38403
rect 30975 38400 30987 38403
rect 31202 38400 31208 38412
rect 30975 38372 31208 38400
rect 30975 38369 30987 38372
rect 30929 38363 30987 38369
rect 31202 38360 31208 38372
rect 31260 38400 31266 38412
rect 31662 38400 31668 38412
rect 31260 38372 31668 38400
rect 31260 38360 31266 38372
rect 31662 38360 31668 38372
rect 31720 38360 31726 38412
rect 19337 38335 19395 38341
rect 17184 38304 17229 38332
rect 17184 38292 17190 38304
rect 19337 38301 19349 38335
rect 19383 38301 19395 38335
rect 19337 38295 19395 38301
rect 19426 38292 19432 38344
rect 19484 38332 19490 38344
rect 19843 38335 19901 38341
rect 19484 38304 19529 38332
rect 19484 38292 19490 38304
rect 19843 38301 19855 38335
rect 19889 38332 19901 38335
rect 20254 38332 20260 38344
rect 19889 38304 20260 38332
rect 19889 38301 19901 38304
rect 19843 38295 19901 38301
rect 20254 38292 20260 38304
rect 20312 38292 20318 38344
rect 24581 38335 24639 38341
rect 24581 38301 24593 38335
rect 24627 38332 24639 38335
rect 24670 38332 24676 38344
rect 24627 38304 24676 38332
rect 24627 38301 24639 38304
rect 24581 38295 24639 38301
rect 24670 38292 24676 38304
rect 24728 38292 24734 38344
rect 28261 38335 28319 38341
rect 28261 38301 28273 38335
rect 28307 38332 28319 38335
rect 28626 38332 28632 38344
rect 28307 38304 28632 38332
rect 28307 38301 28319 38304
rect 28261 38295 28319 38301
rect 28626 38292 28632 38304
rect 28684 38292 28690 38344
rect 30190 38292 30196 38344
rect 30248 38332 30254 38344
rect 31573 38335 31631 38341
rect 30248 38304 30788 38332
rect 30248 38292 30254 38304
rect 6638 38264 6644 38276
rect 6485 38236 6644 38264
rect 6638 38224 6644 38236
rect 6696 38224 6702 38276
rect 9306 38264 9312 38276
rect 9267 38236 9312 38264
rect 9306 38224 9312 38236
rect 9364 38224 9370 38276
rect 15930 38264 15936 38276
rect 15843 38236 15936 38264
rect 15930 38224 15936 38236
rect 15988 38264 15994 38276
rect 16945 38267 17003 38273
rect 15988 38236 16252 38264
rect 15988 38224 15994 38236
rect 6362 38196 6368 38208
rect 3476 38168 6368 38196
rect 3476 38156 3482 38168
rect 6362 38156 6368 38168
rect 6420 38156 6426 38208
rect 6454 38156 6460 38208
rect 6512 38196 6518 38208
rect 7285 38199 7343 38205
rect 7285 38196 7297 38199
rect 6512 38168 7297 38196
rect 6512 38156 6518 38168
rect 7285 38165 7297 38168
rect 7331 38196 7343 38199
rect 8018 38196 8024 38208
rect 7331 38168 8024 38196
rect 7331 38165 7343 38168
rect 7285 38159 7343 38165
rect 8018 38156 8024 38168
rect 8076 38156 8082 38208
rect 9214 38156 9220 38208
rect 9272 38196 9278 38208
rect 10226 38196 10232 38208
rect 9272 38168 10232 38196
rect 9272 38156 9278 38168
rect 10226 38156 10232 38168
rect 10284 38196 10290 38208
rect 10597 38199 10655 38205
rect 10597 38196 10609 38199
rect 10284 38168 10609 38196
rect 10284 38156 10290 38168
rect 10597 38165 10609 38168
rect 10643 38165 10655 38199
rect 16224 38196 16252 38236
rect 16945 38233 16957 38267
rect 16991 38233 17003 38267
rect 16945 38227 17003 38233
rect 16960 38196 16988 38227
rect 19242 38224 19248 38276
rect 19300 38264 19306 38276
rect 19613 38267 19671 38273
rect 19613 38264 19625 38267
rect 19300 38236 19625 38264
rect 19300 38224 19306 38236
rect 19613 38233 19625 38236
rect 19659 38233 19671 38267
rect 19613 38227 19671 38233
rect 19705 38267 19763 38273
rect 19705 38233 19717 38267
rect 19751 38264 19763 38267
rect 20622 38264 20628 38276
rect 19751 38236 20628 38264
rect 19751 38233 19763 38236
rect 19705 38227 19763 38233
rect 20622 38224 20628 38236
rect 20680 38224 20686 38276
rect 24394 38224 24400 38276
rect 24452 38264 24458 38276
rect 24826 38267 24884 38273
rect 24826 38264 24838 38267
rect 24452 38236 24838 38264
rect 24452 38224 24458 38236
rect 24826 38233 24838 38236
rect 24872 38233 24884 38267
rect 24826 38227 24884 38233
rect 28445 38267 28503 38273
rect 28445 38233 28457 38267
rect 28491 38264 28503 38267
rect 29086 38264 29092 38276
rect 28491 38236 29092 38264
rect 28491 38233 28503 38236
rect 28445 38227 28503 38233
rect 29086 38224 29092 38236
rect 29144 38264 29150 38276
rect 30208 38264 30236 38292
rect 29144 38236 30236 38264
rect 29144 38224 29150 38236
rect 30374 38224 30380 38276
rect 30432 38264 30438 38276
rect 30662 38267 30720 38273
rect 30662 38264 30674 38267
rect 30432 38236 30674 38264
rect 30432 38224 30438 38236
rect 30662 38233 30674 38236
rect 30708 38233 30720 38267
rect 30760 38264 30788 38304
rect 31573 38301 31585 38335
rect 31619 38332 31631 38335
rect 31938 38332 31944 38344
rect 31619 38304 31944 38332
rect 31619 38301 31631 38304
rect 31573 38295 31631 38301
rect 31938 38292 31944 38304
rect 31996 38292 32002 38344
rect 31754 38264 31760 38276
rect 30760 38236 31760 38264
rect 30662 38227 30720 38233
rect 31754 38224 31760 38236
rect 31812 38264 31818 38276
rect 31812 38236 31857 38264
rect 31812 38224 31818 38236
rect 17310 38196 17316 38208
rect 16224 38168 16988 38196
rect 17271 38168 17316 38196
rect 10597 38159 10655 38165
rect 17310 38156 17316 38168
rect 17368 38156 17374 38208
rect 19981 38199 20039 38205
rect 19981 38165 19993 38199
rect 20027 38196 20039 38199
rect 21082 38196 21088 38208
rect 20027 38168 21088 38196
rect 20027 38165 20039 38168
rect 19981 38159 20039 38165
rect 21082 38156 21088 38168
rect 21140 38156 21146 38208
rect 25958 38196 25964 38208
rect 25919 38168 25964 38196
rect 25958 38156 25964 38168
rect 26016 38156 26022 38208
rect 29546 38196 29552 38208
rect 29507 38168 29552 38196
rect 29546 38156 29552 38168
rect 29604 38156 29610 38208
rect 30466 38156 30472 38208
rect 30524 38196 30530 38208
rect 31389 38199 31447 38205
rect 31389 38196 31401 38199
rect 30524 38168 31401 38196
rect 30524 38156 30530 38168
rect 31389 38165 31401 38168
rect 31435 38165 31447 38199
rect 32306 38196 32312 38208
rect 32267 38168 32312 38196
rect 31389 38159 31447 38165
rect 32306 38156 32312 38168
rect 32364 38156 32370 38208
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 3050 37992 3056 38004
rect 3011 37964 3056 37992
rect 3050 37952 3056 37964
rect 3108 37952 3114 38004
rect 6362 37952 6368 38004
rect 6420 37992 6426 38004
rect 8297 37995 8355 38001
rect 8297 37992 8309 37995
rect 6420 37964 8309 37992
rect 6420 37952 6426 37964
rect 8297 37961 8309 37964
rect 8343 37961 8355 37995
rect 8297 37955 8355 37961
rect 10042 37952 10048 38004
rect 10100 37992 10106 38004
rect 10229 37995 10287 38001
rect 10229 37992 10241 37995
rect 10100 37964 10241 37992
rect 10100 37952 10106 37964
rect 10229 37961 10241 37964
rect 10275 37961 10287 37995
rect 12526 37992 12532 38004
rect 10229 37955 10287 37961
rect 11716 37964 12532 37992
rect 3418 37924 3424 37936
rect 3379 37896 3424 37924
rect 3418 37884 3424 37896
rect 3476 37884 3482 37936
rect 10410 37924 10416 37936
rect 10371 37896 10416 37924
rect 10410 37884 10416 37896
rect 10468 37884 10474 37936
rect 10597 37927 10655 37933
rect 10597 37893 10609 37927
rect 10643 37924 10655 37927
rect 11054 37924 11060 37936
rect 10643 37896 11060 37924
rect 10643 37893 10655 37896
rect 10597 37887 10655 37893
rect 11054 37884 11060 37896
rect 11112 37884 11118 37936
rect 11716 37933 11744 37964
rect 12526 37952 12532 37964
rect 12584 37992 12590 38004
rect 15930 37992 15936 38004
rect 12584 37964 15936 37992
rect 12584 37952 12590 37964
rect 15930 37952 15936 37964
rect 15988 37952 15994 38004
rect 19242 37992 19248 38004
rect 17604 37964 19248 37992
rect 11701 37927 11759 37933
rect 11701 37893 11713 37927
rect 11747 37893 11759 37927
rect 11701 37887 11759 37893
rect 11793 37927 11851 37933
rect 11793 37893 11805 37927
rect 11839 37924 11851 37927
rect 12434 37924 12440 37936
rect 11839 37896 12440 37924
rect 11839 37893 11851 37896
rect 11793 37887 11851 37893
rect 12434 37884 12440 37896
rect 12492 37884 12498 37936
rect 17604 37933 17632 37964
rect 19242 37952 19248 37964
rect 19300 37992 19306 38004
rect 19610 37992 19616 38004
rect 19300 37964 19616 37992
rect 19300 37952 19306 37964
rect 19610 37952 19616 37964
rect 19668 37952 19674 38004
rect 24394 37992 24400 38004
rect 24355 37964 24400 37992
rect 24394 37952 24400 37964
rect 24452 37952 24458 38004
rect 25869 37995 25927 38001
rect 25869 37992 25881 37995
rect 24504 37964 25544 37992
rect 17589 37927 17647 37933
rect 17589 37893 17601 37927
rect 17635 37893 17647 37927
rect 17589 37887 17647 37893
rect 17681 37927 17739 37933
rect 17681 37893 17693 37927
rect 17727 37924 17739 37927
rect 19978 37924 19984 37936
rect 17727 37896 19984 37924
rect 17727 37893 17739 37896
rect 17681 37887 17739 37893
rect 19978 37884 19984 37896
rect 20036 37884 20042 37936
rect 23474 37884 23480 37936
rect 23532 37924 23538 37936
rect 24504 37924 24532 37964
rect 23532 37896 24532 37924
rect 23532 37884 23538 37896
rect 3234 37856 3240 37868
rect 3195 37828 3240 37856
rect 3234 37816 3240 37828
rect 3292 37816 3298 37868
rect 8481 37859 8539 37865
rect 8481 37825 8493 37859
rect 8527 37856 8539 37859
rect 8527 37828 10364 37856
rect 8527 37825 8539 37828
rect 8481 37819 8539 37825
rect 10336 37788 10364 37828
rect 11238 37816 11244 37868
rect 11296 37856 11302 37868
rect 11517 37859 11575 37865
rect 11517 37856 11529 37859
rect 11296 37828 11529 37856
rect 11296 37816 11302 37828
rect 11517 37825 11529 37828
rect 11563 37825 11575 37859
rect 11882 37856 11888 37868
rect 11843 37828 11888 37856
rect 11517 37819 11575 37825
rect 11882 37816 11888 37828
rect 11940 37856 11946 37868
rect 16114 37856 16120 37868
rect 11940 37828 16120 37856
rect 11940 37816 11946 37828
rect 16114 37816 16120 37828
rect 16172 37856 16178 37868
rect 17126 37856 17132 37868
rect 16172 37828 17132 37856
rect 16172 37816 16178 37828
rect 17126 37816 17132 37828
rect 17184 37816 17190 37868
rect 17310 37856 17316 37868
rect 17271 37828 17316 37856
rect 17310 37816 17316 37828
rect 17368 37816 17374 37868
rect 17402 37816 17408 37868
rect 17460 37856 17466 37868
rect 17819 37859 17877 37865
rect 17460 37828 17505 37856
rect 17460 37816 17466 37828
rect 17819 37825 17831 37859
rect 17865 37856 17877 37859
rect 17865 37828 18184 37856
rect 17865 37825 17877 37828
rect 17819 37819 17877 37825
rect 12894 37788 12900 37800
rect 10336 37760 12900 37788
rect 12894 37748 12900 37760
rect 12952 37748 12958 37800
rect 12069 37723 12127 37729
rect 12069 37689 12081 37723
rect 12115 37720 12127 37723
rect 17862 37720 17868 37732
rect 12115 37692 17868 37720
rect 12115 37689 12127 37692
rect 12069 37683 12127 37689
rect 17862 37680 17868 37692
rect 17920 37680 17926 37732
rect 2866 37612 2872 37664
rect 2924 37652 2930 37664
rect 3973 37655 4031 37661
rect 3973 37652 3985 37655
rect 2924 37624 3985 37652
rect 2924 37612 2930 37624
rect 3973 37621 3985 37624
rect 4019 37652 4031 37655
rect 5626 37652 5632 37664
rect 4019 37624 5632 37652
rect 4019 37621 4031 37624
rect 3973 37615 4031 37621
rect 5626 37612 5632 37624
rect 5684 37612 5690 37664
rect 8294 37612 8300 37664
rect 8352 37652 8358 37664
rect 9125 37655 9183 37661
rect 9125 37652 9137 37655
rect 8352 37624 9137 37652
rect 8352 37612 8358 37624
rect 9125 37621 9137 37624
rect 9171 37652 9183 37655
rect 9306 37652 9312 37664
rect 9171 37624 9312 37652
rect 9171 37621 9183 37624
rect 9125 37615 9183 37621
rect 9306 37612 9312 37624
rect 9364 37612 9370 37664
rect 17954 37652 17960 37664
rect 17915 37624 17960 37652
rect 17954 37612 17960 37624
rect 18012 37612 18018 37664
rect 18156 37652 18184 37828
rect 18322 37816 18328 37868
rect 18380 37856 18386 37868
rect 18417 37859 18475 37865
rect 18417 37856 18429 37859
rect 18380 37828 18429 37856
rect 18380 37816 18386 37828
rect 18417 37825 18429 37828
rect 18463 37825 18475 37859
rect 18417 37819 18475 37825
rect 18506 37816 18512 37868
rect 18564 37856 18570 37868
rect 18673 37859 18731 37865
rect 18673 37856 18685 37859
rect 18564 37828 18685 37856
rect 18564 37816 18570 37828
rect 18673 37825 18685 37828
rect 18719 37825 18731 37859
rect 18673 37819 18731 37825
rect 20070 37816 20076 37868
rect 20128 37856 20134 37868
rect 20257 37859 20315 37865
rect 20257 37856 20269 37859
rect 20128 37828 20269 37856
rect 20128 37816 20134 37828
rect 20257 37825 20269 37828
rect 20303 37825 20315 37859
rect 20438 37856 20444 37868
rect 20399 37828 20444 37856
rect 20257 37819 20315 37825
rect 20438 37816 20444 37828
rect 20496 37816 20502 37868
rect 24118 37816 24124 37868
rect 24176 37856 24182 37868
rect 24673 37859 24731 37865
rect 24673 37856 24685 37859
rect 24176 37828 24685 37856
rect 24176 37816 24182 37828
rect 24673 37825 24685 37828
rect 24719 37825 24731 37859
rect 24673 37819 24731 37825
rect 24765 37859 24823 37865
rect 24765 37825 24777 37859
rect 24811 37825 24823 37859
rect 24765 37819 24823 37825
rect 24857 37859 24915 37865
rect 24857 37825 24869 37859
rect 24903 37825 24915 37859
rect 24857 37819 24915 37825
rect 20254 37720 20260 37732
rect 19352 37692 20260 37720
rect 19352 37652 19380 37692
rect 20254 37680 20260 37692
rect 20312 37680 20318 37732
rect 24670 37680 24676 37732
rect 24728 37720 24734 37732
rect 24780 37720 24808 37819
rect 24872 37788 24900 37819
rect 24946 37816 24952 37868
rect 25004 37856 25010 37868
rect 25516 37865 25544 37964
rect 25608 37964 25881 37992
rect 25041 37859 25099 37865
rect 25041 37856 25053 37859
rect 25004 37828 25053 37856
rect 25004 37816 25010 37828
rect 25041 37825 25053 37828
rect 25087 37825 25099 37859
rect 25041 37819 25099 37825
rect 25501 37859 25559 37865
rect 25501 37825 25513 37859
rect 25547 37825 25559 37859
rect 25501 37819 25559 37825
rect 25608 37788 25636 37964
rect 25869 37961 25881 37964
rect 25915 37961 25927 37995
rect 25869 37955 25927 37961
rect 25685 37927 25743 37933
rect 25685 37893 25697 37927
rect 25731 37924 25743 37927
rect 25958 37924 25964 37936
rect 25731 37896 25964 37924
rect 25731 37893 25743 37896
rect 25685 37887 25743 37893
rect 24872 37760 25636 37788
rect 24728 37692 24808 37720
rect 24728 37680 24734 37692
rect 18156 37624 19380 37652
rect 19426 37612 19432 37664
rect 19484 37652 19490 37664
rect 19797 37655 19855 37661
rect 19797 37652 19809 37655
rect 19484 37624 19809 37652
rect 19484 37612 19490 37624
rect 19797 37621 19809 37624
rect 19843 37621 19855 37655
rect 19797 37615 19855 37621
rect 19978 37612 19984 37664
rect 20036 37652 20042 37664
rect 20625 37655 20683 37661
rect 20625 37652 20637 37655
rect 20036 37624 20637 37652
rect 20036 37612 20042 37624
rect 20625 37621 20637 37624
rect 20671 37621 20683 37655
rect 20625 37615 20683 37621
rect 23014 37612 23020 37664
rect 23072 37652 23078 37664
rect 23293 37655 23351 37661
rect 23293 37652 23305 37655
rect 23072 37624 23305 37652
rect 23072 37612 23078 37624
rect 23293 37621 23305 37624
rect 23339 37621 23351 37655
rect 23293 37615 23351 37621
rect 23937 37655 23995 37661
rect 23937 37621 23949 37655
rect 23983 37652 23995 37655
rect 24118 37652 24124 37664
rect 23983 37624 24124 37652
rect 23983 37621 23995 37624
rect 23937 37615 23995 37621
rect 24118 37612 24124 37624
rect 24176 37612 24182 37664
rect 24578 37612 24584 37664
rect 24636 37652 24642 37664
rect 25700 37652 25728 37887
rect 25958 37884 25964 37896
rect 26016 37884 26022 37936
rect 27801 37859 27859 37865
rect 27801 37825 27813 37859
rect 27847 37856 27859 37859
rect 28810 37856 28816 37868
rect 27847 37828 28816 37856
rect 27847 37825 27859 37828
rect 27801 37819 27859 37825
rect 28810 37816 28816 37828
rect 28868 37816 28874 37868
rect 30282 37856 30288 37868
rect 30243 37828 30288 37856
rect 30282 37816 30288 37828
rect 30340 37816 30346 37868
rect 30466 37856 30472 37868
rect 30427 37828 30472 37856
rect 30466 37816 30472 37828
rect 30524 37816 30530 37868
rect 30561 37859 30619 37865
rect 30561 37825 30573 37859
rect 30607 37825 30619 37859
rect 30561 37819 30619 37825
rect 30576 37788 30604 37819
rect 30650 37816 30656 37868
rect 30708 37856 30714 37868
rect 32582 37865 32588 37868
rect 31389 37859 31447 37865
rect 31389 37856 31401 37859
rect 30708 37828 31401 37856
rect 30708 37816 30714 37828
rect 31389 37825 31401 37828
rect 31435 37825 31447 37859
rect 31389 37819 31447 37825
rect 32576 37819 32588 37865
rect 32640 37856 32646 37868
rect 32640 37828 32676 37856
rect 32582 37816 32588 37819
rect 32640 37816 32646 37828
rect 31110 37788 31116 37800
rect 30576 37760 31116 37788
rect 31110 37748 31116 37760
rect 31168 37748 31174 37800
rect 31662 37748 31668 37800
rect 31720 37788 31726 37800
rect 32309 37791 32367 37797
rect 32309 37788 32321 37791
rect 31720 37760 32321 37788
rect 31720 37748 31726 37760
rect 32309 37757 32321 37760
rect 32355 37757 32367 37791
rect 32309 37751 32367 37757
rect 24636 37624 25728 37652
rect 24636 37612 24642 37624
rect 27430 37612 27436 37664
rect 27488 37652 27494 37664
rect 28902 37652 28908 37664
rect 27488 37624 28908 37652
rect 27488 37612 27494 37624
rect 28902 37612 28908 37624
rect 28960 37652 28966 37664
rect 29089 37655 29147 37661
rect 29089 37652 29101 37655
rect 28960 37624 29101 37652
rect 28960 37612 28966 37624
rect 29089 37621 29101 37624
rect 29135 37621 29147 37655
rect 30926 37652 30932 37664
rect 30887 37624 30932 37652
rect 29089 37615 29147 37621
rect 30926 37612 30932 37624
rect 30984 37612 30990 37664
rect 33689 37655 33747 37661
rect 33689 37621 33701 37655
rect 33735 37652 33747 37655
rect 33778 37652 33784 37664
rect 33735 37624 33784 37652
rect 33735 37621 33747 37624
rect 33689 37615 33747 37621
rect 33778 37612 33784 37624
rect 33836 37612 33842 37664
rect 34609 37655 34667 37661
rect 34609 37621 34621 37655
rect 34655 37652 34667 37655
rect 35526 37652 35532 37664
rect 34655 37624 35532 37652
rect 34655 37621 34667 37624
rect 34609 37615 34667 37621
rect 35526 37612 35532 37624
rect 35584 37612 35590 37664
rect 58158 37652 58164 37664
rect 58119 37624 58164 37652
rect 58158 37612 58164 37624
rect 58216 37612 58222 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 16758 37448 16764 37460
rect 16671 37420 16764 37448
rect 16758 37408 16764 37420
rect 16816 37448 16822 37460
rect 17402 37448 17408 37460
rect 16816 37420 17408 37448
rect 16816 37408 16822 37420
rect 17402 37408 17408 37420
rect 17460 37408 17466 37460
rect 18233 37451 18291 37457
rect 18233 37417 18245 37451
rect 18279 37448 18291 37451
rect 18506 37448 18512 37460
rect 18279 37420 18512 37448
rect 18279 37417 18291 37420
rect 18233 37411 18291 37417
rect 18506 37408 18512 37420
rect 18564 37408 18570 37460
rect 20438 37448 20444 37460
rect 20399 37420 20444 37448
rect 20438 37408 20444 37420
rect 20496 37408 20502 37460
rect 7009 37383 7067 37389
rect 7009 37349 7021 37383
rect 7055 37349 7067 37383
rect 7009 37343 7067 37349
rect 7024 37312 7052 37343
rect 17862 37340 17868 37392
rect 17920 37380 17926 37392
rect 17920 37352 19380 37380
rect 17920 37340 17926 37352
rect 18966 37312 18972 37324
rect 7024 37284 7512 37312
rect 7484 37256 7512 37284
rect 15212 37284 15516 37312
rect 1857 37247 1915 37253
rect 1857 37213 1869 37247
rect 1903 37244 1915 37247
rect 2590 37244 2596 37256
rect 1903 37216 2596 37244
rect 1903 37213 1915 37216
rect 1857 37207 1915 37213
rect 2590 37204 2596 37216
rect 2648 37204 2654 37256
rect 5629 37247 5687 37253
rect 5629 37213 5641 37247
rect 5675 37244 5687 37247
rect 5675 37216 7420 37244
rect 5675 37213 5687 37216
rect 5629 37207 5687 37213
rect 2130 37185 2136 37188
rect 2124 37176 2136 37185
rect 2091 37148 2136 37176
rect 2124 37139 2136 37148
rect 2130 37136 2136 37139
rect 2188 37136 2194 37188
rect 5896 37179 5954 37185
rect 5896 37145 5908 37179
rect 5942 37176 5954 37179
rect 7006 37176 7012 37188
rect 5942 37148 7012 37176
rect 5942 37145 5954 37148
rect 5896 37139 5954 37145
rect 7006 37136 7012 37148
rect 7064 37136 7070 37188
rect 3234 37108 3240 37120
rect 3195 37080 3240 37108
rect 3234 37068 3240 37080
rect 3292 37068 3298 37120
rect 7392 37108 7420 37216
rect 7466 37204 7472 37256
rect 7524 37244 7530 37256
rect 7742 37244 7748 37256
rect 7524 37216 7617 37244
rect 7703 37216 7748 37244
rect 7524 37204 7530 37216
rect 7742 37204 7748 37216
rect 7800 37204 7806 37256
rect 7834 37204 7840 37256
rect 7892 37244 7898 37256
rect 11882 37244 11888 37256
rect 7892 37216 11888 37244
rect 7892 37204 7898 37216
rect 11882 37204 11888 37216
rect 11940 37244 11946 37256
rect 13170 37244 13176 37256
rect 11940 37216 13176 37244
rect 11940 37204 11946 37216
rect 13170 37204 13176 37216
rect 13228 37204 13234 37256
rect 14093 37247 14151 37253
rect 14093 37213 14105 37247
rect 14139 37244 14151 37247
rect 15212 37244 15240 37284
rect 15378 37244 15384 37256
rect 14139 37216 15240 37244
rect 15339 37216 15384 37244
rect 14139 37213 14151 37216
rect 14093 37207 14151 37213
rect 15378 37204 15384 37216
rect 15436 37204 15442 37256
rect 15488 37244 15516 37284
rect 17972 37284 18972 37312
rect 17034 37244 17040 37256
rect 15488 37216 17040 37244
rect 17034 37204 17040 37216
rect 17092 37204 17098 37256
rect 17586 37204 17592 37256
rect 17644 37253 17650 37256
rect 17644 37244 17653 37253
rect 17770 37244 17776 37256
rect 17644 37216 17689 37244
rect 17731 37216 17776 37244
rect 17644 37207 17653 37216
rect 17644 37204 17650 37207
rect 17770 37204 17776 37216
rect 17828 37204 17834 37256
rect 17972 37253 18000 37284
rect 18966 37272 18972 37284
rect 19024 37272 19030 37324
rect 19352 37253 19380 37352
rect 20456 37312 20484 37408
rect 23014 37340 23020 37392
rect 23072 37380 23078 37392
rect 24397 37383 24455 37389
rect 24397 37380 24409 37383
rect 23072 37352 24409 37380
rect 23072 37340 23078 37352
rect 24397 37349 24409 37352
rect 24443 37349 24455 37383
rect 24397 37343 24455 37349
rect 31662 37340 31668 37392
rect 31720 37380 31726 37392
rect 33689 37383 33747 37389
rect 33689 37380 33701 37383
rect 31720 37352 33701 37380
rect 31720 37340 31726 37352
rect 33689 37349 33701 37352
rect 33735 37380 33747 37383
rect 34882 37380 34888 37392
rect 33735 37352 34888 37380
rect 33735 37349 33747 37352
rect 33689 37343 33747 37349
rect 34882 37340 34888 37352
rect 34940 37340 34946 37392
rect 19720 37284 20484 37312
rect 19720 37253 19748 37284
rect 17865 37247 17923 37253
rect 17865 37213 17877 37247
rect 17911 37213 17923 37247
rect 17972 37247 18035 37253
rect 17972 37216 17989 37247
rect 17865 37207 17923 37213
rect 17977 37213 17989 37216
rect 18023 37213 18035 37247
rect 17977 37207 18035 37213
rect 19337 37247 19395 37253
rect 19337 37213 19349 37247
rect 19383 37213 19395 37247
rect 19337 37207 19395 37213
rect 19430 37247 19488 37253
rect 19430 37213 19442 37247
rect 19476 37213 19488 37247
rect 19430 37207 19488 37213
rect 19705 37247 19763 37253
rect 19705 37213 19717 37247
rect 19751 37213 19763 37247
rect 19705 37207 19763 37213
rect 19843 37247 19901 37253
rect 19843 37213 19855 37247
rect 19889 37244 19901 37247
rect 20254 37244 20260 37256
rect 19889 37216 20260 37244
rect 19889 37213 19901 37216
rect 19843 37207 19901 37213
rect 7650 37176 7656 37188
rect 7611 37148 7656 37176
rect 7650 37136 7656 37148
rect 7708 37136 7714 37188
rect 10226 37176 10232 37188
rect 7760 37148 10232 37176
rect 7760 37108 7788 37148
rect 10226 37136 10232 37148
rect 10284 37136 10290 37188
rect 14277 37179 14335 37185
rect 14277 37145 14289 37179
rect 14323 37176 14335 37179
rect 14642 37176 14648 37188
rect 14323 37148 14648 37176
rect 14323 37145 14335 37148
rect 14277 37139 14335 37145
rect 14642 37136 14648 37148
rect 14700 37176 14706 37188
rect 14700 37148 15424 37176
rect 14700 37136 14706 37148
rect 7392 37080 7788 37108
rect 8021 37111 8079 37117
rect 8021 37077 8033 37111
rect 8067 37108 8079 37111
rect 8386 37108 8392 37120
rect 8067 37080 8392 37108
rect 8067 37077 8079 37080
rect 8021 37071 8079 37077
rect 8386 37068 8392 37080
rect 8444 37068 8450 37120
rect 14461 37111 14519 37117
rect 14461 37077 14473 37111
rect 14507 37108 14519 37111
rect 14550 37108 14556 37120
rect 14507 37080 14556 37108
rect 14507 37077 14519 37080
rect 14461 37071 14519 37077
rect 14550 37068 14556 37080
rect 14608 37068 14614 37120
rect 15396 37108 15424 37148
rect 15470 37136 15476 37188
rect 15528 37176 15534 37188
rect 15626 37179 15684 37185
rect 15626 37176 15638 37179
rect 15528 37148 15638 37176
rect 15528 37136 15534 37148
rect 15626 37145 15638 37148
rect 15672 37145 15684 37179
rect 15626 37139 15684 37145
rect 17310 37136 17316 37188
rect 17368 37176 17374 37188
rect 17880 37176 17908 37207
rect 17368 37148 17908 37176
rect 17368 37136 17374 37148
rect 19444 37108 19472 37207
rect 20254 37204 20260 37216
rect 20312 37204 20318 37256
rect 21821 37247 21879 37253
rect 21821 37213 21833 37247
rect 21867 37244 21879 37247
rect 22002 37244 22008 37256
rect 21867 37216 22008 37244
rect 21867 37213 21879 37216
rect 21821 37207 21879 37213
rect 22002 37204 22008 37216
rect 22060 37204 22066 37256
rect 23017 37247 23075 37253
rect 23017 37244 23029 37247
rect 22296 37216 23029 37244
rect 19610 37176 19616 37188
rect 19523 37148 19616 37176
rect 19610 37136 19616 37148
rect 19668 37176 19674 37188
rect 20438 37176 20444 37188
rect 19668 37148 20444 37176
rect 19668 37136 19674 37148
rect 20438 37136 20444 37148
rect 20496 37136 20502 37188
rect 20530 37136 20536 37188
rect 20588 37176 20594 37188
rect 21554 37179 21612 37185
rect 21554 37176 21566 37179
rect 20588 37148 21566 37176
rect 20588 37136 20594 37148
rect 21554 37145 21566 37148
rect 21600 37145 21612 37179
rect 21554 37139 21612 37145
rect 22296 37120 22324 37216
rect 23017 37213 23029 37216
rect 23063 37213 23075 37247
rect 23017 37207 23075 37213
rect 23109 37247 23167 37253
rect 23109 37213 23121 37247
rect 23155 37244 23167 37247
rect 23155 37216 23336 37244
rect 23155 37213 23167 37216
rect 23109 37207 23167 37213
rect 23201 37179 23259 37185
rect 23201 37145 23213 37179
rect 23247 37145 23259 37179
rect 23308 37176 23336 37216
rect 23382 37204 23388 37256
rect 23440 37244 23446 37256
rect 23440 37216 23485 37244
rect 23440 37204 23446 37216
rect 24762 37204 24768 37256
rect 24820 37244 24826 37256
rect 24949 37247 25007 37253
rect 24949 37244 24961 37247
rect 24820 37216 24961 37244
rect 24820 37204 24826 37216
rect 24949 37213 24961 37216
rect 24995 37213 25007 37247
rect 24949 37207 25007 37213
rect 30561 37247 30619 37253
rect 30561 37213 30573 37247
rect 30607 37244 30619 37247
rect 31662 37244 31668 37256
rect 30607 37216 31668 37244
rect 30607 37213 30619 37216
rect 30561 37207 30619 37213
rect 31662 37204 31668 37216
rect 31720 37204 31726 37256
rect 32306 37204 32312 37256
rect 32364 37244 32370 37256
rect 32401 37247 32459 37253
rect 32401 37244 32413 37247
rect 32364 37216 32413 37244
rect 32364 37204 32370 37216
rect 32401 37213 32413 37216
rect 32447 37213 32459 37247
rect 32401 37207 32459 37213
rect 33502 37204 33508 37256
rect 33560 37244 33566 37256
rect 34701 37247 34759 37253
rect 34701 37244 34713 37247
rect 33560 37216 34713 37244
rect 33560 37204 33566 37216
rect 34701 37213 34713 37216
rect 34747 37213 34759 37247
rect 34701 37207 34759 37213
rect 34885 37247 34943 37253
rect 34885 37213 34897 37247
rect 34931 37213 34943 37247
rect 34885 37207 34943 37213
rect 34977 37247 35035 37253
rect 34977 37213 34989 37247
rect 35023 37213 35035 37247
rect 34977 37207 35035 37213
rect 35069 37247 35127 37253
rect 35069 37213 35081 37247
rect 35115 37244 35127 37247
rect 35618 37244 35624 37256
rect 35115 37216 35624 37244
rect 35115 37213 35127 37216
rect 35069 37207 35127 37213
rect 24578 37176 24584 37188
rect 23308 37148 24584 37176
rect 23201 37139 23259 37145
rect 15396 37080 19472 37108
rect 19981 37111 20039 37117
rect 19981 37077 19993 37111
rect 20027 37108 20039 37111
rect 20622 37108 20628 37120
rect 20027 37080 20628 37108
rect 20027 37077 20039 37080
rect 19981 37071 20039 37077
rect 20622 37068 20628 37080
rect 20680 37068 20686 37120
rect 22278 37108 22284 37120
rect 22239 37080 22284 37108
rect 22278 37068 22284 37080
rect 22336 37068 22342 37120
rect 22833 37111 22891 37117
rect 22833 37077 22845 37111
rect 22879 37108 22891 37111
rect 22922 37108 22928 37120
rect 22879 37080 22928 37108
rect 22879 37077 22891 37080
rect 22833 37071 22891 37077
rect 22922 37068 22928 37080
rect 22980 37068 22986 37120
rect 23014 37068 23020 37120
rect 23072 37108 23078 37120
rect 23216 37108 23244 37139
rect 24578 37136 24584 37148
rect 24636 37136 24642 37188
rect 25038 37136 25044 37188
rect 25096 37176 25102 37188
rect 25194 37179 25252 37185
rect 25194 37176 25206 37179
rect 25096 37148 25206 37176
rect 25096 37136 25102 37148
rect 25194 37145 25206 37148
rect 25240 37145 25252 37179
rect 25194 37139 25252 37145
rect 30828 37179 30886 37185
rect 30828 37145 30840 37179
rect 30874 37176 30886 37179
rect 30926 37176 30932 37188
rect 30874 37148 30932 37176
rect 30874 37145 30886 37148
rect 30828 37139 30886 37145
rect 30926 37136 30932 37148
rect 30984 37136 30990 37188
rect 34146 37136 34152 37188
rect 34204 37176 34210 37188
rect 34900 37176 34928 37207
rect 34204 37148 34928 37176
rect 34204 37136 34210 37148
rect 23072 37080 23244 37108
rect 23072 37068 23078 37080
rect 24486 37068 24492 37120
rect 24544 37108 24550 37120
rect 26329 37111 26387 37117
rect 26329 37108 26341 37111
rect 24544 37080 26341 37108
rect 24544 37068 24550 37080
rect 26329 37077 26341 37080
rect 26375 37077 26387 37111
rect 26329 37071 26387 37077
rect 28166 37068 28172 37120
rect 28224 37108 28230 37120
rect 28905 37111 28963 37117
rect 28905 37108 28917 37111
rect 28224 37080 28917 37108
rect 28224 37068 28230 37080
rect 28905 37077 28917 37080
rect 28951 37108 28963 37111
rect 29270 37108 29276 37120
rect 28951 37080 29276 37108
rect 28951 37077 28963 37080
rect 28905 37071 28963 37077
rect 29270 37068 29276 37080
rect 29328 37068 29334 37120
rect 29638 37108 29644 37120
rect 29599 37080 29644 37108
rect 29638 37068 29644 37080
rect 29696 37068 29702 37120
rect 31938 37108 31944 37120
rect 31899 37080 31944 37108
rect 31938 37068 31944 37080
rect 31996 37068 32002 37120
rect 33870 37068 33876 37120
rect 33928 37108 33934 37120
rect 34992 37108 35020 37207
rect 35618 37204 35624 37216
rect 35676 37204 35682 37256
rect 35342 37108 35348 37120
rect 33928 37080 35020 37108
rect 35303 37080 35348 37108
rect 33928 37068 33934 37080
rect 35342 37068 35348 37080
rect 35400 37068 35406 37120
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 7650 36904 7656 36916
rect 6656 36876 7656 36904
rect 2590 36796 2596 36848
rect 2648 36836 2654 36848
rect 3145 36839 3203 36845
rect 3145 36836 3157 36839
rect 2648 36808 3157 36836
rect 2648 36796 2654 36808
rect 3145 36805 3157 36808
rect 3191 36805 3203 36839
rect 3145 36799 3203 36805
rect 5166 36796 5172 36848
rect 5224 36836 5230 36848
rect 5224 36808 6592 36836
rect 5224 36796 5230 36808
rect 6564 36777 6592 36808
rect 4893 36771 4951 36777
rect 4893 36737 4905 36771
rect 4939 36768 4951 36771
rect 6549 36771 6607 36777
rect 4939 36740 5488 36768
rect 4939 36737 4951 36740
rect 4893 36731 4951 36737
rect 5460 36641 5488 36740
rect 6549 36737 6561 36771
rect 6595 36737 6607 36771
rect 6656 36768 6684 36876
rect 7650 36864 7656 36876
rect 7708 36904 7714 36916
rect 12526 36904 12532 36916
rect 7708 36876 12532 36904
rect 7708 36864 7714 36876
rect 12526 36864 12532 36876
rect 12584 36864 12590 36916
rect 14553 36907 14611 36913
rect 14553 36873 14565 36907
rect 14599 36904 14611 36907
rect 14642 36904 14648 36916
rect 14599 36876 14648 36904
rect 14599 36873 14611 36876
rect 14553 36867 14611 36873
rect 14642 36864 14648 36876
rect 14700 36864 14706 36916
rect 15470 36904 15476 36916
rect 15431 36876 15476 36904
rect 15470 36864 15476 36876
rect 15528 36864 15534 36916
rect 17770 36864 17776 36916
rect 17828 36904 17834 36916
rect 18141 36907 18199 36913
rect 18141 36904 18153 36907
rect 17828 36876 18153 36904
rect 17828 36864 17834 36876
rect 18141 36873 18153 36876
rect 18187 36873 18199 36907
rect 18141 36867 18199 36873
rect 18693 36907 18751 36913
rect 18693 36873 18705 36907
rect 18739 36904 18751 36907
rect 18966 36904 18972 36916
rect 18739 36876 18972 36904
rect 18739 36873 18751 36876
rect 18693 36867 18751 36873
rect 18966 36864 18972 36876
rect 19024 36864 19030 36916
rect 20441 36907 20499 36913
rect 20441 36873 20453 36907
rect 20487 36904 20499 36907
rect 20530 36904 20536 36916
rect 20487 36876 20536 36904
rect 20487 36873 20499 36876
rect 20441 36867 20499 36873
rect 20530 36864 20536 36876
rect 20588 36864 20594 36916
rect 24762 36864 24768 36916
rect 24820 36904 24826 36916
rect 24949 36907 25007 36913
rect 24949 36904 24961 36907
rect 24820 36876 24961 36904
rect 24820 36864 24826 36876
rect 24949 36873 24961 36876
rect 24995 36873 25007 36907
rect 24949 36867 25007 36873
rect 29917 36907 29975 36913
rect 29917 36873 29929 36907
rect 29963 36904 29975 36907
rect 30374 36904 30380 36916
rect 29963 36876 30380 36904
rect 29963 36873 29975 36876
rect 29917 36867 29975 36873
rect 30374 36864 30380 36876
rect 30432 36864 30438 36916
rect 32582 36904 32588 36916
rect 32543 36876 32588 36904
rect 32582 36864 32588 36876
rect 32640 36864 32646 36916
rect 33410 36904 33416 36916
rect 32876 36876 33416 36904
rect 6822 36836 6828 36848
rect 6783 36808 6828 36836
rect 6822 36796 6828 36808
rect 6880 36796 6886 36848
rect 7466 36796 7472 36848
rect 7524 36836 7530 36848
rect 7745 36839 7803 36845
rect 7745 36836 7757 36839
rect 7524 36808 7757 36836
rect 7524 36796 7530 36808
rect 7745 36805 7757 36808
rect 7791 36805 7803 36839
rect 7745 36799 7803 36805
rect 13188 36808 14228 36836
rect 6733 36771 6791 36777
rect 6733 36768 6745 36771
rect 6656 36740 6745 36768
rect 6549 36731 6607 36737
rect 6733 36737 6745 36740
rect 6779 36737 6791 36771
rect 6733 36731 6791 36737
rect 6917 36771 6975 36777
rect 6917 36737 6929 36771
rect 6963 36768 6975 36771
rect 7834 36768 7840 36780
rect 6963 36740 7840 36768
rect 6963 36737 6975 36740
rect 6917 36731 6975 36737
rect 7834 36728 7840 36740
rect 7892 36728 7898 36780
rect 7926 36728 7932 36780
rect 7984 36768 7990 36780
rect 7984 36740 8029 36768
rect 7984 36728 7990 36740
rect 9766 36728 9772 36780
rect 9824 36768 9830 36780
rect 13188 36777 13216 36808
rect 12069 36771 12127 36777
rect 12069 36768 12081 36771
rect 9824 36740 12081 36768
rect 9824 36728 9830 36740
rect 12069 36737 12081 36740
rect 12115 36737 12127 36771
rect 12069 36731 12127 36737
rect 13173 36771 13231 36777
rect 13173 36737 13185 36771
rect 13219 36737 13231 36771
rect 13173 36731 13231 36737
rect 13440 36771 13498 36777
rect 13440 36737 13452 36771
rect 13486 36768 13498 36771
rect 13998 36768 14004 36780
rect 13486 36740 14004 36768
rect 13486 36737 13498 36740
rect 13440 36731 13498 36737
rect 13998 36728 14004 36740
rect 14056 36728 14062 36780
rect 14200 36768 14228 36808
rect 16758 36796 16764 36848
rect 16816 36836 16822 36848
rect 16853 36839 16911 36845
rect 16853 36836 16865 36839
rect 16816 36808 16865 36836
rect 16816 36796 16822 36808
rect 16853 36805 16865 36808
rect 16899 36805 16911 36839
rect 16853 36799 16911 36805
rect 17957 36839 18015 36845
rect 17957 36805 17969 36839
rect 18003 36836 18015 36839
rect 19426 36836 19432 36848
rect 18003 36808 19432 36836
rect 18003 36805 18015 36808
rect 17957 36799 18015 36805
rect 19426 36796 19432 36808
rect 19484 36796 19490 36848
rect 23661 36839 23719 36845
rect 19720 36808 20208 36836
rect 15378 36768 15384 36780
rect 14200 36740 15384 36768
rect 15378 36728 15384 36740
rect 15436 36728 15442 36780
rect 15726 36768 15732 36780
rect 15687 36740 15732 36768
rect 15726 36728 15732 36740
rect 15784 36728 15790 36780
rect 15841 36771 15899 36777
rect 15841 36737 15853 36771
rect 15887 36737 15899 36771
rect 15841 36731 15899 36737
rect 15933 36774 15991 36780
rect 15933 36740 15945 36774
rect 15979 36740 15991 36774
rect 15933 36734 15991 36740
rect 15856 36644 15884 36731
rect 15948 36700 15976 36734
rect 16114 36728 16120 36780
rect 16172 36768 16178 36780
rect 17034 36768 17040 36780
rect 16172 36740 16217 36768
rect 16995 36740 17040 36768
rect 16172 36728 16178 36740
rect 17034 36728 17040 36740
rect 17092 36768 17098 36780
rect 17773 36771 17831 36777
rect 17773 36768 17785 36771
rect 17092 36740 17785 36768
rect 17092 36728 17098 36740
rect 17773 36737 17785 36740
rect 17819 36737 17831 36771
rect 17773 36731 17831 36737
rect 17862 36728 17868 36780
rect 17920 36768 17926 36780
rect 19720 36768 19748 36808
rect 17920 36740 19748 36768
rect 17920 36728 17926 36740
rect 19794 36728 19800 36780
rect 19852 36768 19858 36780
rect 19978 36768 19984 36780
rect 19852 36740 19897 36768
rect 19939 36740 19984 36768
rect 19852 36728 19858 36740
rect 19978 36728 19984 36740
rect 20036 36728 20042 36780
rect 20180 36777 20208 36808
rect 23661 36805 23673 36839
rect 23707 36836 23719 36839
rect 25961 36839 26019 36845
rect 25961 36836 25973 36839
rect 23707 36808 25973 36836
rect 23707 36805 23719 36808
rect 23661 36799 23719 36805
rect 25961 36805 25973 36808
rect 26007 36836 26019 36839
rect 28810 36836 28816 36848
rect 26007 36808 28816 36836
rect 26007 36805 26019 36808
rect 25961 36799 26019 36805
rect 28810 36796 28816 36808
rect 28868 36796 28874 36848
rect 32876 36836 32904 36876
rect 33410 36864 33416 36876
rect 33468 36864 33474 36916
rect 35434 36864 35440 36916
rect 35492 36904 35498 36916
rect 36265 36907 36323 36913
rect 36265 36904 36277 36907
rect 35492 36876 36277 36904
rect 35492 36864 35498 36876
rect 36265 36873 36277 36876
rect 36311 36873 36323 36907
rect 36265 36867 36323 36873
rect 33870 36836 33876 36848
rect 28966 36808 32904 36836
rect 20073 36771 20131 36777
rect 20073 36737 20085 36771
rect 20119 36737 20131 36771
rect 20073 36731 20131 36737
rect 20165 36771 20223 36777
rect 20165 36737 20177 36771
rect 20211 36768 20223 36771
rect 20901 36771 20959 36777
rect 20901 36768 20913 36771
rect 20211 36740 20913 36768
rect 20211 36737 20223 36740
rect 20165 36731 20223 36737
rect 20901 36737 20913 36740
rect 20947 36737 20959 36771
rect 20901 36731 20959 36737
rect 15948 36672 16712 36700
rect 5445 36635 5503 36641
rect 5445 36601 5457 36635
rect 5491 36632 5503 36635
rect 8294 36632 8300 36644
rect 5491 36604 8300 36632
rect 5491 36601 5503 36604
rect 5445 36595 5503 36601
rect 8294 36592 8300 36604
rect 8352 36592 8358 36644
rect 15838 36592 15844 36644
rect 15896 36592 15902 36644
rect 16684 36641 16712 36672
rect 18690 36660 18696 36712
rect 18748 36700 18754 36712
rect 19242 36700 19248 36712
rect 18748 36672 19248 36700
rect 18748 36660 18754 36672
rect 19242 36660 19248 36672
rect 19300 36700 19306 36712
rect 20088 36700 20116 36731
rect 19300 36672 20116 36700
rect 19300 36660 19306 36672
rect 16669 36635 16727 36641
rect 16669 36601 16681 36635
rect 16715 36601 16727 36635
rect 16669 36595 16727 36601
rect 19978 36592 19984 36644
rect 20036 36632 20042 36644
rect 20254 36632 20260 36644
rect 20036 36604 20260 36632
rect 20036 36592 20042 36604
rect 20254 36592 20260 36604
rect 20312 36592 20318 36644
rect 20916 36632 20944 36731
rect 22278 36728 22284 36780
rect 22336 36768 22342 36780
rect 22833 36771 22891 36777
rect 22833 36768 22845 36771
rect 22336 36740 22845 36768
rect 22336 36728 22342 36740
rect 22833 36737 22845 36740
rect 22879 36737 22891 36771
rect 22833 36731 22891 36737
rect 22925 36771 22983 36777
rect 22925 36737 22937 36771
rect 22971 36737 22983 36771
rect 22925 36731 22983 36737
rect 22940 36700 22968 36731
rect 23014 36728 23020 36780
rect 23072 36768 23078 36780
rect 23201 36771 23259 36777
rect 23072 36740 23117 36768
rect 23072 36728 23078 36740
rect 23201 36737 23213 36771
rect 23247 36768 23259 36771
rect 23566 36768 23572 36780
rect 23247 36740 23572 36768
rect 23247 36737 23259 36740
rect 23201 36731 23259 36737
rect 23566 36728 23572 36740
rect 23624 36728 23630 36780
rect 27430 36768 27436 36780
rect 27391 36740 27436 36768
rect 27430 36728 27436 36740
rect 27488 36728 27494 36780
rect 27522 36728 27528 36780
rect 27580 36768 27586 36780
rect 27689 36771 27747 36777
rect 27689 36768 27701 36771
rect 27580 36740 27701 36768
rect 27580 36728 27586 36740
rect 27689 36737 27701 36740
rect 27735 36737 27747 36771
rect 27689 36731 27747 36737
rect 27982 36728 27988 36780
rect 28040 36768 28046 36780
rect 28966 36768 28994 36808
rect 29270 36768 29276 36780
rect 28040 36740 28994 36768
rect 29231 36740 29276 36768
rect 28040 36728 28046 36740
rect 29270 36728 29276 36740
rect 29328 36728 29334 36780
rect 29454 36768 29460 36780
rect 29415 36740 29460 36768
rect 29454 36728 29460 36740
rect 29512 36728 29518 36780
rect 29549 36771 29607 36777
rect 29549 36737 29561 36771
rect 29595 36737 29607 36771
rect 29549 36731 29607 36737
rect 24486 36700 24492 36712
rect 22940 36672 24492 36700
rect 24486 36660 24492 36672
rect 24544 36660 24550 36712
rect 28994 36660 29000 36712
rect 29052 36700 29058 36712
rect 29564 36700 29592 36731
rect 29638 36728 29644 36780
rect 29696 36768 29702 36780
rect 29696 36740 29741 36768
rect 29696 36728 29702 36740
rect 30282 36728 30288 36780
rect 30340 36768 30346 36780
rect 32876 36777 32904 36808
rect 32968 36808 33876 36836
rect 32968 36777 32996 36808
rect 33870 36796 33876 36808
rect 33928 36836 33934 36848
rect 34425 36839 34483 36845
rect 33928 36808 34100 36836
rect 33928 36796 33934 36808
rect 31113 36771 31171 36777
rect 31113 36768 31125 36771
rect 30340 36740 31125 36768
rect 30340 36728 30346 36740
rect 31113 36737 31125 36740
rect 31159 36768 31171 36771
rect 32861 36771 32919 36777
rect 31159 36740 31754 36768
rect 31159 36737 31171 36740
rect 31113 36731 31171 36737
rect 31386 36700 31392 36712
rect 29052 36672 29592 36700
rect 31347 36672 31392 36700
rect 29052 36660 29058 36672
rect 31386 36660 31392 36672
rect 31444 36660 31450 36712
rect 31726 36700 31754 36740
rect 32861 36737 32873 36771
rect 32907 36737 32919 36771
rect 32861 36731 32919 36737
rect 32953 36771 33011 36777
rect 32953 36737 32965 36771
rect 32999 36737 33011 36771
rect 32953 36731 33011 36737
rect 33045 36771 33103 36777
rect 33045 36737 33057 36771
rect 33091 36768 33103 36771
rect 33134 36768 33140 36780
rect 33091 36740 33140 36768
rect 33091 36737 33103 36740
rect 33045 36731 33103 36737
rect 33134 36728 33140 36740
rect 33192 36728 33198 36780
rect 33229 36771 33287 36777
rect 33229 36737 33241 36771
rect 33275 36737 33287 36771
rect 33229 36731 33287 36737
rect 33244 36700 33272 36731
rect 33502 36728 33508 36780
rect 33560 36768 33566 36780
rect 34072 36777 34100 36808
rect 34425 36805 34437 36839
rect 34471 36836 34483 36839
rect 35130 36839 35188 36845
rect 35130 36836 35142 36839
rect 34471 36808 35142 36836
rect 34471 36805 34483 36808
rect 34425 36799 34483 36805
rect 35130 36805 35142 36808
rect 35176 36805 35188 36839
rect 35130 36799 35188 36805
rect 33781 36771 33839 36777
rect 33781 36768 33793 36771
rect 33560 36740 33793 36768
rect 33560 36728 33566 36740
rect 33781 36737 33793 36740
rect 33827 36737 33839 36771
rect 33781 36731 33839 36737
rect 33965 36771 34023 36777
rect 33965 36737 33977 36771
rect 34011 36737 34023 36771
rect 33965 36731 34023 36737
rect 34057 36771 34115 36777
rect 34057 36737 34069 36771
rect 34103 36737 34115 36771
rect 34057 36731 34115 36737
rect 34149 36771 34207 36777
rect 34149 36737 34161 36771
rect 34195 36768 34207 36771
rect 34238 36768 34244 36780
rect 34195 36740 34244 36768
rect 34195 36737 34207 36740
rect 34149 36731 34207 36737
rect 31726 36672 33272 36700
rect 33980 36700 34008 36731
rect 34238 36728 34244 36740
rect 34296 36728 34302 36780
rect 34882 36768 34888 36780
rect 34843 36740 34888 36768
rect 34882 36728 34888 36740
rect 34940 36728 34946 36780
rect 34698 36700 34704 36712
rect 33980 36672 34704 36700
rect 34698 36660 34704 36672
rect 34756 36660 34762 36712
rect 25222 36632 25228 36644
rect 20916 36604 25228 36632
rect 25222 36592 25228 36604
rect 25280 36592 25286 36644
rect 7098 36564 7104 36576
rect 7059 36536 7104 36564
rect 7098 36524 7104 36536
rect 7156 36524 7162 36576
rect 7466 36524 7472 36576
rect 7524 36564 7530 36576
rect 7561 36567 7619 36573
rect 7561 36564 7573 36567
rect 7524 36536 7573 36564
rect 7524 36524 7530 36536
rect 7561 36533 7573 36536
rect 7607 36533 7619 36567
rect 7561 36527 7619 36533
rect 12161 36567 12219 36573
rect 12161 36533 12173 36567
rect 12207 36564 12219 36567
rect 15470 36564 15476 36576
rect 12207 36536 15476 36564
rect 12207 36533 12219 36536
rect 12161 36527 12219 36533
rect 15470 36524 15476 36536
rect 15528 36564 15534 36576
rect 16114 36564 16120 36576
rect 15528 36536 16120 36564
rect 15528 36524 15534 36536
rect 16114 36524 16120 36536
rect 16172 36564 16178 36576
rect 17586 36564 17592 36576
rect 16172 36536 17592 36564
rect 16172 36524 16178 36536
rect 17586 36524 17592 36536
rect 17644 36524 17650 36576
rect 19337 36567 19395 36573
rect 19337 36533 19349 36567
rect 19383 36564 19395 36567
rect 19426 36564 19432 36576
rect 19383 36536 19432 36564
rect 19383 36533 19395 36536
rect 19337 36527 19395 36533
rect 19426 36524 19432 36536
rect 19484 36564 19490 36576
rect 19794 36564 19800 36576
rect 19484 36536 19800 36564
rect 19484 36524 19490 36536
rect 19794 36524 19800 36536
rect 19852 36564 19858 36576
rect 20346 36564 20352 36576
rect 19852 36536 20352 36564
rect 19852 36524 19858 36536
rect 20346 36524 20352 36536
rect 20404 36524 20410 36576
rect 22189 36567 22247 36573
rect 22189 36533 22201 36567
rect 22235 36564 22247 36567
rect 22278 36564 22284 36576
rect 22235 36536 22284 36564
rect 22235 36533 22247 36536
rect 22189 36527 22247 36533
rect 22278 36524 22284 36536
rect 22336 36524 22342 36576
rect 22646 36564 22652 36576
rect 22607 36536 22652 36564
rect 22646 36524 22652 36536
rect 22704 36524 22710 36576
rect 28442 36524 28448 36576
rect 28500 36564 28506 36576
rect 28813 36567 28871 36573
rect 28813 36564 28825 36567
rect 28500 36536 28825 36564
rect 28500 36524 28506 36536
rect 28813 36533 28825 36536
rect 28859 36533 28871 36567
rect 28813 36527 28871 36533
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 5166 36360 5172 36372
rect 5127 36332 5172 36360
rect 5166 36320 5172 36332
rect 5224 36320 5230 36372
rect 7006 36360 7012 36372
rect 6967 36332 7012 36360
rect 7006 36320 7012 36332
rect 7064 36320 7070 36372
rect 9677 36363 9735 36369
rect 9677 36329 9689 36363
rect 9723 36360 9735 36363
rect 11054 36360 11060 36372
rect 9723 36332 11060 36360
rect 9723 36329 9735 36332
rect 9677 36323 9735 36329
rect 11054 36320 11060 36332
rect 11112 36320 11118 36372
rect 12526 36360 12532 36372
rect 12487 36332 12532 36360
rect 12526 36320 12532 36332
rect 12584 36320 12590 36372
rect 13998 36320 14004 36372
rect 14056 36360 14062 36372
rect 14093 36363 14151 36369
rect 14093 36360 14105 36363
rect 14056 36332 14105 36360
rect 14056 36320 14062 36332
rect 14093 36329 14105 36332
rect 14139 36329 14151 36363
rect 14093 36323 14151 36329
rect 14366 36320 14372 36372
rect 14424 36360 14430 36372
rect 15102 36360 15108 36372
rect 14424 36332 15108 36360
rect 14424 36320 14430 36332
rect 15102 36320 15108 36332
rect 15160 36360 15166 36372
rect 15197 36363 15255 36369
rect 15197 36360 15209 36363
rect 15160 36332 15209 36360
rect 15160 36320 15166 36332
rect 15197 36329 15209 36332
rect 15243 36329 15255 36363
rect 15197 36323 15255 36329
rect 15746 36320 15752 36372
rect 15804 36360 15810 36372
rect 16298 36360 16304 36372
rect 15804 36332 16304 36360
rect 15804 36320 15810 36332
rect 16298 36320 16304 36332
rect 16356 36320 16362 36372
rect 27062 36360 27068 36372
rect 27023 36332 27068 36360
rect 27062 36320 27068 36332
rect 27120 36320 27126 36372
rect 27522 36360 27528 36372
rect 27483 36332 27528 36360
rect 27522 36320 27528 36332
rect 27580 36320 27586 36372
rect 29454 36320 29460 36372
rect 29512 36360 29518 36372
rect 29549 36363 29607 36369
rect 29549 36360 29561 36363
rect 29512 36332 29561 36360
rect 29512 36320 29518 36332
rect 29549 36329 29561 36332
rect 29595 36329 29607 36363
rect 34146 36360 34152 36372
rect 34107 36332 34152 36360
rect 29549 36323 29607 36329
rect 34146 36320 34152 36332
rect 34204 36320 34210 36372
rect 34698 36320 34704 36372
rect 34756 36360 34762 36372
rect 35069 36363 35127 36369
rect 35069 36360 35081 36363
rect 34756 36332 35081 36360
rect 34756 36320 34762 36332
rect 35069 36329 35081 36332
rect 35115 36329 35127 36363
rect 35069 36323 35127 36329
rect 23658 36252 23664 36304
rect 23716 36292 23722 36304
rect 25133 36295 25191 36301
rect 25133 36292 25145 36295
rect 23716 36264 25145 36292
rect 23716 36252 23722 36264
rect 25133 36261 25145 36264
rect 25179 36261 25191 36295
rect 25133 36255 25191 36261
rect 28810 36252 28816 36304
rect 28868 36292 28874 36304
rect 32306 36292 32312 36304
rect 28868 36264 32312 36292
rect 28868 36252 28874 36264
rect 32306 36252 32312 36264
rect 32364 36252 32370 36304
rect 2590 36184 2596 36236
rect 2648 36224 2654 36236
rect 3789 36227 3847 36233
rect 3789 36224 3801 36227
rect 2648 36196 3801 36224
rect 2648 36184 2654 36196
rect 3789 36193 3801 36196
rect 3835 36193 3847 36227
rect 3789 36187 3847 36193
rect 5350 36184 5356 36236
rect 5408 36224 5414 36236
rect 5408 36196 7417 36224
rect 5408 36184 5414 36196
rect 7285 36159 7343 36165
rect 7389 36159 7417 36196
rect 20990 36184 20996 36236
rect 21048 36224 21054 36236
rect 26513 36227 26571 36233
rect 21048 36196 22692 36224
rect 21048 36184 21054 36196
rect 7285 36125 7297 36159
rect 7331 36125 7343 36159
rect 7285 36119 7343 36125
rect 7374 36153 7432 36159
rect 7374 36119 7386 36153
rect 7420 36119 7432 36153
rect 4056 36091 4114 36097
rect 4056 36057 4068 36091
rect 4102 36088 4114 36091
rect 4614 36088 4620 36100
rect 4102 36060 4620 36088
rect 4102 36057 4114 36060
rect 4056 36051 4114 36057
rect 4614 36048 4620 36060
rect 4672 36048 4678 36100
rect 6549 36023 6607 36029
rect 6549 35989 6561 36023
rect 6595 36020 6607 36023
rect 6638 36020 6644 36032
rect 6595 35992 6644 36020
rect 6595 35989 6607 35992
rect 6549 35983 6607 35989
rect 6638 35980 6644 35992
rect 6696 36020 6702 36032
rect 7300 36020 7328 36119
rect 7374 36113 7432 36119
rect 7466 36116 7472 36168
rect 7524 36156 7530 36168
rect 7653 36159 7711 36165
rect 7524 36128 7569 36156
rect 7524 36116 7530 36128
rect 7653 36125 7665 36159
rect 7699 36125 7711 36159
rect 7653 36119 7711 36125
rect 6696 35992 7328 36020
rect 7389 36020 7417 36113
rect 7668 36088 7696 36119
rect 9306 36116 9312 36168
rect 9364 36156 9370 36168
rect 9493 36159 9551 36165
rect 9493 36156 9505 36159
rect 9364 36128 9505 36156
rect 9364 36116 9370 36128
rect 9493 36125 9505 36128
rect 9539 36125 9551 36159
rect 9493 36119 9551 36125
rect 10137 36159 10195 36165
rect 10137 36125 10149 36159
rect 10183 36156 10195 36159
rect 10226 36156 10232 36168
rect 10183 36128 10232 36156
rect 10183 36125 10195 36128
rect 10137 36119 10195 36125
rect 10226 36116 10232 36128
rect 10284 36116 10290 36168
rect 14366 36156 14372 36168
rect 14327 36128 14372 36156
rect 14366 36116 14372 36128
rect 14424 36116 14430 36168
rect 14461 36159 14519 36165
rect 14461 36125 14473 36159
rect 14507 36125 14519 36159
rect 14461 36119 14519 36125
rect 10410 36097 10416 36100
rect 7668 36060 10180 36088
rect 10152 36032 10180 36060
rect 10404 36051 10416 36097
rect 10468 36088 10474 36100
rect 12621 36091 12679 36097
rect 10468 36060 10504 36088
rect 10410 36048 10416 36051
rect 10468 36048 10474 36060
rect 12621 36057 12633 36091
rect 12667 36088 12679 36091
rect 13078 36088 13084 36100
rect 12667 36060 13084 36088
rect 12667 36057 12679 36060
rect 12621 36051 12679 36057
rect 13078 36048 13084 36060
rect 13136 36048 13142 36100
rect 13354 36088 13360 36100
rect 13315 36060 13360 36088
rect 13354 36048 13360 36060
rect 13412 36088 13418 36100
rect 13814 36088 13820 36100
rect 13412 36060 13820 36088
rect 13412 36048 13418 36060
rect 13814 36048 13820 36060
rect 13872 36048 13878 36100
rect 14274 36048 14280 36100
rect 14332 36088 14338 36100
rect 14476 36088 14504 36119
rect 14550 36116 14556 36168
rect 14608 36156 14614 36168
rect 14608 36128 14653 36156
rect 14608 36116 14614 36128
rect 14734 36116 14740 36168
rect 14792 36156 14798 36168
rect 22278 36156 22284 36168
rect 14792 36128 14837 36156
rect 22239 36128 22284 36156
rect 14792 36116 14798 36128
rect 22278 36116 22284 36128
rect 22336 36116 22342 36168
rect 22664 36165 22692 36196
rect 26513 36193 26525 36227
rect 26559 36224 26571 36227
rect 27430 36224 27436 36236
rect 26559 36196 27436 36224
rect 26559 36193 26571 36196
rect 26513 36187 26571 36193
rect 27430 36184 27436 36196
rect 27488 36184 27494 36236
rect 28629 36227 28687 36233
rect 28629 36224 28641 36227
rect 28000 36196 28641 36224
rect 22649 36159 22707 36165
rect 22649 36125 22661 36159
rect 22695 36125 22707 36159
rect 23474 36156 23480 36168
rect 23435 36128 23480 36156
rect 22649 36119 22707 36125
rect 23474 36116 23480 36128
rect 23532 36116 23538 36168
rect 23661 36159 23719 36165
rect 23661 36125 23673 36159
rect 23707 36156 23719 36159
rect 24486 36156 24492 36168
rect 23707 36128 24492 36156
rect 23707 36125 23719 36128
rect 23661 36119 23719 36125
rect 24486 36116 24492 36128
rect 24544 36116 24550 36168
rect 27062 36116 27068 36168
rect 27120 36156 27126 36168
rect 28000 36165 28028 36196
rect 28629 36193 28641 36196
rect 28675 36193 28687 36227
rect 28629 36187 28687 36193
rect 34790 36184 34796 36236
rect 34848 36224 34854 36236
rect 35621 36227 35679 36233
rect 35621 36224 35633 36227
rect 34848 36196 35633 36224
rect 34848 36184 34854 36196
rect 35621 36193 35633 36196
rect 35667 36193 35679 36227
rect 35621 36187 35679 36193
rect 27801 36159 27859 36165
rect 27801 36156 27813 36159
rect 27120 36128 27813 36156
rect 27120 36116 27126 36128
rect 27801 36125 27813 36128
rect 27847 36125 27859 36159
rect 27801 36119 27859 36125
rect 27893 36159 27951 36165
rect 27893 36125 27905 36159
rect 27939 36125 27951 36159
rect 27893 36119 27951 36125
rect 27985 36159 28043 36165
rect 27985 36125 27997 36159
rect 28031 36125 28043 36159
rect 28166 36156 28172 36168
rect 28127 36128 28172 36156
rect 27985 36119 28043 36125
rect 15838 36088 15844 36100
rect 14332 36060 15844 36088
rect 14332 36048 14338 36060
rect 15838 36048 15844 36060
rect 15896 36088 15902 36100
rect 17310 36088 17316 36100
rect 15896 36060 17316 36088
rect 15896 36048 15902 36060
rect 17310 36048 17316 36060
rect 17368 36048 17374 36100
rect 22373 36091 22431 36097
rect 22373 36057 22385 36091
rect 22419 36057 22431 36091
rect 22373 36051 22431 36057
rect 22465 36091 22523 36097
rect 22465 36057 22477 36091
rect 22511 36088 22523 36091
rect 23014 36088 23020 36100
rect 22511 36060 23020 36088
rect 22511 36057 22523 36060
rect 22465 36051 22523 36057
rect 9490 36020 9496 36032
rect 7389 35992 9496 36020
rect 6696 35980 6702 35992
rect 9490 35980 9496 35992
rect 9548 35980 9554 36032
rect 10134 35980 10140 36032
rect 10192 35980 10198 36032
rect 11517 36023 11575 36029
rect 11517 35989 11529 36023
rect 11563 36020 11575 36023
rect 11698 36020 11704 36032
rect 11563 35992 11704 36020
rect 11563 35989 11575 35992
rect 11517 35983 11575 35989
rect 11698 35980 11704 35992
rect 11756 35980 11762 36032
rect 13449 36023 13507 36029
rect 13449 35989 13461 36023
rect 13495 36020 13507 36023
rect 13998 36020 14004 36032
rect 13495 35992 14004 36020
rect 13495 35989 13507 35992
rect 13449 35983 13507 35989
rect 13998 35980 14004 35992
rect 14056 35980 14062 36032
rect 22094 35980 22100 36032
rect 22152 36020 22158 36032
rect 22388 36020 22416 36051
rect 23014 36048 23020 36060
rect 23072 36048 23078 36100
rect 23842 36088 23848 36100
rect 23803 36060 23848 36088
rect 23842 36048 23848 36060
rect 23900 36048 23906 36100
rect 26234 36088 26240 36100
rect 26292 36097 26298 36100
rect 26204 36060 26240 36088
rect 26234 36048 26240 36060
rect 26292 36051 26304 36097
rect 26292 36048 26298 36051
rect 23658 36020 23664 36032
rect 22152 35992 22197 36020
rect 22388 35992 23664 36020
rect 22152 35980 22158 35992
rect 23658 35980 23664 35992
rect 23716 35980 23722 36032
rect 24394 36020 24400 36032
rect 24355 35992 24400 36020
rect 24394 35980 24400 35992
rect 24452 35980 24458 36032
rect 27908 36020 27936 36119
rect 28166 36116 28172 36128
rect 28224 36116 28230 36168
rect 28997 36159 29055 36165
rect 28997 36125 29009 36159
rect 29043 36156 29055 36159
rect 31386 36156 31392 36168
rect 29043 36128 29960 36156
rect 31299 36128 31392 36156
rect 29043 36125 29055 36128
rect 28997 36119 29055 36125
rect 28442 36048 28448 36100
rect 28500 36088 28506 36100
rect 28813 36091 28871 36097
rect 28813 36088 28825 36091
rect 28500 36060 28825 36088
rect 28500 36048 28506 36060
rect 28813 36057 28825 36060
rect 28859 36057 28871 36091
rect 28813 36051 28871 36057
rect 29454 36048 29460 36100
rect 29512 36088 29518 36100
rect 29932 36097 29960 36128
rect 31386 36116 31392 36128
rect 31444 36156 31450 36168
rect 31941 36159 31999 36165
rect 31941 36156 31953 36159
rect 31444 36128 31953 36156
rect 31444 36116 31450 36128
rect 31941 36125 31953 36128
rect 31987 36125 31999 36159
rect 31941 36119 31999 36125
rect 32217 36159 32275 36165
rect 32217 36125 32229 36159
rect 32263 36156 32275 36159
rect 33502 36156 33508 36168
rect 32263 36128 33508 36156
rect 32263 36125 32275 36128
rect 32217 36119 32275 36125
rect 33502 36116 33508 36128
rect 33560 36116 33566 36168
rect 34701 36159 34759 36165
rect 34701 36156 34713 36159
rect 33796 36128 34713 36156
rect 29733 36091 29791 36097
rect 29733 36088 29745 36091
rect 29512 36060 29745 36088
rect 29512 36048 29518 36060
rect 29733 36057 29745 36060
rect 29779 36057 29791 36091
rect 29733 36051 29791 36057
rect 29917 36091 29975 36097
rect 29917 36057 29929 36091
rect 29963 36088 29975 36091
rect 30466 36088 30472 36100
rect 29963 36060 30472 36088
rect 29963 36057 29975 36060
rect 29917 36051 29975 36057
rect 30466 36048 30472 36060
rect 30524 36048 30530 36100
rect 28994 36020 29000 36032
rect 27908 35992 29000 36020
rect 28994 35980 29000 35992
rect 29052 35980 29058 36032
rect 30374 36020 30380 36032
rect 30335 35992 30380 36020
rect 30374 35980 30380 35992
rect 30432 36020 30438 36032
rect 31404 36029 31432 36116
rect 33686 36048 33692 36100
rect 33744 36088 33750 36100
rect 33796 36097 33824 36128
rect 34701 36125 34713 36128
rect 34747 36125 34759 36159
rect 34701 36119 34759 36125
rect 35342 36116 35348 36168
rect 35400 36156 35406 36168
rect 35877 36159 35935 36165
rect 35877 36156 35889 36159
rect 35400 36128 35889 36156
rect 35400 36116 35406 36128
rect 35877 36125 35889 36128
rect 35923 36125 35935 36159
rect 58158 36156 58164 36168
rect 58119 36128 58164 36156
rect 35877 36119 35935 36125
rect 58158 36116 58164 36128
rect 58216 36116 58222 36168
rect 33781 36091 33839 36097
rect 33781 36088 33793 36091
rect 33744 36060 33793 36088
rect 33744 36048 33750 36060
rect 33781 36057 33793 36060
rect 33827 36057 33839 36091
rect 33781 36051 33839 36057
rect 33965 36091 34023 36097
rect 33965 36057 33977 36091
rect 34011 36057 34023 36091
rect 33965 36051 34023 36057
rect 34885 36091 34943 36097
rect 34885 36057 34897 36091
rect 34931 36088 34943 36091
rect 35434 36088 35440 36100
rect 34931 36060 35440 36088
rect 34931 36057 34943 36060
rect 34885 36051 34943 36057
rect 31389 36023 31447 36029
rect 31389 36020 31401 36023
rect 30432 35992 31401 36020
rect 30432 35980 30438 35992
rect 31389 35989 31401 35992
rect 31435 35989 31447 36023
rect 31389 35983 31447 35989
rect 33321 36023 33379 36029
rect 33321 35989 33333 36023
rect 33367 36020 33379 36023
rect 33410 36020 33416 36032
rect 33367 35992 33416 36020
rect 33367 35989 33379 35992
rect 33321 35983 33379 35989
rect 33410 35980 33416 35992
rect 33468 35980 33474 36032
rect 33980 36020 34008 36051
rect 35434 36048 35440 36060
rect 35492 36048 35498 36100
rect 34698 36020 34704 36032
rect 33980 35992 34704 36020
rect 34698 35980 34704 35992
rect 34756 36020 34762 36032
rect 37001 36023 37059 36029
rect 37001 36020 37013 36023
rect 34756 35992 37013 36020
rect 34756 35980 34762 35992
rect 37001 35989 37013 35992
rect 37047 35989 37059 36023
rect 37001 35983 37059 35989
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 12713 35819 12771 35825
rect 12713 35785 12725 35819
rect 12759 35816 12771 35819
rect 13354 35816 13360 35828
rect 12759 35788 13360 35816
rect 12759 35785 12771 35788
rect 12713 35779 12771 35785
rect 13354 35776 13360 35788
rect 13412 35776 13418 35828
rect 24670 35776 24676 35828
rect 24728 35816 24734 35828
rect 25133 35819 25191 35825
rect 24728 35788 24854 35816
rect 24728 35776 24734 35788
rect 4525 35751 4583 35757
rect 4525 35717 4537 35751
rect 4571 35748 4583 35751
rect 5166 35748 5172 35760
rect 4571 35720 5172 35748
rect 4571 35717 4583 35720
rect 4525 35711 4583 35717
rect 5166 35708 5172 35720
rect 5224 35708 5230 35760
rect 6104 35720 7604 35748
rect 2866 35640 2872 35692
rect 2924 35680 2930 35692
rect 4341 35683 4399 35689
rect 4341 35680 4353 35683
rect 2924 35652 4353 35680
rect 2924 35640 2930 35652
rect 4341 35649 4353 35652
rect 4387 35680 4399 35683
rect 6104 35680 6132 35720
rect 4387 35652 6132 35680
rect 4387 35649 4399 35652
rect 4341 35643 4399 35649
rect 7190 35640 7196 35692
rect 7248 35680 7254 35692
rect 7478 35683 7536 35689
rect 7478 35680 7490 35683
rect 7248 35652 7490 35680
rect 7248 35640 7254 35652
rect 7478 35649 7490 35652
rect 7524 35649 7536 35683
rect 7576 35680 7604 35720
rect 11054 35708 11060 35760
rect 11112 35748 11118 35760
rect 11514 35748 11520 35760
rect 11112 35720 11520 35748
rect 11112 35708 11118 35720
rect 11514 35708 11520 35720
rect 11572 35708 11578 35760
rect 13170 35748 13176 35760
rect 13131 35720 13176 35748
rect 13170 35708 13176 35720
rect 13228 35708 13234 35760
rect 23474 35748 23480 35760
rect 23435 35720 23480 35748
rect 23474 35708 23480 35720
rect 23532 35708 23538 35760
rect 24826 35695 24854 35788
rect 25133 35785 25145 35819
rect 25179 35816 25191 35819
rect 26234 35816 26240 35828
rect 25179 35788 26240 35816
rect 25179 35785 25191 35788
rect 25133 35779 25191 35785
rect 26234 35776 26240 35788
rect 26292 35776 26298 35828
rect 28258 35776 28264 35828
rect 28316 35816 28322 35828
rect 30650 35816 30656 35828
rect 28316 35788 30656 35816
rect 28316 35776 28322 35788
rect 30650 35776 30656 35788
rect 30708 35776 30714 35828
rect 33134 35776 33140 35828
rect 33192 35816 33198 35828
rect 33321 35819 33379 35825
rect 33321 35816 33333 35819
rect 33192 35788 33333 35816
rect 33192 35776 33198 35788
rect 33321 35785 33333 35788
rect 33367 35785 33379 35819
rect 33321 35779 33379 35785
rect 27982 35748 27988 35760
rect 7745 35683 7803 35689
rect 7576 35652 7696 35680
rect 7478 35643 7536 35649
rect 7668 35612 7696 35652
rect 7745 35649 7757 35683
rect 7791 35680 7803 35683
rect 10226 35680 10232 35692
rect 7791 35652 10232 35680
rect 7791 35649 7803 35652
rect 7745 35643 7803 35649
rect 10226 35640 10232 35652
rect 10284 35640 10290 35692
rect 11701 35683 11759 35689
rect 11701 35649 11713 35683
rect 11747 35680 11759 35683
rect 11974 35680 11980 35692
rect 11747 35652 11980 35680
rect 11747 35649 11759 35652
rect 11701 35643 11759 35649
rect 11974 35640 11980 35652
rect 12032 35640 12038 35692
rect 13357 35683 13415 35689
rect 13357 35649 13369 35683
rect 13403 35680 13415 35683
rect 13446 35680 13452 35692
rect 13403 35652 13452 35680
rect 13403 35649 13415 35652
rect 13357 35643 13415 35649
rect 13446 35640 13452 35652
rect 13504 35640 13510 35692
rect 16482 35640 16488 35692
rect 16540 35680 16546 35692
rect 17034 35680 17040 35692
rect 16540 35652 17040 35680
rect 16540 35640 16546 35652
rect 17034 35640 17040 35652
rect 17092 35680 17098 35692
rect 17405 35683 17463 35689
rect 17405 35680 17417 35683
rect 17092 35652 17417 35680
rect 17092 35640 17098 35652
rect 17405 35649 17417 35652
rect 17451 35649 17463 35683
rect 17405 35643 17463 35649
rect 17589 35683 17647 35689
rect 17589 35649 17601 35683
rect 17635 35680 17647 35683
rect 18506 35680 18512 35692
rect 17635 35652 18512 35680
rect 17635 35649 17647 35652
rect 17589 35643 17647 35649
rect 18506 35640 18512 35652
rect 18564 35640 18570 35692
rect 23658 35680 23664 35692
rect 23619 35652 23664 35680
rect 23658 35640 23664 35652
rect 23716 35640 23722 35692
rect 24394 35640 24400 35692
rect 24452 35680 24458 35692
rect 24784 35689 24854 35695
rect 27586 35720 27988 35748
rect 24489 35683 24547 35689
rect 24489 35680 24501 35683
rect 24452 35652 24501 35680
rect 24452 35640 24458 35652
rect 24489 35649 24501 35652
rect 24535 35649 24547 35683
rect 24489 35643 24547 35649
rect 24673 35683 24731 35689
rect 24673 35649 24685 35683
rect 24719 35649 24731 35683
rect 24784 35655 24796 35689
rect 24830 35658 24854 35689
rect 24903 35683 24961 35689
rect 24830 35655 24842 35658
rect 24784 35649 24842 35655
rect 24903 35649 24915 35683
rect 24949 35680 24961 35683
rect 25222 35680 25228 35692
rect 24949 35652 25228 35680
rect 24949 35649 24961 35652
rect 24673 35643 24731 35649
rect 24903 35643 24961 35649
rect 7926 35612 7932 35624
rect 7668 35584 7932 35612
rect 7926 35572 7932 35584
rect 7984 35612 7990 35624
rect 9033 35615 9091 35621
rect 9033 35612 9045 35615
rect 7984 35584 9045 35612
rect 7984 35572 7990 35584
rect 9033 35581 9045 35584
rect 9079 35581 9091 35615
rect 9306 35612 9312 35624
rect 9267 35584 9312 35612
rect 9033 35575 9091 35581
rect 9306 35572 9312 35584
rect 9364 35572 9370 35624
rect 9766 35612 9772 35624
rect 9727 35584 9772 35612
rect 9766 35572 9772 35584
rect 9824 35572 9830 35624
rect 10045 35615 10103 35621
rect 10045 35581 10057 35615
rect 10091 35612 10103 35615
rect 10134 35612 10140 35624
rect 10091 35584 10140 35612
rect 10091 35581 10103 35584
rect 10045 35575 10103 35581
rect 10134 35572 10140 35584
rect 10192 35612 10198 35624
rect 10686 35612 10692 35624
rect 10192 35584 10692 35612
rect 10192 35572 10198 35584
rect 10686 35572 10692 35584
rect 10744 35572 10750 35624
rect 23845 35615 23903 35621
rect 23845 35581 23857 35615
rect 23891 35612 23903 35615
rect 24688 35612 24716 35643
rect 25222 35640 25228 35652
rect 25280 35680 25286 35692
rect 25593 35683 25651 35689
rect 25593 35680 25605 35683
rect 25280 35652 25605 35680
rect 25280 35640 25286 35652
rect 25593 35649 25605 35652
rect 25639 35680 25651 35683
rect 27586 35680 27614 35720
rect 27982 35708 27988 35720
rect 28040 35708 28046 35760
rect 33505 35751 33563 35757
rect 33505 35717 33517 35751
rect 33551 35748 33563 35751
rect 33778 35748 33784 35760
rect 33551 35720 33784 35748
rect 33551 35717 33563 35720
rect 33505 35711 33563 35717
rect 33778 35708 33784 35720
rect 33836 35708 33842 35760
rect 25639 35652 27614 35680
rect 25639 35649 25651 35652
rect 25593 35643 25651 35649
rect 31754 35640 31760 35692
rect 31812 35680 31818 35692
rect 32217 35683 32275 35689
rect 32217 35680 32229 35683
rect 31812 35652 32229 35680
rect 31812 35640 31818 35652
rect 32217 35649 32229 35652
rect 32263 35649 32275 35683
rect 33686 35680 33692 35692
rect 33647 35652 33692 35680
rect 32217 35643 32275 35649
rect 33686 35640 33692 35652
rect 33744 35640 33750 35692
rect 23891 35584 24716 35612
rect 23891 35581 23903 35584
rect 23845 35575 23903 35581
rect 13998 35504 14004 35556
rect 14056 35544 14062 35556
rect 27157 35547 27215 35553
rect 27157 35544 27169 35547
rect 14056 35516 27169 35544
rect 14056 35504 14062 35516
rect 27157 35513 27169 35516
rect 27203 35544 27215 35547
rect 28166 35544 28172 35556
rect 27203 35516 28172 35544
rect 27203 35513 27215 35516
rect 27157 35507 27215 35513
rect 28166 35504 28172 35516
rect 28224 35504 28230 35556
rect 34149 35547 34207 35553
rect 34149 35544 34161 35547
rect 32324 35516 34161 35544
rect 4706 35476 4712 35488
rect 4667 35448 4712 35476
rect 4706 35436 4712 35448
rect 4764 35436 4770 35488
rect 5261 35479 5319 35485
rect 5261 35445 5273 35479
rect 5307 35476 5319 35479
rect 6086 35476 6092 35488
rect 5307 35448 6092 35476
rect 5307 35445 5319 35448
rect 5261 35439 5319 35445
rect 6086 35436 6092 35448
rect 6144 35436 6150 35488
rect 6365 35479 6423 35485
rect 6365 35445 6377 35479
rect 6411 35476 6423 35479
rect 6546 35476 6552 35488
rect 6411 35448 6552 35476
rect 6411 35445 6423 35448
rect 6365 35439 6423 35445
rect 6546 35436 6552 35448
rect 6604 35436 6610 35488
rect 10594 35436 10600 35488
rect 10652 35476 10658 35488
rect 11885 35479 11943 35485
rect 11885 35476 11897 35479
rect 10652 35448 11897 35476
rect 10652 35436 10658 35448
rect 11885 35445 11897 35448
rect 11931 35445 11943 35479
rect 13906 35476 13912 35488
rect 13867 35448 13912 35476
rect 11885 35439 11943 35445
rect 13906 35436 13912 35448
rect 13964 35476 13970 35488
rect 14734 35476 14740 35488
rect 13964 35448 14740 35476
rect 13964 35436 13970 35448
rect 14734 35436 14740 35448
rect 14792 35436 14798 35488
rect 17770 35476 17776 35488
rect 17731 35448 17776 35476
rect 17770 35436 17776 35448
rect 17828 35436 17834 35488
rect 22370 35476 22376 35488
rect 22331 35448 22376 35476
rect 22370 35436 22376 35448
rect 22428 35436 22434 35488
rect 23014 35476 23020 35488
rect 22975 35448 23020 35476
rect 23014 35436 23020 35448
rect 23072 35436 23078 35488
rect 25866 35436 25872 35488
rect 25924 35476 25930 35488
rect 32324 35476 32352 35516
rect 34149 35513 34161 35516
rect 34195 35544 34207 35547
rect 34238 35544 34244 35556
rect 34195 35516 34244 35544
rect 34195 35513 34207 35516
rect 34149 35507 34207 35513
rect 34238 35504 34244 35516
rect 34296 35544 34302 35556
rect 36446 35544 36452 35556
rect 34296 35516 36452 35544
rect 34296 35504 34302 35516
rect 36446 35504 36452 35516
rect 36504 35504 36510 35556
rect 25924 35448 32352 35476
rect 32401 35479 32459 35485
rect 25924 35436 25930 35448
rect 32401 35445 32413 35479
rect 32447 35476 32459 35479
rect 33686 35476 33692 35488
rect 32447 35448 33692 35476
rect 32447 35445 32459 35448
rect 32401 35439 32459 35445
rect 33686 35436 33692 35448
rect 33744 35436 33750 35488
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 4249 35275 4307 35281
rect 4249 35241 4261 35275
rect 4295 35272 4307 35275
rect 4614 35272 4620 35284
rect 4295 35244 4620 35272
rect 4295 35241 4307 35244
rect 4249 35235 4307 35241
rect 4614 35232 4620 35244
rect 4672 35232 4678 35284
rect 6086 35272 6092 35284
rect 4724 35244 6092 35272
rect 4724 35136 4752 35244
rect 6086 35232 6092 35244
rect 6144 35232 6150 35284
rect 7190 35272 7196 35284
rect 7151 35244 7196 35272
rect 7190 35232 7196 35244
rect 7248 35232 7254 35284
rect 8389 35275 8447 35281
rect 7392 35244 7696 35272
rect 4982 35204 4988 35216
rect 4540 35108 4752 35136
rect 4908 35176 4988 35204
rect 4540 35077 4568 35108
rect 4525 35071 4583 35077
rect 4525 35037 4537 35071
rect 4571 35037 4583 35071
rect 4525 35031 4583 35037
rect 4617 35071 4675 35077
rect 4617 35037 4629 35071
rect 4663 35037 4675 35071
rect 4617 35031 4675 35037
rect 2682 34960 2688 35012
rect 2740 35000 2746 35012
rect 4632 35000 4660 35031
rect 4706 35028 4712 35080
rect 4764 35068 4770 35080
rect 4908 35077 4936 35176
rect 4982 35164 4988 35176
rect 5040 35164 5046 35216
rect 6733 35207 6791 35213
rect 6733 35173 6745 35207
rect 6779 35204 6791 35207
rect 7392 35204 7420 35244
rect 7558 35204 7564 35216
rect 6779 35176 7420 35204
rect 7464 35176 7564 35204
rect 6779 35173 6791 35176
rect 6733 35167 6791 35173
rect 7464 35077 7492 35176
rect 7558 35164 7564 35176
rect 7616 35164 7622 35216
rect 7668 35077 7696 35244
rect 8389 35241 8401 35275
rect 8435 35272 8447 35275
rect 11974 35272 11980 35284
rect 8435 35244 11560 35272
rect 11935 35244 11980 35272
rect 8435 35241 8447 35244
rect 8389 35235 8447 35241
rect 4893 35071 4951 35077
rect 4764 35040 4809 35068
rect 4764 35028 4770 35040
rect 4893 35037 4905 35071
rect 4939 35037 4951 35071
rect 4893 35031 4951 35037
rect 7449 35071 7507 35077
rect 7449 35037 7461 35071
rect 7495 35037 7507 35071
rect 7449 35031 7507 35037
rect 7561 35071 7619 35077
rect 7561 35037 7573 35071
rect 7607 35037 7619 35071
rect 7561 35031 7619 35037
rect 7653 35071 7711 35077
rect 7653 35037 7665 35071
rect 7699 35037 7711 35071
rect 7653 35031 7711 35037
rect 7837 35071 7895 35077
rect 7837 35037 7849 35071
rect 7883 35068 7895 35071
rect 8404 35068 8432 35235
rect 11532 35204 11560 35244
rect 11974 35232 11980 35244
rect 12032 35232 12038 35284
rect 19150 35272 19156 35284
rect 12406 35244 19156 35272
rect 12406 35204 12434 35244
rect 19150 35232 19156 35244
rect 19208 35272 19214 35284
rect 19426 35272 19432 35284
rect 19208 35244 19432 35272
rect 19208 35232 19214 35244
rect 19426 35232 19432 35244
rect 19484 35232 19490 35284
rect 25038 35272 25044 35284
rect 24999 35244 25044 35272
rect 25038 35232 25044 35244
rect 25096 35232 25102 35284
rect 25958 35204 25964 35216
rect 11532 35176 12434 35204
rect 25516 35176 25964 35204
rect 9861 35139 9919 35145
rect 9861 35105 9873 35139
rect 9907 35136 9919 35139
rect 10042 35136 10048 35148
rect 9907 35108 10048 35136
rect 9907 35105 9919 35108
rect 9861 35099 9919 35105
rect 10042 35096 10048 35108
rect 10100 35096 10106 35148
rect 10226 35096 10232 35148
rect 10284 35136 10290 35148
rect 10597 35139 10655 35145
rect 10597 35136 10609 35139
rect 10284 35108 10609 35136
rect 10284 35096 10290 35108
rect 10597 35105 10609 35108
rect 10643 35105 10655 35139
rect 10597 35099 10655 35105
rect 15378 35096 15384 35148
rect 15436 35136 15442 35148
rect 17129 35139 17187 35145
rect 17129 35136 17141 35139
rect 15436 35108 17141 35136
rect 15436 35096 15442 35108
rect 17129 35105 17141 35108
rect 17175 35105 17187 35139
rect 17129 35099 17187 35105
rect 18598 35096 18604 35148
rect 18656 35136 18662 35148
rect 21637 35139 21695 35145
rect 18656 35108 20668 35136
rect 18656 35096 18662 35108
rect 7883 35040 8432 35068
rect 7883 35037 7895 35040
rect 7837 35031 7895 35037
rect 5350 35000 5356 35012
rect 2740 34972 5356 35000
rect 2740 34960 2746 34972
rect 5350 34960 5356 34972
rect 5408 34960 5414 35012
rect 6362 35000 6368 35012
rect 6323 34972 6368 35000
rect 6362 34960 6368 34972
rect 6420 34960 6426 35012
rect 6546 35000 6552 35012
rect 6507 34972 6552 35000
rect 6546 34960 6552 34972
rect 6604 34960 6610 35012
rect 6730 34960 6736 35012
rect 6788 35000 6794 35012
rect 7576 35000 7604 35031
rect 9950 35028 9956 35080
rect 10008 35068 10014 35080
rect 10137 35071 10195 35077
rect 10137 35068 10149 35071
rect 10008 35040 10149 35068
rect 10008 35028 10014 35040
rect 10137 35037 10149 35040
rect 10183 35037 10195 35071
rect 10137 35031 10195 35037
rect 11974 35028 11980 35080
rect 12032 35068 12038 35080
rect 13009 35071 13067 35077
rect 13009 35068 13021 35071
rect 12032 35040 13021 35068
rect 12032 35028 12038 35040
rect 13009 35037 13021 35040
rect 13055 35037 13067 35071
rect 13009 35031 13067 35037
rect 13357 35071 13415 35077
rect 13357 35037 13369 35071
rect 13403 35068 13415 35071
rect 13446 35068 13452 35080
rect 13403 35040 13452 35068
rect 13403 35037 13415 35040
rect 13357 35031 13415 35037
rect 13446 35028 13452 35040
rect 13504 35028 13510 35080
rect 17678 35028 17684 35080
rect 17736 35068 17742 35080
rect 20530 35068 20536 35080
rect 17736 35040 20536 35068
rect 17736 35028 17742 35040
rect 20530 35028 20536 35040
rect 20588 35028 20594 35080
rect 20640 35068 20668 35108
rect 21637 35105 21649 35139
rect 21683 35136 21695 35139
rect 22002 35136 22008 35148
rect 21683 35108 22008 35136
rect 21683 35105 21695 35108
rect 21637 35099 21695 35105
rect 22002 35096 22008 35108
rect 22060 35096 22066 35148
rect 23842 35096 23848 35148
rect 23900 35136 23906 35148
rect 23900 35108 24532 35136
rect 23900 35096 23906 35108
rect 22097 35071 22155 35077
rect 22097 35068 22109 35071
rect 20640 35040 22109 35068
rect 22097 35037 22109 35040
rect 22143 35068 22155 35071
rect 22738 35068 22744 35080
rect 22143 35040 22744 35068
rect 22143 35037 22155 35040
rect 22097 35031 22155 35037
rect 22738 35028 22744 35040
rect 22796 35028 22802 35080
rect 24394 35068 24400 35080
rect 23952 35040 24400 35068
rect 6788 34972 7604 35000
rect 10864 35003 10922 35009
rect 6788 34960 6794 34972
rect 10864 34969 10876 35003
rect 10910 35000 10922 35003
rect 11054 35000 11060 35012
rect 10910 34972 11060 35000
rect 10910 34969 10922 34972
rect 10864 34963 10922 34969
rect 11054 34960 11060 34972
rect 11112 34960 11118 35012
rect 13170 35000 13176 35012
rect 13131 34972 13176 35000
rect 13170 34960 13176 34972
rect 13228 34960 13234 35012
rect 13265 35003 13323 35009
rect 13265 34969 13277 35003
rect 13311 35000 13323 35003
rect 14090 35000 14096 35012
rect 13311 34972 14096 35000
rect 13311 34969 13323 34972
rect 13265 34963 13323 34969
rect 14090 34960 14096 34972
rect 14148 34960 14154 35012
rect 17126 34960 17132 35012
rect 17184 35000 17190 35012
rect 17374 35003 17432 35009
rect 17374 35000 17386 35003
rect 17184 34972 17386 35000
rect 17184 34960 17190 34972
rect 17374 34969 17386 34972
rect 17420 34969 17432 35003
rect 17374 34963 17432 34969
rect 20346 34960 20352 35012
rect 20404 35000 20410 35012
rect 21370 35003 21428 35009
rect 21370 35000 21382 35003
rect 20404 34972 21382 35000
rect 20404 34960 20410 34972
rect 21370 34969 21382 34972
rect 21416 34969 21428 35003
rect 21370 34963 21428 34969
rect 23952 34944 23980 35040
rect 24394 35028 24400 35040
rect 24452 35028 24458 35080
rect 24504 35068 24532 35108
rect 24581 35071 24639 35077
rect 24581 35068 24593 35071
rect 24504 35040 24593 35068
rect 24581 35037 24593 35040
rect 24627 35037 24639 35071
rect 24581 35031 24639 35037
rect 24670 35028 24676 35080
rect 24728 35068 24734 35080
rect 24811 35071 24869 35077
rect 24728 35040 24773 35068
rect 24728 35028 24734 35040
rect 24811 35037 24823 35071
rect 24857 35037 24869 35071
rect 24811 35031 24869 35037
rect 5445 34935 5503 34941
rect 5445 34901 5457 34935
rect 5491 34932 5503 34935
rect 5626 34932 5632 34944
rect 5491 34904 5632 34932
rect 5491 34901 5503 34904
rect 5445 34895 5503 34901
rect 5626 34892 5632 34904
rect 5684 34892 5690 34944
rect 13541 34935 13599 34941
rect 13541 34901 13553 34935
rect 13587 34932 13599 34935
rect 15102 34932 15108 34944
rect 13587 34904 15108 34932
rect 13587 34901 13599 34904
rect 13541 34895 13599 34901
rect 15102 34892 15108 34904
rect 15160 34892 15166 34944
rect 18506 34932 18512 34944
rect 18467 34904 18512 34932
rect 18506 34892 18512 34904
rect 18564 34892 18570 34944
rect 20254 34932 20260 34944
rect 20215 34904 20260 34932
rect 20254 34892 20260 34904
rect 20312 34892 20318 34944
rect 22186 34892 22192 34944
rect 22244 34932 22250 34944
rect 22554 34932 22560 34944
rect 22244 34904 22560 34932
rect 22244 34892 22250 34904
rect 22554 34892 22560 34904
rect 22612 34892 22618 34944
rect 23845 34935 23903 34941
rect 23845 34901 23857 34935
rect 23891 34932 23903 34935
rect 23934 34932 23940 34944
rect 23891 34904 23940 34932
rect 23891 34901 23903 34904
rect 23845 34895 23903 34901
rect 23934 34892 23940 34904
rect 23992 34892 23998 34944
rect 24302 34892 24308 34944
rect 24360 34932 24366 34944
rect 24841 34932 24869 35031
rect 25516 34941 25544 35176
rect 25958 35164 25964 35176
rect 26016 35204 26022 35216
rect 33318 35204 33324 35216
rect 26016 35176 33324 35204
rect 26016 35164 26022 35176
rect 33318 35164 33324 35176
rect 33376 35164 33382 35216
rect 29270 35028 29276 35080
rect 29328 35068 29334 35080
rect 30190 35068 30196 35080
rect 29328 35040 30196 35068
rect 29328 35028 29334 35040
rect 30190 35028 30196 35040
rect 30248 35068 30254 35080
rect 31481 35071 31539 35077
rect 31481 35068 31493 35071
rect 30248 35040 31493 35068
rect 30248 35028 30254 35040
rect 31481 35037 31493 35040
rect 31527 35037 31539 35071
rect 31481 35031 31539 35037
rect 31754 35028 31760 35080
rect 31812 35068 31818 35080
rect 58158 35068 58164 35080
rect 31812 35040 31857 35068
rect 58119 35040 58164 35068
rect 31812 35028 31818 35040
rect 58158 35028 58164 35040
rect 58216 35028 58222 35080
rect 28902 34960 28908 35012
rect 28960 35000 28966 35012
rect 29822 35000 29828 35012
rect 28960 34972 29828 35000
rect 28960 34960 28966 34972
rect 29822 34960 29828 34972
rect 29880 34960 29886 35012
rect 30285 35003 30343 35009
rect 30285 34969 30297 35003
rect 30331 34969 30343 35003
rect 30285 34963 30343 34969
rect 25501 34935 25559 34941
rect 25501 34932 25513 34935
rect 24360 34904 25513 34932
rect 24360 34892 24366 34904
rect 25501 34901 25513 34904
rect 25547 34901 25559 34935
rect 25501 34895 25559 34901
rect 29546 34892 29552 34944
rect 29604 34932 29610 34944
rect 30101 34935 30159 34941
rect 30101 34932 30113 34935
rect 29604 34904 30113 34932
rect 29604 34892 29610 34904
rect 30101 34901 30113 34904
rect 30147 34901 30159 34935
rect 30300 34932 30328 34963
rect 30466 34960 30472 35012
rect 30524 35000 30530 35012
rect 31202 35000 31208 35012
rect 30524 34972 31208 35000
rect 30524 34960 30530 34972
rect 31202 34960 31208 34972
rect 31260 34960 31266 35012
rect 31570 34932 31576 34944
rect 30300 34904 31576 34932
rect 30101 34895 30159 34901
rect 31570 34892 31576 34904
rect 31628 34892 31634 34944
rect 33689 34935 33747 34941
rect 33689 34901 33701 34935
rect 33735 34932 33747 34935
rect 34238 34932 34244 34944
rect 33735 34904 34244 34932
rect 33735 34901 33747 34904
rect 33689 34895 33747 34901
rect 34238 34892 34244 34904
rect 34296 34892 34302 34944
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 3973 34731 4031 34737
rect 3973 34697 3985 34731
rect 4019 34728 4031 34731
rect 4614 34728 4620 34740
rect 4019 34700 4620 34728
rect 4019 34697 4031 34700
rect 3973 34691 4031 34697
rect 4614 34688 4620 34700
rect 4672 34688 4678 34740
rect 5626 34728 5632 34740
rect 4724 34700 5632 34728
rect 2860 34663 2918 34669
rect 2860 34629 2872 34663
rect 2906 34660 2918 34663
rect 4433 34663 4491 34669
rect 4433 34660 4445 34663
rect 2906 34632 4445 34660
rect 2906 34629 2918 34632
rect 2860 34623 2918 34629
rect 4433 34629 4445 34632
rect 4479 34629 4491 34663
rect 4724 34660 4752 34700
rect 5626 34688 5632 34700
rect 5684 34688 5690 34740
rect 9033 34731 9091 34737
rect 9033 34697 9045 34731
rect 9079 34728 9091 34731
rect 9122 34728 9128 34740
rect 9079 34700 9128 34728
rect 9079 34697 9091 34700
rect 9033 34691 9091 34697
rect 9122 34688 9128 34700
rect 9180 34688 9186 34740
rect 10321 34731 10379 34737
rect 10321 34697 10333 34731
rect 10367 34728 10379 34731
rect 10410 34728 10416 34740
rect 10367 34700 10416 34728
rect 10367 34697 10379 34700
rect 10321 34691 10379 34697
rect 10410 34688 10416 34700
rect 10468 34688 10474 34740
rect 12437 34731 12495 34737
rect 12437 34728 12449 34731
rect 10591 34700 12449 34728
rect 4433 34623 4491 34629
rect 4540 34632 4752 34660
rect 4908 34632 5028 34660
rect 2590 34592 2596 34604
rect 2551 34564 2596 34592
rect 2590 34552 2596 34564
rect 2648 34552 2654 34604
rect 4540 34592 4568 34632
rect 4908 34601 4936 34632
rect 4709 34595 4767 34601
rect 4632 34592 4721 34595
rect 4540 34567 4721 34592
rect 4540 34564 4660 34567
rect 4709 34561 4721 34567
rect 4755 34561 4767 34595
rect 4709 34555 4767 34561
rect 4798 34595 4856 34601
rect 4798 34561 4810 34595
rect 4844 34561 4856 34595
rect 4798 34555 4856 34561
rect 4893 34595 4951 34601
rect 4893 34561 4905 34595
rect 4939 34561 4951 34595
rect 4893 34555 4951 34561
rect 4813 34524 4841 34555
rect 4632 34496 4841 34524
rect 4632 34388 4660 34496
rect 4706 34416 4712 34468
rect 4764 34456 4770 34468
rect 5000 34456 5028 34632
rect 6546 34620 6552 34672
rect 6604 34660 6610 34672
rect 8757 34663 8815 34669
rect 8757 34660 8769 34663
rect 6604 34632 8769 34660
rect 6604 34620 6610 34632
rect 8757 34629 8769 34632
rect 8803 34629 8815 34663
rect 9490 34660 9496 34672
rect 9451 34632 9496 34660
rect 8757 34623 8815 34629
rect 9490 34620 9496 34632
rect 9548 34620 9554 34672
rect 5077 34595 5135 34601
rect 5077 34561 5089 34595
rect 5123 34592 5135 34595
rect 5442 34592 5448 34604
rect 5123 34564 5448 34592
rect 5123 34561 5135 34564
rect 5077 34555 5135 34561
rect 5442 34552 5448 34564
rect 5500 34552 5506 34604
rect 7558 34552 7564 34604
rect 7616 34592 7622 34604
rect 7837 34595 7895 34601
rect 7837 34592 7849 34595
rect 7616 34564 7849 34592
rect 7616 34552 7622 34564
rect 7837 34561 7849 34564
rect 7883 34561 7895 34595
rect 8386 34592 8392 34604
rect 8347 34564 8392 34592
rect 7837 34555 7895 34561
rect 8386 34552 8392 34564
rect 8444 34552 8450 34604
rect 8482 34595 8540 34601
rect 8482 34561 8494 34595
rect 8528 34561 8540 34595
rect 8662 34592 8668 34604
rect 8623 34564 8668 34592
rect 8482 34555 8540 34561
rect 8018 34484 8024 34536
rect 8076 34524 8082 34536
rect 8496 34524 8524 34555
rect 8662 34552 8668 34564
rect 8720 34552 8726 34604
rect 8895 34595 8953 34601
rect 8895 34561 8907 34595
rect 8941 34592 8953 34595
rect 9582 34592 9588 34604
rect 8941 34564 9588 34592
rect 8941 34561 8953 34564
rect 8895 34555 8953 34561
rect 9582 34552 9588 34564
rect 9640 34552 9646 34604
rect 9677 34595 9735 34601
rect 9677 34561 9689 34595
rect 9723 34592 9735 34595
rect 9950 34592 9956 34604
rect 9723 34564 9956 34592
rect 9723 34561 9735 34564
rect 9677 34555 9735 34561
rect 9950 34552 9956 34564
rect 10008 34552 10014 34604
rect 10591 34601 10619 34700
rect 12437 34697 12449 34700
rect 12483 34728 12495 34731
rect 13633 34731 13691 34737
rect 12483 34700 13492 34728
rect 12483 34697 12495 34700
rect 12437 34691 12495 34697
rect 11885 34663 11943 34669
rect 11885 34660 11897 34663
rect 10796 34632 11897 34660
rect 10796 34601 10824 34632
rect 11885 34629 11897 34632
rect 11931 34629 11943 34663
rect 11885 34623 11943 34629
rect 12802 34620 12808 34672
rect 12860 34660 12866 34672
rect 13357 34663 13415 34669
rect 13357 34660 13369 34663
rect 12860 34632 13369 34660
rect 12860 34620 12866 34632
rect 13357 34629 13369 34632
rect 13403 34629 13415 34663
rect 13464 34660 13492 34700
rect 13633 34697 13645 34731
rect 13679 34728 13691 34731
rect 16114 34728 16120 34740
rect 13679 34700 16120 34728
rect 13679 34697 13691 34700
rect 13633 34691 13691 34697
rect 16114 34688 16120 34700
rect 16172 34688 16178 34740
rect 17126 34728 17132 34740
rect 17087 34700 17132 34728
rect 17126 34688 17132 34700
rect 17184 34688 17190 34740
rect 17586 34688 17592 34740
rect 17644 34728 17650 34740
rect 20070 34728 20076 34740
rect 17644 34700 17816 34728
rect 17644 34688 17650 34700
rect 16298 34660 16304 34672
rect 13464 34632 16304 34660
rect 13357 34623 13415 34629
rect 16298 34620 16304 34632
rect 16356 34620 16362 34672
rect 17310 34620 17316 34672
rect 17368 34660 17374 34672
rect 17368 34632 17540 34660
rect 17368 34620 17374 34632
rect 10577 34595 10635 34601
rect 10577 34561 10589 34595
rect 10623 34561 10635 34595
rect 10577 34555 10635 34561
rect 10670 34595 10728 34601
rect 10670 34561 10682 34595
rect 10716 34561 10728 34595
rect 10670 34555 10728 34561
rect 10781 34595 10839 34601
rect 10781 34561 10793 34595
rect 10827 34561 10839 34595
rect 10962 34592 10968 34604
rect 10923 34564 10968 34592
rect 10781 34555 10839 34561
rect 8076 34496 8524 34524
rect 8076 34484 8082 34496
rect 10042 34484 10048 34536
rect 10100 34524 10106 34536
rect 10685 34524 10713 34555
rect 10962 34552 10968 34564
rect 11020 34552 11026 34604
rect 11514 34592 11520 34604
rect 11475 34564 11520 34592
rect 11514 34552 11520 34564
rect 11572 34552 11578 34604
rect 11698 34592 11704 34604
rect 11659 34564 11704 34592
rect 11698 34552 11704 34564
rect 11756 34592 11762 34604
rect 13081 34595 13139 34601
rect 13081 34592 13093 34595
rect 11756 34564 13093 34592
rect 11756 34552 11762 34564
rect 13081 34561 13093 34564
rect 13127 34561 13139 34595
rect 13262 34592 13268 34604
rect 13223 34564 13268 34592
rect 13081 34555 13139 34561
rect 13262 34552 13268 34564
rect 13320 34552 13326 34604
rect 13446 34552 13452 34604
rect 13504 34592 13510 34604
rect 16758 34592 16764 34604
rect 13504 34564 13597 34592
rect 16040 34564 16764 34592
rect 13504 34552 13510 34564
rect 10100 34496 10713 34524
rect 10100 34484 10106 34496
rect 13170 34484 13176 34536
rect 13228 34524 13234 34536
rect 13464 34524 13492 34552
rect 13228 34496 13492 34524
rect 13228 34484 13234 34496
rect 4764 34428 5028 34456
rect 4764 34416 4770 34428
rect 11514 34416 11520 34468
rect 11572 34456 11578 34468
rect 16040 34465 16068 34564
rect 16758 34552 16764 34564
rect 16816 34592 16822 34604
rect 17512 34601 17540 34632
rect 17405 34595 17463 34601
rect 17405 34592 17417 34595
rect 16816 34564 17417 34592
rect 16816 34552 16822 34564
rect 17405 34561 17417 34564
rect 17451 34561 17463 34595
rect 17405 34555 17463 34561
rect 17497 34595 17555 34601
rect 17497 34561 17509 34595
rect 17543 34561 17555 34595
rect 17497 34555 17555 34561
rect 17589 34595 17647 34601
rect 17589 34561 17601 34595
rect 17635 34592 17647 34595
rect 17678 34592 17684 34604
rect 17635 34564 17684 34592
rect 17635 34561 17647 34564
rect 17589 34555 17647 34561
rect 17678 34552 17684 34564
rect 17736 34552 17742 34604
rect 17788 34601 17816 34700
rect 18800 34700 20076 34728
rect 17773 34595 17831 34601
rect 17773 34561 17785 34595
rect 17819 34592 17831 34595
rect 17862 34592 17868 34604
rect 17819 34564 17868 34592
rect 17819 34561 17831 34564
rect 17773 34555 17831 34561
rect 17862 34552 17868 34564
rect 17920 34552 17926 34604
rect 18690 34552 18696 34604
rect 18748 34592 18754 34604
rect 18800 34601 18828 34700
rect 20070 34688 20076 34700
rect 20128 34688 20134 34740
rect 20257 34731 20315 34737
rect 20257 34697 20269 34731
rect 20303 34728 20315 34731
rect 20346 34728 20352 34740
rect 20303 34700 20352 34728
rect 20303 34697 20315 34700
rect 20257 34691 20315 34697
rect 20346 34688 20352 34700
rect 20404 34688 20410 34740
rect 20809 34731 20867 34737
rect 20809 34697 20821 34731
rect 20855 34728 20867 34731
rect 25866 34728 25872 34740
rect 20855 34700 25872 34728
rect 20855 34697 20867 34700
rect 20809 34691 20867 34697
rect 18969 34663 19027 34669
rect 18969 34629 18981 34663
rect 19015 34660 19027 34663
rect 20530 34660 20536 34672
rect 19015 34632 20300 34660
rect 20443 34632 20536 34660
rect 19015 34629 19027 34632
rect 18969 34623 19027 34629
rect 20272 34604 20300 34632
rect 20530 34620 20536 34632
rect 20588 34660 20594 34672
rect 20824 34660 20852 34691
rect 25866 34688 25872 34700
rect 25924 34688 25930 34740
rect 30558 34728 30564 34740
rect 29012 34700 30564 34728
rect 20588 34632 20852 34660
rect 20588 34620 20594 34632
rect 21818 34620 21824 34672
rect 21876 34660 21882 34672
rect 27893 34663 27951 34669
rect 21876 34632 22324 34660
rect 21876 34620 21882 34632
rect 18785 34595 18843 34601
rect 18785 34592 18797 34595
rect 18748 34564 18797 34592
rect 18748 34552 18754 34564
rect 18785 34561 18797 34564
rect 18831 34561 18843 34595
rect 18785 34555 18843 34561
rect 19426 34552 19432 34604
rect 19484 34592 19490 34604
rect 19613 34595 19671 34601
rect 19613 34592 19625 34595
rect 19484 34564 19625 34592
rect 19484 34552 19490 34564
rect 19613 34561 19625 34564
rect 19659 34561 19671 34595
rect 19613 34555 19671 34561
rect 19797 34595 19855 34601
rect 19797 34561 19809 34595
rect 19843 34561 19855 34595
rect 19797 34555 19855 34561
rect 19889 34595 19947 34601
rect 19889 34561 19901 34595
rect 19935 34561 19947 34595
rect 19889 34555 19947 34561
rect 19981 34595 20039 34601
rect 19981 34561 19993 34595
rect 20027 34561 20039 34595
rect 19981 34555 20039 34561
rect 18046 34484 18052 34536
rect 18104 34524 18110 34536
rect 19153 34527 19211 34533
rect 18104 34496 19104 34524
rect 18104 34484 18110 34496
rect 16025 34459 16083 34465
rect 16025 34456 16037 34459
rect 11572 34428 16037 34456
rect 11572 34416 11578 34428
rect 16025 34425 16037 34428
rect 16071 34425 16083 34459
rect 16025 34419 16083 34425
rect 16298 34416 16304 34468
rect 16356 34456 16362 34468
rect 17494 34456 17500 34468
rect 16356 34428 17500 34456
rect 16356 34416 16362 34428
rect 17494 34416 17500 34428
rect 17552 34456 17558 34468
rect 18598 34456 18604 34468
rect 17552 34428 18604 34456
rect 17552 34416 17558 34428
rect 18598 34416 18604 34428
rect 18656 34416 18662 34468
rect 19076 34456 19104 34496
rect 19153 34493 19165 34527
rect 19199 34524 19211 34527
rect 19812 34524 19840 34555
rect 19199 34496 19840 34524
rect 19199 34493 19211 34496
rect 19153 34487 19211 34493
rect 19242 34456 19248 34468
rect 19076 34428 19248 34456
rect 19242 34416 19248 34428
rect 19300 34456 19306 34468
rect 19904 34456 19932 34555
rect 19996 34524 20024 34555
rect 20254 34552 20260 34604
rect 20312 34552 20318 34604
rect 20548 34524 20576 34620
rect 20622 34552 20628 34604
rect 20680 34592 20686 34604
rect 21726 34592 21732 34604
rect 20680 34564 21732 34592
rect 20680 34552 20686 34564
rect 21726 34552 21732 34564
rect 21784 34552 21790 34604
rect 22186 34592 22192 34604
rect 22147 34564 22192 34592
rect 22186 34552 22192 34564
rect 22244 34552 22250 34604
rect 22296 34592 22324 34632
rect 27893 34629 27905 34663
rect 27939 34660 27951 34663
rect 28350 34660 28356 34672
rect 27939 34632 28356 34660
rect 27939 34629 27951 34632
rect 27893 34623 27951 34629
rect 28350 34620 28356 34632
rect 28408 34620 28414 34672
rect 29012 34660 29040 34700
rect 30558 34688 30564 34700
rect 30616 34688 30622 34740
rect 31570 34728 31576 34740
rect 31531 34700 31576 34728
rect 31570 34688 31576 34700
rect 31628 34688 31634 34740
rect 33962 34688 33968 34740
rect 34020 34688 34026 34740
rect 28828 34632 29040 34660
rect 29089 34663 29147 34669
rect 22352 34595 22410 34601
rect 22468 34598 22526 34604
rect 22468 34595 22480 34598
rect 22352 34592 22364 34595
rect 22296 34564 22364 34592
rect 22352 34561 22364 34564
rect 22398 34561 22410 34595
rect 22352 34555 22410 34561
rect 22467 34564 22480 34595
rect 22514 34564 22526 34598
rect 22467 34558 22526 34564
rect 22557 34595 22615 34601
rect 22557 34561 22569 34595
rect 22603 34592 22692 34595
rect 22738 34592 22744 34604
rect 22603 34567 22744 34592
rect 22603 34561 22615 34567
rect 22664 34564 22744 34567
rect 19996 34496 20576 34524
rect 21542 34484 21548 34536
rect 21600 34524 21606 34536
rect 22094 34524 22100 34536
rect 21600 34496 22100 34524
rect 21600 34484 21606 34496
rect 22094 34484 22100 34496
rect 22152 34484 22158 34536
rect 22467 34468 22495 34558
rect 22557 34555 22615 34561
rect 22738 34552 22744 34564
rect 22796 34552 22802 34604
rect 28077 34595 28135 34601
rect 28077 34561 28089 34595
rect 28123 34592 28135 34595
rect 28828 34592 28856 34632
rect 29089 34629 29101 34663
rect 29135 34660 29147 34663
rect 30438 34663 30496 34669
rect 30438 34660 30450 34663
rect 29135 34632 30450 34660
rect 29135 34629 29147 34632
rect 29089 34623 29147 34629
rect 30438 34629 30450 34632
rect 30484 34629 30496 34663
rect 33980 34660 34008 34688
rect 33980 34632 34100 34660
rect 30438 34623 30496 34629
rect 34072 34604 34100 34632
rect 29365 34595 29423 34601
rect 29365 34592 29377 34595
rect 28123 34564 28856 34592
rect 28920 34564 29377 34592
rect 28123 34561 28135 34564
rect 28077 34555 28135 34561
rect 28258 34484 28264 34536
rect 28316 34524 28322 34536
rect 28537 34527 28595 34533
rect 28537 34524 28549 34527
rect 28316 34496 28549 34524
rect 28316 34484 28322 34496
rect 28537 34493 28549 34496
rect 28583 34524 28595 34527
rect 28920 34524 28948 34564
rect 29365 34561 29377 34564
rect 29411 34561 29423 34595
rect 29365 34555 29423 34561
rect 29457 34595 29515 34601
rect 29457 34561 29469 34595
rect 29503 34561 29515 34595
rect 29457 34555 29515 34561
rect 28583 34496 28948 34524
rect 28583 34493 28595 34496
rect 28537 34487 28595 34493
rect 19300 34428 19932 34456
rect 19300 34416 19306 34428
rect 22462 34416 22468 34468
rect 22520 34416 22526 34468
rect 28994 34416 29000 34468
rect 29052 34456 29058 34468
rect 29472 34456 29500 34555
rect 29546 34552 29552 34604
rect 29604 34592 29610 34604
rect 29604 34564 29649 34592
rect 29604 34552 29610 34564
rect 29730 34552 29736 34604
rect 29788 34592 29794 34604
rect 29788 34564 29833 34592
rect 29788 34552 29794 34564
rect 33502 34552 33508 34604
rect 33560 34592 33566 34604
rect 33781 34595 33839 34601
rect 33781 34592 33793 34595
rect 33560 34564 33793 34592
rect 33560 34552 33566 34564
rect 33781 34561 33793 34564
rect 33827 34561 33839 34595
rect 33781 34555 33839 34561
rect 33965 34595 34023 34601
rect 33965 34561 33977 34595
rect 34011 34561 34023 34595
rect 33965 34555 34023 34561
rect 34060 34598 34118 34604
rect 34060 34564 34072 34598
rect 34106 34564 34118 34598
rect 34060 34558 34118 34564
rect 34149 34595 34207 34601
rect 34149 34561 34161 34595
rect 34195 34592 34207 34595
rect 34238 34592 34244 34604
rect 34195 34564 34244 34592
rect 34195 34561 34207 34564
rect 34149 34555 34207 34561
rect 29822 34484 29828 34536
rect 29880 34524 29886 34536
rect 30193 34527 30251 34533
rect 30193 34524 30205 34527
rect 29880 34496 30205 34524
rect 29880 34484 29886 34496
rect 30193 34493 30205 34496
rect 30239 34493 30251 34527
rect 33980 34524 34008 34555
rect 34238 34552 34244 34564
rect 34296 34552 34302 34604
rect 34425 34527 34483 34533
rect 33980 34496 34376 34524
rect 30193 34487 30251 34493
rect 34348 34456 34376 34496
rect 34425 34493 34437 34527
rect 34471 34524 34483 34527
rect 35802 34524 35808 34536
rect 34471 34496 35808 34524
rect 34471 34493 34483 34496
rect 34425 34487 34483 34493
rect 35802 34484 35808 34496
rect 35860 34484 35866 34536
rect 34790 34456 34796 34468
rect 29052 34428 30236 34456
rect 34348 34428 34796 34456
rect 29052 34416 29058 34428
rect 30208 34400 30236 34428
rect 34790 34416 34796 34428
rect 34848 34416 34854 34468
rect 4890 34388 4896 34400
rect 4632 34360 4896 34388
rect 4890 34348 4896 34360
rect 4948 34348 4954 34400
rect 5442 34348 5448 34400
rect 5500 34388 5506 34400
rect 5537 34391 5595 34397
rect 5537 34388 5549 34391
rect 5500 34360 5549 34388
rect 5500 34348 5506 34360
rect 5537 34357 5549 34360
rect 5583 34357 5595 34391
rect 5537 34351 5595 34357
rect 7558 34348 7564 34400
rect 7616 34388 7622 34400
rect 11790 34388 11796 34400
rect 7616 34360 11796 34388
rect 7616 34348 7622 34360
rect 11790 34348 11796 34360
rect 11848 34348 11854 34400
rect 14550 34348 14556 34400
rect 14608 34388 14614 34400
rect 19794 34388 19800 34400
rect 14608 34360 19800 34388
rect 14608 34348 14614 34360
rect 19794 34348 19800 34360
rect 19852 34348 19858 34400
rect 22830 34388 22836 34400
rect 22791 34360 22836 34388
rect 22830 34348 22836 34360
rect 22888 34348 22894 34400
rect 24762 34388 24768 34400
rect 24723 34360 24768 34388
rect 24762 34348 24768 34360
rect 24820 34348 24826 34400
rect 27706 34388 27712 34400
rect 27667 34360 27712 34388
rect 27706 34348 27712 34360
rect 27764 34348 27770 34400
rect 30190 34348 30196 34400
rect 30248 34348 30254 34400
rect 33318 34388 33324 34400
rect 33231 34360 33324 34388
rect 33318 34348 33324 34360
rect 33376 34388 33382 34400
rect 33870 34388 33876 34400
rect 33376 34360 33876 34388
rect 33376 34348 33382 34360
rect 33870 34348 33876 34360
rect 33928 34348 33934 34400
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 5442 34144 5448 34196
rect 5500 34184 5506 34196
rect 5721 34187 5779 34193
rect 5721 34184 5733 34187
rect 5500 34156 5733 34184
rect 5500 34144 5506 34156
rect 5721 34153 5733 34156
rect 5767 34153 5779 34187
rect 11054 34184 11060 34196
rect 11015 34156 11060 34184
rect 5721 34147 5779 34153
rect 11054 34144 11060 34156
rect 11112 34144 11118 34196
rect 14550 34144 14556 34196
rect 14608 34184 14614 34196
rect 14608 34156 14653 34184
rect 14608 34144 14614 34156
rect 15102 34144 15108 34196
rect 15160 34184 15166 34196
rect 18509 34187 18567 34193
rect 15160 34156 18184 34184
rect 15160 34144 15166 34156
rect 5074 34116 5080 34128
rect 4080 34088 5080 34116
rect 4080 33989 4108 34088
rect 5074 34076 5080 34088
rect 5132 34076 5138 34128
rect 13541 34119 13599 34125
rect 13541 34085 13553 34119
rect 13587 34116 13599 34119
rect 14274 34116 14280 34128
rect 13587 34088 14280 34116
rect 13587 34085 13599 34088
rect 13541 34079 13599 34085
rect 14274 34076 14280 34088
rect 14332 34076 14338 34128
rect 17310 34076 17316 34128
rect 17368 34076 17374 34128
rect 4890 34048 4896 34060
rect 4172 34020 4896 34048
rect 4172 33989 4200 34020
rect 4890 34008 4896 34020
rect 4948 34048 4954 34060
rect 6730 34048 6736 34060
rect 4948 34020 6736 34048
rect 4948 34008 4954 34020
rect 6730 34008 6736 34020
rect 6788 34008 6794 34060
rect 10042 34008 10048 34060
rect 10100 34048 10106 34060
rect 17328 34048 17356 34076
rect 10100 34020 10732 34048
rect 17328 34020 17724 34048
rect 10100 34008 10106 34020
rect 4065 33983 4123 33989
rect 4065 33949 4077 33983
rect 4111 33949 4123 33983
rect 4065 33943 4123 33949
rect 4157 33983 4215 33989
rect 4157 33949 4169 33983
rect 4203 33949 4215 33983
rect 4157 33943 4215 33949
rect 4249 33983 4307 33989
rect 4249 33949 4261 33983
rect 4295 33949 4307 33983
rect 4249 33943 4307 33949
rect 4433 33983 4491 33989
rect 4433 33949 4445 33983
rect 4479 33980 4491 33983
rect 5442 33980 5448 33992
rect 4479 33952 5448 33980
rect 4479 33949 4491 33952
rect 4433 33943 4491 33949
rect 4264 33912 4292 33943
rect 5442 33940 5448 33952
rect 5500 33940 5506 33992
rect 10134 33940 10140 33992
rect 10192 33980 10198 33992
rect 10594 33989 10600 33992
rect 10413 33983 10471 33989
rect 10413 33980 10425 33983
rect 10192 33952 10425 33980
rect 10192 33940 10198 33952
rect 10413 33949 10425 33952
rect 10459 33949 10471 33983
rect 10413 33943 10471 33949
rect 10576 33983 10600 33989
rect 10576 33949 10588 33983
rect 10576 33943 10600 33949
rect 10594 33940 10600 33943
rect 10652 33940 10658 33992
rect 10704 33989 10732 34020
rect 10689 33983 10747 33989
rect 10689 33949 10701 33983
rect 10735 33949 10747 33983
rect 10689 33943 10747 33949
rect 10827 33983 10885 33989
rect 10827 33949 10839 33983
rect 10873 33980 10885 33983
rect 11514 33980 11520 33992
rect 10873 33952 11520 33980
rect 10873 33949 10885 33952
rect 10827 33943 10885 33949
rect 11514 33940 11520 33952
rect 11572 33940 11578 33992
rect 13357 33983 13415 33989
rect 13357 33949 13369 33983
rect 13403 33980 13415 33983
rect 14918 33980 14924 33992
rect 13403 33952 14924 33980
rect 13403 33949 13415 33952
rect 13357 33943 13415 33949
rect 4893 33915 4951 33921
rect 4893 33912 4905 33915
rect 4264 33884 4905 33912
rect 4893 33881 4905 33884
rect 4939 33881 4951 33915
rect 5074 33912 5080 33924
rect 5035 33884 5080 33912
rect 4893 33875 4951 33881
rect 5074 33872 5080 33884
rect 5132 33872 5138 33924
rect 5261 33915 5319 33921
rect 5261 33881 5273 33915
rect 5307 33912 5319 33915
rect 5534 33912 5540 33924
rect 5307 33884 5540 33912
rect 5307 33881 5319 33884
rect 5261 33875 5319 33881
rect 5534 33872 5540 33884
rect 5592 33912 5598 33924
rect 6362 33912 6368 33924
rect 5592 33884 6368 33912
rect 5592 33872 5598 33884
rect 6362 33872 6368 33884
rect 6420 33872 6426 33924
rect 3786 33844 3792 33856
rect 3747 33816 3792 33844
rect 3786 33804 3792 33816
rect 3844 33804 3850 33856
rect 7374 33804 7380 33856
rect 7432 33844 7438 33856
rect 7561 33847 7619 33853
rect 7561 33844 7573 33847
rect 7432 33816 7573 33844
rect 7432 33804 7438 33816
rect 7561 33813 7573 33816
rect 7607 33844 7619 33847
rect 8110 33844 8116 33856
rect 7607 33816 8116 33844
rect 7607 33813 7619 33816
rect 7561 33807 7619 33813
rect 8110 33804 8116 33816
rect 8168 33804 8174 33856
rect 8386 33804 8392 33856
rect 8444 33844 8450 33856
rect 13372 33844 13400 33943
rect 14918 33940 14924 33952
rect 14976 33940 14982 33992
rect 16853 33983 16911 33989
rect 16853 33949 16865 33983
rect 16899 33980 16911 33983
rect 17034 33980 17040 33992
rect 16899 33952 17040 33980
rect 16899 33949 16911 33952
rect 16853 33943 16911 33949
rect 17034 33940 17040 33952
rect 17092 33980 17098 33992
rect 17092 33952 17448 33980
rect 17092 33940 17098 33952
rect 14642 33912 14648 33924
rect 14603 33884 14648 33912
rect 14642 33872 14648 33884
rect 14700 33872 14706 33924
rect 16597 33915 16655 33921
rect 16597 33881 16609 33915
rect 16643 33912 16655 33915
rect 17313 33915 17371 33921
rect 17313 33912 17325 33915
rect 16643 33884 17325 33912
rect 16643 33881 16655 33884
rect 16597 33875 16655 33881
rect 17313 33881 17325 33884
rect 17359 33881 17371 33915
rect 17420 33912 17448 33952
rect 17494 33940 17500 33992
rect 17552 33980 17558 33992
rect 17696 33989 17724 34020
rect 17862 34008 17868 34060
rect 17920 34048 17926 34060
rect 17920 34020 18000 34048
rect 17920 34008 17926 34020
rect 17589 33983 17647 33989
rect 17589 33980 17601 33983
rect 17552 33952 17601 33980
rect 17552 33940 17558 33952
rect 17589 33949 17601 33952
rect 17635 33949 17647 33983
rect 17589 33943 17647 33949
rect 17681 33983 17739 33989
rect 17681 33949 17693 33983
rect 17727 33949 17739 33983
rect 17681 33943 17739 33949
rect 17770 33940 17776 33992
rect 17828 33980 17834 33992
rect 17972 33989 18000 34020
rect 17957 33983 18015 33989
rect 17828 33952 17873 33980
rect 17828 33940 17834 33952
rect 17957 33949 17969 33983
rect 18003 33949 18015 33983
rect 18156 33980 18184 34156
rect 18509 34153 18521 34187
rect 18555 34184 18567 34187
rect 18598 34184 18604 34196
rect 18555 34156 18604 34184
rect 18555 34153 18567 34156
rect 18509 34147 18567 34153
rect 18598 34144 18604 34156
rect 18656 34144 18662 34196
rect 21818 34184 21824 34196
rect 21779 34156 21824 34184
rect 21818 34144 21824 34156
rect 21876 34144 21882 34196
rect 25866 34184 25872 34196
rect 25827 34156 25872 34184
rect 25866 34144 25872 34156
rect 25924 34144 25930 34196
rect 34790 34144 34796 34196
rect 34848 34184 34854 34196
rect 35069 34187 35127 34193
rect 35069 34184 35081 34187
rect 34848 34156 35081 34184
rect 34848 34144 34854 34156
rect 35069 34153 35081 34156
rect 35115 34153 35127 34187
rect 35069 34147 35127 34153
rect 33686 34116 33692 34128
rect 32692 34088 33692 34116
rect 18506 34008 18512 34060
rect 18564 34048 18570 34060
rect 20438 34048 20444 34060
rect 18564 34020 19472 34048
rect 18564 34008 18570 34020
rect 19444 33989 19472 34020
rect 19628 34020 20444 34048
rect 19337 33983 19395 33989
rect 19337 33980 19349 33983
rect 18156 33952 19349 33980
rect 17957 33943 18015 33949
rect 19337 33949 19349 33952
rect 19383 33949 19395 33983
rect 19337 33943 19395 33949
rect 19430 33983 19488 33989
rect 19430 33949 19442 33983
rect 19476 33949 19488 33983
rect 19430 33943 19488 33949
rect 17862 33912 17868 33924
rect 17420 33884 17868 33912
rect 17313 33875 17371 33881
rect 17862 33872 17868 33884
rect 17920 33872 17926 33924
rect 19628 33921 19656 34020
rect 20438 34008 20444 34020
rect 20496 34008 20502 34060
rect 22002 34008 22008 34060
rect 22060 34048 22066 34060
rect 22281 34051 22339 34057
rect 22281 34048 22293 34051
rect 22060 34020 22293 34048
rect 22060 34008 22066 34020
rect 22281 34017 22293 34020
rect 22327 34017 22339 34051
rect 22281 34011 22339 34017
rect 29730 34008 29736 34060
rect 29788 34048 29794 34060
rect 30193 34051 30251 34057
rect 30193 34048 30205 34051
rect 29788 34020 30205 34048
rect 29788 34008 29794 34020
rect 30193 34017 30205 34020
rect 30239 34048 30251 34051
rect 30742 34048 30748 34060
rect 30239 34020 30748 34048
rect 30239 34017 30251 34020
rect 30193 34011 30251 34017
rect 30742 34008 30748 34020
rect 30800 34008 30806 34060
rect 19794 33940 19800 33992
rect 19852 33989 19858 33992
rect 19852 33980 19860 33989
rect 22548 33983 22606 33989
rect 19852 33952 19897 33980
rect 19852 33943 19860 33952
rect 22548 33949 22560 33983
rect 22594 33980 22606 33983
rect 22830 33980 22836 33992
rect 22594 33952 22836 33980
rect 22594 33949 22606 33952
rect 22548 33943 22606 33949
rect 19852 33940 19858 33943
rect 22830 33940 22836 33952
rect 22888 33940 22894 33992
rect 23474 33940 23480 33992
rect 23532 33980 23538 33992
rect 24857 33983 24915 33989
rect 24857 33980 24869 33983
rect 23532 33952 24869 33980
rect 23532 33940 23538 33952
rect 24857 33949 24869 33952
rect 24903 33949 24915 33983
rect 24857 33943 24915 33949
rect 26973 33983 27031 33989
rect 26973 33949 26985 33983
rect 27019 33980 27031 33983
rect 27062 33980 27068 33992
rect 27019 33952 27068 33980
rect 27019 33949 27031 33952
rect 26973 33943 27031 33949
rect 27062 33940 27068 33952
rect 27120 33940 27126 33992
rect 28997 33983 29055 33989
rect 28997 33949 29009 33983
rect 29043 33980 29055 33983
rect 29914 33980 29920 33992
rect 29043 33952 29920 33980
rect 29043 33949 29055 33952
rect 28997 33943 29055 33949
rect 29914 33940 29920 33952
rect 29972 33980 29978 33992
rect 30374 33980 30380 33992
rect 29972 33952 30380 33980
rect 29972 33940 29978 33952
rect 30374 33940 30380 33952
rect 30432 33940 30438 33992
rect 32692 33989 32720 34088
rect 33686 34076 33692 34088
rect 33744 34116 33750 34128
rect 33744 34088 34560 34116
rect 33744 34076 33750 34088
rect 33045 34051 33103 34057
rect 33045 34017 33057 34051
rect 33091 34048 33103 34051
rect 33962 34048 33968 34060
rect 33091 34020 33732 34048
rect 33091 34017 33103 34020
rect 33045 34011 33103 34017
rect 32677 33983 32735 33989
rect 32677 33949 32689 33983
rect 32723 33949 32735 33983
rect 33502 33980 33508 33992
rect 33463 33952 33508 33980
rect 32677 33943 32735 33949
rect 33502 33940 33508 33952
rect 33560 33940 33566 33992
rect 33704 33989 33732 34020
rect 33796 34020 33968 34048
rect 33796 33989 33824 34020
rect 33962 34008 33968 34020
rect 34020 34008 34026 34060
rect 33689 33983 33747 33989
rect 33689 33949 33701 33983
rect 33735 33949 33747 33983
rect 33689 33943 33747 33949
rect 33781 33983 33839 33989
rect 33781 33949 33793 33983
rect 33827 33949 33839 33983
rect 33781 33943 33839 33949
rect 33870 33940 33876 33992
rect 33928 33980 33934 33992
rect 33928 33952 33973 33980
rect 33928 33940 33934 33952
rect 19613 33915 19671 33921
rect 19613 33881 19625 33915
rect 19659 33881 19671 33915
rect 19613 33875 19671 33881
rect 19705 33915 19763 33921
rect 19705 33881 19717 33915
rect 19751 33912 19763 33915
rect 20254 33912 20260 33924
rect 19751 33884 20260 33912
rect 19751 33881 19763 33884
rect 19705 33875 19763 33881
rect 8444 33816 13400 33844
rect 15473 33847 15531 33853
rect 8444 33804 8450 33816
rect 15473 33813 15485 33847
rect 15519 33844 15531 33847
rect 15930 33844 15936 33856
rect 15519 33816 15936 33844
rect 15519 33813 15531 33816
rect 15473 33807 15531 33813
rect 15930 33804 15936 33816
rect 15988 33804 15994 33856
rect 16942 33804 16948 33856
rect 17000 33844 17006 33856
rect 19628 33844 19656 33875
rect 20254 33872 20260 33884
rect 20312 33872 20318 33924
rect 21450 33912 21456 33924
rect 21411 33884 21456 33912
rect 21450 33872 21456 33884
rect 21508 33872 21514 33924
rect 21637 33915 21695 33921
rect 21637 33881 21649 33915
rect 21683 33912 21695 33915
rect 25038 33912 25044 33924
rect 21683 33884 22094 33912
rect 24999 33884 25044 33912
rect 21683 33881 21695 33884
rect 21637 33875 21695 33881
rect 19978 33844 19984 33856
rect 17000 33816 19656 33844
rect 19939 33816 19984 33844
rect 17000 33804 17006 33816
rect 19978 33804 19984 33816
rect 20036 33804 20042 33856
rect 22066 33844 22094 33884
rect 25038 33872 25044 33884
rect 25096 33872 25102 33924
rect 27246 33921 27252 33924
rect 27240 33875 27252 33921
rect 27304 33912 27310 33924
rect 31202 33912 31208 33924
rect 27304 33884 27340 33912
rect 31163 33884 31208 33912
rect 27246 33872 27252 33875
rect 27304 33872 27310 33884
rect 31202 33872 31208 33884
rect 31260 33872 31266 33924
rect 31386 33912 31392 33924
rect 31347 33884 31392 33912
rect 31386 33872 31392 33884
rect 31444 33872 31450 33924
rect 32861 33915 32919 33921
rect 32861 33881 32873 33915
rect 32907 33912 32919 33915
rect 34422 33912 34428 33924
rect 32907 33884 34428 33912
rect 32907 33881 32919 33884
rect 32861 33875 32919 33881
rect 34422 33872 34428 33884
rect 34480 33872 34486 33924
rect 34532 33912 34560 34088
rect 34606 33940 34612 33992
rect 34664 33980 34670 33992
rect 34885 33983 34943 33989
rect 34885 33980 34897 33983
rect 34664 33952 34897 33980
rect 34664 33940 34670 33952
rect 34885 33949 34897 33952
rect 34931 33949 34943 33983
rect 34885 33943 34943 33949
rect 34701 33915 34759 33921
rect 34701 33912 34713 33915
rect 34532 33884 34713 33912
rect 34701 33881 34713 33884
rect 34747 33881 34759 33915
rect 34701 33875 34759 33881
rect 23661 33847 23719 33853
rect 23661 33844 23673 33847
rect 22066 33816 23673 33844
rect 23661 33813 23673 33816
rect 23707 33844 23719 33847
rect 24486 33844 24492 33856
rect 23707 33816 24492 33844
rect 23707 33813 23719 33816
rect 23661 33807 23719 33813
rect 24486 33804 24492 33816
rect 24544 33804 24550 33856
rect 25222 33844 25228 33856
rect 25183 33816 25228 33844
rect 25222 33804 25228 33816
rect 25280 33804 25286 33856
rect 28350 33844 28356 33856
rect 28311 33816 28356 33844
rect 28350 33804 28356 33816
rect 28408 33804 28414 33856
rect 30558 33804 30564 33856
rect 30616 33844 30622 33856
rect 31573 33847 31631 33853
rect 31573 33844 31585 33847
rect 30616 33816 31585 33844
rect 30616 33804 30622 33816
rect 31573 33813 31585 33816
rect 31619 33813 31631 33847
rect 34146 33844 34152 33856
rect 34107 33816 34152 33844
rect 31573 33807 31631 33813
rect 34146 33804 34152 33816
rect 34204 33804 34210 33856
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 4433 33643 4491 33649
rect 4433 33609 4445 33643
rect 4479 33640 4491 33643
rect 4706 33640 4712 33652
rect 4479 33612 4712 33640
rect 4479 33609 4491 33612
rect 4433 33603 4491 33609
rect 4706 33600 4712 33612
rect 4764 33600 4770 33652
rect 5166 33600 5172 33652
rect 5224 33640 5230 33652
rect 5261 33643 5319 33649
rect 5261 33640 5273 33643
rect 5224 33612 5273 33640
rect 5224 33600 5230 33612
rect 5261 33609 5273 33612
rect 5307 33609 5319 33643
rect 5261 33603 5319 33609
rect 6454 33600 6460 33652
rect 6512 33640 6518 33652
rect 7098 33640 7104 33652
rect 6512 33612 7104 33640
rect 6512 33600 6518 33612
rect 7098 33600 7104 33612
rect 7156 33600 7162 33652
rect 8018 33640 8024 33652
rect 7979 33612 8024 33640
rect 8018 33600 8024 33612
rect 8076 33600 8082 33652
rect 8110 33600 8116 33652
rect 8168 33640 8174 33652
rect 17037 33643 17095 33649
rect 8168 33612 12434 33640
rect 8168 33600 8174 33612
rect 2860 33575 2918 33581
rect 2860 33541 2872 33575
rect 2906 33572 2918 33575
rect 3786 33572 3792 33584
rect 2906 33544 3792 33572
rect 2906 33541 2918 33544
rect 2860 33535 2918 33541
rect 3786 33532 3792 33544
rect 3844 33532 3850 33584
rect 4614 33572 4620 33584
rect 4527 33544 4620 33572
rect 4614 33532 4620 33544
rect 4672 33572 4678 33584
rect 5350 33572 5356 33584
rect 4672 33544 5356 33572
rect 4672 33532 4678 33544
rect 5350 33532 5356 33544
rect 5408 33532 5414 33584
rect 12406 33572 12434 33612
rect 17037 33609 17049 33643
rect 17083 33640 17095 33643
rect 17770 33640 17776 33652
rect 17083 33612 17776 33640
rect 17083 33609 17095 33612
rect 17037 33603 17095 33609
rect 17770 33600 17776 33612
rect 17828 33600 17834 33652
rect 27246 33640 27252 33652
rect 27207 33612 27252 33640
rect 27246 33600 27252 33612
rect 27304 33600 27310 33652
rect 30650 33640 30656 33652
rect 30116 33612 30656 33640
rect 13906 33572 13912 33584
rect 12406 33544 13912 33572
rect 13906 33532 13912 33544
rect 13964 33532 13970 33584
rect 14124 33575 14182 33581
rect 14124 33541 14136 33575
rect 14170 33572 14182 33575
rect 14829 33575 14887 33581
rect 14829 33572 14841 33575
rect 14170 33544 14841 33572
rect 14170 33541 14182 33544
rect 14124 33535 14182 33541
rect 14829 33541 14841 33544
rect 14875 33541 14887 33575
rect 14829 33535 14887 33541
rect 14918 33532 14924 33584
rect 14976 33572 14982 33584
rect 14976 33544 15240 33572
rect 14976 33532 14982 33544
rect 2590 33504 2596 33516
rect 2551 33476 2596 33504
rect 2590 33464 2596 33476
rect 2648 33464 2654 33516
rect 4801 33507 4859 33513
rect 4801 33473 4813 33507
rect 4847 33504 4859 33507
rect 5534 33504 5540 33516
rect 4847 33476 5540 33504
rect 4847 33473 4859 33476
rect 4801 33467 4859 33473
rect 5534 33464 5540 33476
rect 5592 33464 5598 33516
rect 6914 33513 6920 33516
rect 6908 33467 6920 33513
rect 6972 33504 6978 33516
rect 6972 33476 7008 33504
rect 6914 33464 6920 33467
rect 6972 33464 6978 33476
rect 11698 33464 11704 33516
rect 11756 33504 11762 33516
rect 12437 33507 12495 33513
rect 12437 33504 12449 33507
rect 11756 33476 12449 33504
rect 11756 33464 11762 33476
rect 12437 33473 12449 33476
rect 12483 33473 12495 33507
rect 12437 33467 12495 33473
rect 15010 33464 15016 33516
rect 15068 33504 15074 33516
rect 15212 33513 15240 33544
rect 15930 33532 15936 33584
rect 15988 33572 15994 33584
rect 16298 33572 16304 33584
rect 15988 33544 16304 33572
rect 15988 33532 15994 33544
rect 16298 33532 16304 33544
rect 16356 33572 16362 33584
rect 16853 33575 16911 33581
rect 16853 33572 16865 33575
rect 16356 33544 16865 33572
rect 16356 33532 16362 33544
rect 16853 33541 16865 33544
rect 16899 33541 16911 33575
rect 19150 33572 19156 33584
rect 19111 33544 19156 33572
rect 16853 33535 16911 33541
rect 19150 33532 19156 33544
rect 19208 33532 19214 33584
rect 22088 33575 22146 33581
rect 22088 33541 22100 33575
rect 22134 33572 22146 33575
rect 23937 33575 23995 33581
rect 23937 33572 23949 33575
rect 22134 33544 23949 33572
rect 22134 33541 22146 33544
rect 22088 33535 22146 33541
rect 23937 33541 23949 33544
rect 23983 33541 23995 33575
rect 24670 33572 24676 33584
rect 23937 33535 23995 33541
rect 24320 33544 24676 33572
rect 15105 33507 15163 33513
rect 15105 33504 15117 33507
rect 15068 33476 15117 33504
rect 15068 33464 15074 33476
rect 15105 33473 15117 33476
rect 15151 33473 15163 33507
rect 15105 33467 15163 33473
rect 15197 33507 15255 33513
rect 15197 33473 15209 33507
rect 15243 33473 15255 33507
rect 15197 33467 15255 33473
rect 15286 33464 15292 33516
rect 15344 33504 15350 33516
rect 15344 33476 15389 33504
rect 15344 33464 15350 33476
rect 15470 33464 15476 33516
rect 15528 33504 15534 33516
rect 15528 33476 15573 33504
rect 15528 33464 15534 33476
rect 16482 33464 16488 33516
rect 16540 33504 16546 33516
rect 16669 33507 16727 33513
rect 16669 33504 16681 33507
rect 16540 33476 16681 33504
rect 16540 33464 16546 33476
rect 16669 33473 16681 33476
rect 16715 33473 16727 33507
rect 16669 33467 16727 33473
rect 17865 33507 17923 33513
rect 17865 33473 17877 33507
rect 17911 33504 17923 33507
rect 18509 33507 18567 33513
rect 18509 33504 18521 33507
rect 17911 33476 18521 33504
rect 17911 33473 17923 33476
rect 17865 33467 17923 33473
rect 18509 33473 18521 33476
rect 18555 33504 18567 33507
rect 19337 33507 19395 33513
rect 19337 33504 19349 33507
rect 18555 33476 19349 33504
rect 18555 33473 18567 33476
rect 18509 33467 18567 33473
rect 19337 33473 19349 33476
rect 19383 33504 19395 33507
rect 21821 33507 21879 33513
rect 19383 33476 20024 33504
rect 19383 33473 19395 33476
rect 19337 33467 19395 33473
rect 6641 33439 6699 33445
rect 6641 33405 6653 33439
rect 6687 33405 6699 33439
rect 6641 33399 6699 33405
rect 14369 33439 14427 33445
rect 14369 33405 14381 33439
rect 14415 33436 14427 33439
rect 17034 33436 17040 33448
rect 14415 33408 17040 33436
rect 14415 33405 14427 33408
rect 14369 33399 14427 33405
rect 3973 33303 4031 33309
rect 3973 33269 3985 33303
rect 4019 33300 4031 33303
rect 5074 33300 5080 33312
rect 4019 33272 5080 33300
rect 4019 33269 4031 33272
rect 3973 33263 4031 33269
rect 5074 33260 5080 33272
rect 5132 33260 5138 33312
rect 6656 33300 6684 33399
rect 17034 33396 17040 33408
rect 17092 33396 17098 33448
rect 8662 33328 8668 33380
rect 8720 33368 8726 33380
rect 12253 33371 12311 33377
rect 12253 33368 12265 33371
rect 8720 33340 12265 33368
rect 8720 33328 8726 33340
rect 12253 33337 12265 33340
rect 12299 33368 12311 33371
rect 18322 33368 18328 33380
rect 12299 33340 13124 33368
rect 18283 33340 18328 33368
rect 12299 33337 12311 33340
rect 12253 33331 12311 33337
rect 7006 33300 7012 33312
rect 6656 33272 7012 33300
rect 7006 33260 7012 33272
rect 7064 33260 7070 33312
rect 10962 33260 10968 33312
rect 11020 33300 11026 33312
rect 11517 33303 11575 33309
rect 11517 33300 11529 33303
rect 11020 33272 11529 33300
rect 11020 33260 11026 33272
rect 11517 33269 11529 33272
rect 11563 33269 11575 33303
rect 12986 33300 12992 33312
rect 12947 33272 12992 33300
rect 11517 33263 11575 33269
rect 12986 33260 12992 33272
rect 13044 33260 13050 33312
rect 13096 33300 13124 33340
rect 18322 33328 18328 33340
rect 18380 33328 18386 33380
rect 16942 33300 16948 33312
rect 13096 33272 16948 33300
rect 16942 33260 16948 33272
rect 17000 33260 17006 33312
rect 19996 33309 20024 33476
rect 21821 33473 21833 33507
rect 21867 33504 21879 33507
rect 21910 33504 21916 33516
rect 21867 33476 21916 33504
rect 21867 33473 21879 33476
rect 21821 33467 21879 33473
rect 21910 33464 21916 33476
rect 21968 33464 21974 33516
rect 24320 33513 24348 33544
rect 24670 33532 24676 33544
rect 24728 33572 24734 33584
rect 24728 33544 25360 33572
rect 24728 33532 24734 33544
rect 24213 33507 24271 33513
rect 24213 33473 24225 33507
rect 24259 33473 24271 33507
rect 24213 33467 24271 33473
rect 24305 33507 24363 33513
rect 24305 33473 24317 33507
rect 24351 33473 24363 33507
rect 24305 33467 24363 33473
rect 24228 33436 24256 33467
rect 24394 33464 24400 33516
rect 24452 33504 24458 33516
rect 24581 33507 24639 33513
rect 24452 33476 24497 33504
rect 24452 33464 24458 33476
rect 24581 33473 24593 33507
rect 24627 33504 24639 33507
rect 24946 33504 24952 33516
rect 24627 33476 24952 33504
rect 24627 33473 24639 33476
rect 24581 33467 24639 33473
rect 24946 33464 24952 33476
rect 25004 33504 25010 33516
rect 25041 33507 25099 33513
rect 25041 33504 25053 33507
rect 25004 33476 25053 33504
rect 25004 33464 25010 33476
rect 25041 33473 25053 33476
rect 25087 33473 25099 33507
rect 25222 33504 25228 33516
rect 25183 33476 25228 33504
rect 25041 33467 25099 33473
rect 25222 33464 25228 33476
rect 25280 33464 25286 33516
rect 25332 33513 25360 33544
rect 25317 33507 25375 33513
rect 25317 33473 25329 33507
rect 25363 33473 25375 33507
rect 25317 33467 25375 33473
rect 25455 33507 25513 33513
rect 25455 33473 25467 33507
rect 25501 33504 25513 33507
rect 25866 33504 25872 33516
rect 25501 33476 25872 33504
rect 25501 33473 25513 33476
rect 25455 33467 25513 33473
rect 25866 33464 25872 33476
rect 25924 33464 25930 33516
rect 27525 33507 27583 33513
rect 27525 33473 27537 33507
rect 27571 33473 27583 33507
rect 27525 33467 27583 33473
rect 27617 33507 27675 33513
rect 27617 33473 27629 33507
rect 27663 33473 27675 33507
rect 27617 33467 27675 33473
rect 24762 33436 24768 33448
rect 24228 33408 24768 33436
rect 24762 33396 24768 33408
rect 24820 33396 24826 33448
rect 23842 33368 23848 33380
rect 23124 33340 23848 33368
rect 19981 33303 20039 33309
rect 19981 33269 19993 33303
rect 20027 33300 20039 33303
rect 23124 33300 23152 33340
rect 23842 33328 23848 33340
rect 23900 33368 23906 33380
rect 24302 33368 24308 33380
rect 23900 33340 24308 33368
rect 23900 33328 23906 33340
rect 24302 33328 24308 33340
rect 24360 33328 24366 33380
rect 25685 33371 25743 33377
rect 25685 33337 25697 33371
rect 25731 33368 25743 33371
rect 26878 33368 26884 33380
rect 25731 33340 26884 33368
rect 25731 33337 25743 33340
rect 25685 33331 25743 33337
rect 26878 33328 26884 33340
rect 26936 33328 26942 33380
rect 20027 33272 23152 33300
rect 23201 33303 23259 33309
rect 20027 33269 20039 33272
rect 19981 33263 20039 33269
rect 23201 33269 23213 33303
rect 23247 33300 23259 33303
rect 23658 33300 23664 33312
rect 23247 33272 23664 33300
rect 23247 33269 23259 33272
rect 23201 33263 23259 33269
rect 23658 33260 23664 33272
rect 23716 33260 23722 33312
rect 26234 33260 26240 33312
rect 26292 33300 26298 33312
rect 26329 33303 26387 33309
rect 26329 33300 26341 33303
rect 26292 33272 26341 33300
rect 26292 33260 26298 33272
rect 26329 33269 26341 33272
rect 26375 33300 26387 33303
rect 26970 33300 26976 33312
rect 26375 33272 26976 33300
rect 26375 33269 26387 33272
rect 26329 33263 26387 33269
rect 26970 33260 26976 33272
rect 27028 33300 27034 33312
rect 27540 33300 27568 33467
rect 27632 33436 27660 33467
rect 27706 33464 27712 33516
rect 27764 33504 27770 33516
rect 27893 33507 27951 33513
rect 27764 33476 27809 33504
rect 27764 33464 27770 33476
rect 27893 33473 27905 33507
rect 27939 33504 27951 33507
rect 28166 33504 28172 33516
rect 27939 33476 28172 33504
rect 27939 33473 27951 33476
rect 27893 33467 27951 33473
rect 28166 33464 28172 33476
rect 28224 33464 28230 33516
rect 29546 33464 29552 33516
rect 29604 33504 29610 33516
rect 30116 33504 30144 33612
rect 30650 33600 30656 33612
rect 30708 33600 30714 33652
rect 34422 33600 34428 33652
rect 34480 33640 34486 33652
rect 34517 33643 34575 33649
rect 34517 33640 34529 33643
rect 34480 33612 34529 33640
rect 34480 33600 34486 33612
rect 34517 33609 34529 33612
rect 34563 33609 34575 33643
rect 34517 33603 34575 33609
rect 31389 33575 31447 33581
rect 31389 33541 31401 33575
rect 31435 33572 31447 33575
rect 32306 33572 32312 33584
rect 31435 33544 32312 33572
rect 31435 33541 31447 33544
rect 31389 33535 31447 33541
rect 32306 33532 32312 33544
rect 32364 33532 32370 33584
rect 34146 33532 34152 33584
rect 34204 33572 34210 33584
rect 35630 33575 35688 33581
rect 35630 33572 35642 33575
rect 34204 33544 35642 33572
rect 34204 33532 34210 33544
rect 35630 33541 35642 33544
rect 35676 33541 35688 33575
rect 35630 33535 35688 33541
rect 30377 33507 30435 33513
rect 30377 33504 30389 33507
rect 29604 33476 30389 33504
rect 29604 33464 29610 33476
rect 30377 33473 30389 33476
rect 30423 33473 30435 33507
rect 30377 33467 30435 33473
rect 30469 33507 30527 33513
rect 30469 33473 30481 33507
rect 30515 33473 30527 33507
rect 30469 33467 30527 33473
rect 30282 33436 30288 33448
rect 27632 33408 30288 33436
rect 30282 33396 30288 33408
rect 30340 33436 30346 33448
rect 30484 33436 30512 33467
rect 30558 33464 30564 33516
rect 30616 33504 30622 33516
rect 30616 33476 30661 33504
rect 30616 33464 30622 33476
rect 30742 33464 30748 33516
rect 30800 33504 30806 33516
rect 30800 33476 30845 33504
rect 30800 33464 30806 33476
rect 31662 33464 31668 33516
rect 31720 33504 31726 33516
rect 32950 33513 32956 33516
rect 32677 33507 32735 33513
rect 32677 33504 32689 33507
rect 31720 33476 32689 33504
rect 31720 33464 31726 33476
rect 32677 33473 32689 33476
rect 32723 33473 32735 33507
rect 32677 33467 32735 33473
rect 32944 33467 32956 33513
rect 33008 33504 33014 33516
rect 33008 33476 33044 33504
rect 32950 33464 32956 33467
rect 33008 33464 33014 33476
rect 30340 33408 30512 33436
rect 35897 33439 35955 33445
rect 30340 33396 30346 33408
rect 35897 33405 35909 33439
rect 35943 33436 35955 33439
rect 36078 33436 36084 33448
rect 35943 33408 36084 33436
rect 35943 33405 35955 33408
rect 35897 33399 35955 33405
rect 36078 33396 36084 33408
rect 36136 33396 36142 33448
rect 31110 33328 31116 33380
rect 31168 33368 31174 33380
rect 31205 33371 31263 33377
rect 31205 33368 31217 33371
rect 31168 33340 31217 33368
rect 31168 33328 31174 33340
rect 31205 33337 31217 33340
rect 31251 33337 31263 33371
rect 58158 33368 58164 33380
rect 58119 33340 58164 33368
rect 31205 33331 31263 33337
rect 58158 33328 58164 33340
rect 58216 33328 58222 33380
rect 29546 33300 29552 33312
rect 27028 33272 27568 33300
rect 29507 33272 29552 33300
rect 27028 33260 27034 33272
rect 29546 33260 29552 33272
rect 29604 33260 29610 33312
rect 30098 33300 30104 33312
rect 30059 33272 30104 33300
rect 30098 33260 30104 33272
rect 30156 33260 30162 33312
rect 34057 33303 34115 33309
rect 34057 33269 34069 33303
rect 34103 33300 34115 33303
rect 34146 33300 34152 33312
rect 34103 33272 34152 33300
rect 34103 33269 34115 33272
rect 34057 33263 34115 33269
rect 34146 33260 34152 33272
rect 34204 33260 34210 33312
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 5258 33056 5264 33108
rect 5316 33096 5322 33108
rect 5537 33099 5595 33105
rect 5537 33096 5549 33099
rect 5316 33068 5549 33096
rect 5316 33056 5322 33068
rect 5537 33065 5549 33068
rect 5583 33065 5595 33099
rect 5537 33059 5595 33065
rect 6733 33099 6791 33105
rect 6733 33065 6745 33099
rect 6779 33096 6791 33099
rect 6914 33096 6920 33108
rect 6779 33068 6920 33096
rect 6779 33065 6791 33068
rect 6733 33059 6791 33065
rect 6914 33056 6920 33068
rect 6972 33056 6978 33108
rect 13541 33099 13599 33105
rect 13541 33065 13553 33099
rect 13587 33096 13599 33099
rect 15286 33096 15292 33108
rect 13587 33068 15292 33096
rect 13587 33065 13599 33068
rect 13541 33059 13599 33065
rect 15286 33056 15292 33068
rect 15344 33056 15350 33108
rect 17954 33056 17960 33108
rect 18012 33096 18018 33108
rect 20346 33096 20352 33108
rect 18012 33068 20352 33096
rect 18012 33056 18018 33068
rect 20346 33056 20352 33068
rect 20404 33056 20410 33108
rect 23845 33099 23903 33105
rect 23845 33065 23857 33099
rect 23891 33096 23903 33099
rect 24394 33096 24400 33108
rect 23891 33068 24400 33096
rect 23891 33065 23903 33068
rect 23845 33059 23903 33065
rect 24394 33056 24400 33068
rect 24452 33056 24458 33108
rect 26234 33056 26240 33108
rect 26292 33056 26298 33108
rect 27709 33099 27767 33105
rect 27709 33065 27721 33099
rect 27755 33096 27767 33099
rect 28166 33096 28172 33108
rect 27755 33068 28172 33096
rect 27755 33065 27767 33068
rect 27709 33059 27767 33065
rect 28166 33056 28172 33068
rect 28224 33056 28230 33108
rect 4982 32988 4988 33040
rect 5040 33028 5046 33040
rect 5040 33000 9720 33028
rect 5040 32988 5046 33000
rect 9692 32969 9720 33000
rect 17218 32988 17224 33040
rect 17276 33028 17282 33040
rect 26252 33028 26280 33056
rect 17276 33000 26280 33028
rect 17276 32988 17282 33000
rect 7837 32963 7895 32969
rect 7837 32960 7849 32963
rect 7208 32932 7849 32960
rect 6638 32892 6644 32904
rect 6196 32864 6644 32892
rect 5718 32716 5724 32768
rect 5776 32756 5782 32768
rect 6196 32765 6224 32864
rect 6638 32852 6644 32864
rect 6696 32892 6702 32904
rect 7208 32901 7236 32932
rect 7837 32929 7849 32932
rect 7883 32929 7895 32963
rect 7837 32923 7895 32929
rect 9677 32963 9735 32969
rect 9677 32929 9689 32963
rect 9723 32960 9735 32963
rect 9858 32960 9864 32972
rect 9723 32932 9864 32960
rect 9723 32929 9735 32932
rect 9677 32923 9735 32929
rect 9858 32920 9864 32932
rect 9916 32920 9922 32972
rect 14369 32963 14427 32969
rect 14369 32929 14381 32963
rect 14415 32960 14427 32963
rect 16482 32960 16488 32972
rect 14415 32932 16488 32960
rect 14415 32929 14427 32932
rect 14369 32923 14427 32929
rect 16482 32920 16488 32932
rect 16540 32920 16546 32972
rect 24302 32920 24308 32972
rect 24360 32960 24366 32972
rect 24397 32963 24455 32969
rect 24397 32960 24409 32963
rect 24360 32932 24409 32960
rect 24360 32920 24366 32932
rect 24397 32929 24409 32932
rect 24443 32929 24455 32963
rect 24397 32923 24455 32929
rect 24673 32963 24731 32969
rect 24673 32929 24685 32963
rect 24719 32960 24731 32963
rect 24946 32960 24952 32972
rect 24719 32932 24952 32960
rect 24719 32929 24731 32932
rect 24673 32923 24731 32929
rect 24946 32920 24952 32932
rect 25004 32920 25010 32972
rect 32306 32960 32312 32972
rect 32267 32932 32312 32960
rect 32306 32920 32312 32932
rect 32364 32920 32370 32972
rect 32585 32963 32643 32969
rect 32585 32929 32597 32963
rect 32631 32960 32643 32963
rect 33962 32960 33968 32972
rect 32631 32932 33968 32960
rect 32631 32929 32643 32932
rect 32585 32923 32643 32929
rect 33962 32920 33968 32932
rect 34020 32920 34026 32972
rect 7009 32895 7067 32901
rect 7009 32892 7021 32895
rect 6696 32864 7021 32892
rect 6696 32852 6702 32864
rect 7009 32861 7021 32864
rect 7055 32861 7067 32895
rect 7009 32855 7067 32861
rect 7101 32895 7159 32901
rect 7101 32861 7113 32895
rect 7147 32861 7159 32895
rect 7101 32855 7159 32861
rect 7193 32895 7251 32901
rect 7193 32861 7205 32895
rect 7239 32861 7251 32895
rect 7374 32892 7380 32904
rect 7335 32864 7380 32892
rect 7193 32855 7251 32861
rect 7116 32824 7144 32855
rect 7374 32852 7380 32864
rect 7432 32852 7438 32904
rect 8018 32892 8024 32904
rect 7979 32864 8024 32892
rect 8018 32852 8024 32864
rect 8076 32852 8082 32904
rect 9306 32852 9312 32904
rect 9364 32892 9370 32904
rect 10321 32895 10379 32901
rect 9364 32864 10180 32892
rect 9364 32852 9370 32864
rect 10152 32836 10180 32864
rect 10321 32861 10333 32895
rect 10367 32892 10379 32895
rect 11054 32892 11060 32904
rect 10367 32864 11060 32892
rect 10367 32861 10379 32864
rect 10321 32855 10379 32861
rect 11054 32852 11060 32864
rect 11112 32852 11118 32904
rect 13173 32895 13231 32901
rect 13173 32892 13185 32895
rect 12406 32864 13185 32892
rect 7558 32824 7564 32836
rect 7116 32796 7564 32824
rect 7558 32784 7564 32796
rect 7616 32784 7622 32836
rect 7742 32784 7748 32836
rect 7800 32824 7806 32836
rect 8205 32827 8263 32833
rect 8205 32824 8217 32827
rect 7800 32796 8217 32824
rect 7800 32784 7806 32796
rect 8205 32793 8217 32796
rect 8251 32793 8263 32827
rect 8205 32787 8263 32793
rect 9493 32827 9551 32833
rect 9493 32793 9505 32827
rect 9539 32824 9551 32827
rect 9766 32824 9772 32836
rect 9539 32796 9772 32824
rect 9539 32793 9551 32796
rect 9493 32787 9551 32793
rect 9766 32784 9772 32796
rect 9824 32784 9830 32836
rect 10134 32824 10140 32836
rect 10095 32796 10140 32824
rect 10134 32784 10140 32796
rect 10192 32784 10198 32836
rect 10686 32784 10692 32836
rect 10744 32824 10750 32836
rect 12406 32824 12434 32864
rect 13173 32861 13185 32864
rect 13219 32892 13231 32895
rect 14093 32895 14151 32901
rect 14093 32892 14105 32895
rect 13219 32864 14105 32892
rect 13219 32861 13231 32864
rect 13173 32855 13231 32861
rect 14093 32861 14105 32864
rect 14139 32861 14151 32895
rect 14093 32855 14151 32861
rect 16114 32852 16120 32904
rect 16172 32892 16178 32904
rect 16209 32895 16267 32901
rect 16209 32892 16221 32895
rect 16172 32864 16221 32892
rect 16172 32852 16178 32864
rect 16209 32861 16221 32864
rect 16255 32861 16267 32895
rect 16209 32855 16267 32861
rect 16298 32852 16304 32904
rect 16356 32892 16362 32904
rect 16715 32895 16773 32901
rect 16356 32864 16401 32892
rect 16356 32852 16362 32864
rect 16715 32861 16727 32895
rect 16761 32892 16773 32895
rect 16942 32892 16948 32904
rect 16761 32864 16948 32892
rect 16761 32861 16773 32864
rect 16715 32855 16773 32861
rect 16942 32852 16948 32864
rect 17000 32852 17006 32904
rect 17678 32892 17684 32904
rect 17639 32864 17684 32892
rect 17678 32852 17684 32864
rect 17736 32852 17742 32904
rect 17770 32852 17776 32904
rect 17828 32892 17834 32904
rect 18233 32895 18291 32901
rect 18233 32892 18245 32895
rect 17828 32864 18245 32892
rect 17828 32852 17834 32864
rect 18233 32861 18245 32864
rect 18279 32861 18291 32895
rect 23474 32892 23480 32904
rect 23435 32864 23480 32892
rect 18233 32855 18291 32861
rect 23474 32852 23480 32864
rect 23532 32852 23538 32904
rect 26878 32852 26884 32904
rect 26936 32901 26942 32904
rect 26936 32892 26948 32901
rect 26936 32864 26981 32892
rect 26936 32855 26948 32864
rect 26936 32852 26942 32855
rect 27062 32852 27068 32904
rect 27120 32892 27126 32904
rect 27157 32895 27215 32901
rect 27157 32892 27169 32895
rect 27120 32864 27169 32892
rect 27120 32852 27126 32864
rect 27157 32861 27169 32864
rect 27203 32892 27215 32895
rect 27246 32892 27252 32904
rect 27203 32864 27252 32892
rect 27203 32861 27215 32864
rect 27157 32855 27215 32861
rect 27246 32852 27252 32864
rect 27304 32852 27310 32904
rect 29914 32892 29920 32904
rect 29748 32864 29920 32892
rect 10744 32796 12434 32824
rect 10744 32784 10750 32796
rect 12986 32784 12992 32836
rect 13044 32824 13050 32836
rect 13357 32827 13415 32833
rect 13357 32824 13369 32827
rect 13044 32796 13369 32824
rect 13044 32784 13050 32796
rect 13357 32793 13369 32796
rect 13403 32824 13415 32827
rect 13538 32824 13544 32836
rect 13403 32796 13544 32824
rect 13403 32793 13415 32796
rect 13357 32787 13415 32793
rect 13538 32784 13544 32796
rect 13596 32784 13602 32836
rect 16022 32784 16028 32836
rect 16080 32824 16086 32836
rect 16485 32827 16543 32833
rect 16485 32824 16497 32827
rect 16080 32796 16497 32824
rect 16080 32784 16086 32796
rect 16485 32793 16497 32796
rect 16531 32793 16543 32827
rect 16485 32787 16543 32793
rect 16577 32827 16635 32833
rect 16577 32793 16589 32827
rect 16623 32824 16635 32827
rect 18414 32824 18420 32836
rect 16623 32796 18420 32824
rect 16623 32793 16635 32796
rect 16577 32787 16635 32793
rect 18414 32784 18420 32796
rect 18472 32784 18478 32836
rect 18601 32827 18659 32833
rect 18601 32793 18613 32827
rect 18647 32824 18659 32827
rect 18690 32824 18696 32836
rect 18647 32796 18696 32824
rect 18647 32793 18659 32796
rect 18601 32787 18659 32793
rect 18690 32784 18696 32796
rect 18748 32784 18754 32836
rect 19978 32784 19984 32836
rect 20036 32824 20042 32836
rect 21358 32824 21364 32836
rect 20036 32796 21364 32824
rect 20036 32784 20042 32796
rect 21358 32784 21364 32796
rect 21416 32784 21422 32836
rect 23658 32784 23664 32836
rect 23716 32824 23722 32836
rect 24210 32824 24216 32836
rect 23716 32796 24216 32824
rect 23716 32784 23722 32796
rect 24210 32784 24216 32796
rect 24268 32784 24274 32836
rect 29748 32768 29776 32864
rect 29914 32852 29920 32864
rect 29972 32892 29978 32904
rect 30285 32895 30343 32901
rect 30285 32892 30297 32895
rect 29972 32864 30297 32892
rect 29972 32852 29978 32864
rect 30285 32861 30297 32864
rect 30331 32861 30343 32895
rect 30285 32855 30343 32861
rect 31481 32895 31539 32901
rect 31481 32861 31493 32895
rect 31527 32892 31539 32895
rect 31754 32892 31760 32904
rect 31527 32864 31760 32892
rect 31527 32861 31539 32864
rect 31481 32855 31539 32861
rect 31754 32852 31760 32864
rect 31812 32892 31818 32904
rect 32122 32892 32128 32904
rect 31812 32864 32128 32892
rect 31812 32852 31818 32864
rect 32122 32852 32128 32864
rect 32180 32852 32186 32904
rect 35802 32852 35808 32904
rect 35860 32901 35866 32904
rect 35860 32892 35872 32901
rect 36078 32892 36084 32904
rect 35860 32864 35905 32892
rect 35991 32864 36084 32892
rect 35860 32855 35872 32864
rect 35860 32852 35866 32855
rect 36078 32852 36084 32864
rect 36136 32892 36142 32904
rect 38930 32892 38936 32904
rect 36136 32864 38936 32892
rect 36136 32852 36142 32864
rect 38930 32852 38936 32864
rect 38988 32852 38994 32904
rect 31665 32827 31723 32833
rect 31665 32793 31677 32827
rect 31711 32824 31723 32827
rect 34146 32824 34152 32836
rect 31711 32796 34152 32824
rect 31711 32793 31723 32796
rect 31665 32787 31723 32793
rect 34146 32784 34152 32796
rect 34204 32784 34210 32836
rect 6181 32759 6239 32765
rect 6181 32756 6193 32759
rect 5776 32728 6193 32756
rect 5776 32716 5782 32728
rect 6181 32725 6193 32728
rect 6227 32725 6239 32759
rect 6181 32719 6239 32725
rect 10505 32759 10563 32765
rect 10505 32725 10517 32759
rect 10551 32756 10563 32759
rect 10778 32756 10784 32768
rect 10551 32728 10784 32756
rect 10551 32725 10563 32728
rect 10505 32719 10563 32725
rect 10778 32716 10784 32728
rect 10836 32716 10842 32768
rect 10962 32716 10968 32768
rect 11020 32756 11026 32768
rect 11057 32759 11115 32765
rect 11057 32756 11069 32759
rect 11020 32728 11069 32756
rect 11020 32716 11026 32728
rect 11057 32725 11069 32728
rect 11103 32725 11115 32759
rect 11057 32719 11115 32725
rect 15010 32716 15016 32768
rect 15068 32756 15074 32768
rect 15473 32759 15531 32765
rect 15473 32756 15485 32759
rect 15068 32728 15485 32756
rect 15068 32716 15074 32728
rect 15473 32725 15485 32728
rect 15519 32756 15531 32759
rect 16114 32756 16120 32768
rect 15519 32728 16120 32756
rect 15519 32725 15531 32728
rect 15473 32719 15531 32725
rect 16114 32716 16120 32728
rect 16172 32716 16178 32768
rect 16853 32759 16911 32765
rect 16853 32725 16865 32759
rect 16899 32756 16911 32759
rect 17586 32756 17592 32768
rect 16899 32728 17592 32756
rect 16899 32725 16911 32728
rect 16853 32719 16911 32725
rect 17586 32716 17592 32728
rect 17644 32716 17650 32768
rect 22094 32716 22100 32768
rect 22152 32756 22158 32768
rect 22152 32728 22197 32756
rect 22152 32716 22158 32728
rect 25038 32716 25044 32768
rect 25096 32756 25102 32768
rect 25777 32759 25835 32765
rect 25777 32756 25789 32759
rect 25096 32728 25789 32756
rect 25096 32716 25102 32728
rect 25777 32725 25789 32728
rect 25823 32725 25835 32759
rect 29730 32756 29736 32768
rect 29691 32728 29736 32756
rect 25777 32719 25835 32725
rect 29730 32716 29736 32728
rect 29788 32716 29794 32768
rect 30374 32716 30380 32768
rect 30432 32756 30438 32768
rect 30469 32759 30527 32765
rect 30469 32756 30481 32759
rect 30432 32728 30481 32756
rect 30432 32716 30438 32728
rect 30469 32725 30481 32728
rect 30515 32725 30527 32759
rect 30469 32719 30527 32725
rect 31849 32759 31907 32765
rect 31849 32725 31861 32759
rect 31895 32756 31907 32759
rect 32398 32756 32404 32768
rect 31895 32728 32404 32756
rect 31895 32725 31907 32728
rect 31849 32719 31907 32725
rect 32398 32716 32404 32728
rect 32456 32716 32462 32768
rect 34606 32716 34612 32768
rect 34664 32756 34670 32768
rect 34701 32759 34759 32765
rect 34701 32756 34713 32759
rect 34664 32728 34713 32756
rect 34664 32716 34670 32728
rect 34701 32725 34713 32728
rect 34747 32725 34759 32759
rect 34701 32719 34759 32725
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 5169 32555 5227 32561
rect 5169 32521 5181 32555
rect 5215 32552 5227 32555
rect 5442 32552 5448 32564
rect 5215 32524 5448 32552
rect 5215 32521 5227 32524
rect 5169 32515 5227 32521
rect 5442 32512 5448 32524
rect 5500 32512 5506 32564
rect 5534 32512 5540 32564
rect 5592 32552 5598 32564
rect 5629 32555 5687 32561
rect 5629 32552 5641 32555
rect 5592 32524 5641 32552
rect 5592 32512 5598 32524
rect 5629 32521 5641 32524
rect 5675 32552 5687 32555
rect 5675 32524 6684 32552
rect 5675 32521 5687 32524
rect 5629 32515 5687 32521
rect 6656 32493 6684 32524
rect 12802 32512 12808 32564
rect 12860 32552 12866 32564
rect 13998 32552 14004 32564
rect 12860 32524 14004 32552
rect 12860 32512 12866 32524
rect 13998 32512 14004 32524
rect 14056 32552 14062 32564
rect 14734 32552 14740 32564
rect 14056 32524 14740 32552
rect 14056 32512 14062 32524
rect 14734 32512 14740 32524
rect 14792 32512 14798 32564
rect 17678 32512 17684 32564
rect 17736 32552 17742 32564
rect 17954 32552 17960 32564
rect 17736 32524 17960 32552
rect 17736 32512 17742 32524
rect 17954 32512 17960 32524
rect 18012 32512 18018 32564
rect 18414 32512 18420 32564
rect 18472 32552 18478 32564
rect 20073 32555 20131 32561
rect 20073 32552 20085 32555
rect 18472 32524 20085 32552
rect 18472 32512 18478 32524
rect 20073 32521 20085 32524
rect 20119 32521 20131 32555
rect 20073 32515 20131 32521
rect 24302 32512 24308 32564
rect 24360 32552 24366 32564
rect 25317 32555 25375 32561
rect 25317 32552 25329 32555
rect 24360 32524 25329 32552
rect 24360 32512 24366 32524
rect 25317 32521 25329 32524
rect 25363 32521 25375 32555
rect 29546 32552 29552 32564
rect 25317 32515 25375 32521
rect 28276 32524 29552 32552
rect 6641 32487 6699 32493
rect 6641 32453 6653 32487
rect 6687 32453 6699 32487
rect 6641 32447 6699 32453
rect 9398 32444 9404 32496
rect 9456 32484 9462 32496
rect 9950 32484 9956 32496
rect 9456 32456 9956 32484
rect 9456 32444 9462 32456
rect 9950 32444 9956 32456
rect 10008 32484 10014 32496
rect 18233 32487 18291 32493
rect 10008 32456 10732 32484
rect 10008 32444 10014 32456
rect 2130 32376 2136 32428
rect 2188 32416 2194 32428
rect 2481 32419 2539 32425
rect 2481 32416 2493 32419
rect 2188 32388 2493 32416
rect 2188 32376 2194 32388
rect 2481 32385 2493 32388
rect 2527 32385 2539 32419
rect 2481 32379 2539 32385
rect 5813 32419 5871 32425
rect 5813 32385 5825 32419
rect 5859 32385 5871 32419
rect 5813 32379 5871 32385
rect 6825 32419 6883 32425
rect 6825 32385 6837 32419
rect 6871 32416 6883 32419
rect 7098 32416 7104 32428
rect 6871 32388 7104 32416
rect 6871 32385 6883 32388
rect 6825 32379 6883 32385
rect 1854 32308 1860 32360
rect 1912 32348 1918 32360
rect 2225 32351 2283 32357
rect 2225 32348 2237 32351
rect 1912 32320 2237 32348
rect 1912 32308 1918 32320
rect 2225 32317 2237 32320
rect 2271 32317 2283 32351
rect 2225 32311 2283 32317
rect 5828 32280 5856 32379
rect 7098 32376 7104 32388
rect 7156 32376 7162 32428
rect 7742 32376 7748 32428
rect 7800 32416 7806 32428
rect 10704 32425 10732 32456
rect 17604 32456 18184 32484
rect 9585 32419 9643 32425
rect 10597 32419 10655 32425
rect 9585 32416 9597 32419
rect 7800 32388 9597 32416
rect 7800 32376 7806 32388
rect 9585 32385 9597 32388
rect 9631 32385 9643 32419
rect 9585 32379 9643 32385
rect 10520 32391 10609 32419
rect 6546 32308 6552 32360
rect 6604 32348 6610 32360
rect 8297 32351 8355 32357
rect 8297 32348 8309 32351
rect 6604 32320 8309 32348
rect 6604 32308 6610 32320
rect 8297 32317 8309 32320
rect 8343 32317 8355 32351
rect 8570 32348 8576 32360
rect 8531 32320 8576 32348
rect 8297 32311 8355 32317
rect 8570 32308 8576 32320
rect 8628 32308 8634 32360
rect 9861 32351 9919 32357
rect 9861 32317 9873 32351
rect 9907 32348 9919 32351
rect 10410 32348 10416 32360
rect 9907 32320 10416 32348
rect 9907 32317 9919 32320
rect 9861 32311 9919 32317
rect 10410 32308 10416 32320
rect 10468 32308 10474 32360
rect 10520 32348 10548 32391
rect 10597 32385 10609 32391
rect 10643 32385 10655 32419
rect 10597 32379 10655 32385
rect 10689 32419 10747 32425
rect 10689 32385 10701 32419
rect 10735 32385 10747 32419
rect 10689 32379 10747 32385
rect 10778 32376 10784 32428
rect 10836 32416 10842 32428
rect 10836 32388 10881 32416
rect 10836 32376 10842 32388
rect 10962 32376 10968 32428
rect 11020 32416 11026 32428
rect 11609 32419 11667 32425
rect 11020 32388 11065 32416
rect 11020 32376 11026 32388
rect 11609 32385 11621 32419
rect 11655 32416 11667 32419
rect 14918 32416 14924 32428
rect 11655 32388 14924 32416
rect 11655 32385 11667 32388
rect 11609 32379 11667 32385
rect 11624 32348 11652 32379
rect 14918 32376 14924 32388
rect 14976 32376 14982 32428
rect 15010 32376 15016 32428
rect 15068 32416 15074 32428
rect 17604 32425 17632 32456
rect 17589 32419 17647 32425
rect 17589 32416 17601 32419
rect 15068 32388 17601 32416
rect 15068 32376 15074 32388
rect 17589 32385 17601 32388
rect 17635 32385 17647 32419
rect 17770 32416 17776 32428
rect 17731 32388 17776 32416
rect 17589 32379 17647 32385
rect 17770 32376 17776 32388
rect 17828 32376 17834 32428
rect 17865 32419 17923 32425
rect 17865 32385 17877 32419
rect 17911 32385 17923 32419
rect 17865 32379 17923 32385
rect 10520 32320 11652 32348
rect 15378 32308 15384 32360
rect 15436 32348 15442 32360
rect 17678 32348 17684 32360
rect 15436 32320 17684 32348
rect 15436 32308 15442 32320
rect 17678 32308 17684 32320
rect 17736 32308 17742 32360
rect 17880 32280 17908 32379
rect 17954 32376 17960 32428
rect 18012 32416 18018 32428
rect 18156 32416 18184 32456
rect 18233 32453 18245 32487
rect 18279 32484 18291 32487
rect 18938 32487 18996 32493
rect 18938 32484 18950 32487
rect 18279 32456 18950 32484
rect 18279 32453 18291 32456
rect 18233 32447 18291 32453
rect 18938 32453 18950 32456
rect 18984 32453 18996 32487
rect 18938 32447 18996 32453
rect 20530 32444 20536 32496
rect 20588 32484 20594 32496
rect 28276 32484 28304 32524
rect 29546 32512 29552 32524
rect 29604 32512 29610 32564
rect 30561 32555 30619 32561
rect 30561 32521 30573 32555
rect 30607 32552 30619 32555
rect 31202 32552 31208 32564
rect 30607 32524 31208 32552
rect 30607 32521 30619 32524
rect 30561 32515 30619 32521
rect 31202 32512 31208 32524
rect 31260 32512 31266 32564
rect 32861 32555 32919 32561
rect 32861 32521 32873 32555
rect 32907 32552 32919 32555
rect 32950 32552 32956 32564
rect 32907 32524 32956 32552
rect 32907 32521 32919 32524
rect 32861 32515 32919 32521
rect 32950 32512 32956 32524
rect 33008 32512 33014 32564
rect 28442 32484 28448 32496
rect 20588 32456 28304 32484
rect 28403 32456 28448 32484
rect 20588 32444 20594 32456
rect 28442 32444 28448 32456
rect 28500 32444 28506 32496
rect 32306 32444 32312 32496
rect 32364 32484 32370 32496
rect 32364 32456 32536 32484
rect 32364 32444 32370 32456
rect 18322 32416 18328 32428
rect 18012 32388 18057 32416
rect 18156 32388 18328 32416
rect 18012 32376 18018 32388
rect 18322 32376 18328 32388
rect 18380 32376 18386 32428
rect 22094 32376 22100 32428
rect 22152 32416 22158 32428
rect 22189 32419 22247 32425
rect 22189 32416 22201 32419
rect 22152 32388 22201 32416
rect 22152 32376 22158 32388
rect 22189 32385 22201 32388
rect 22235 32416 22247 32419
rect 24026 32416 24032 32428
rect 22235 32388 24032 32416
rect 22235 32385 22247 32388
rect 22189 32379 22247 32385
rect 24026 32376 24032 32388
rect 24084 32376 24090 32428
rect 24302 32416 24308 32428
rect 24263 32388 24308 32416
rect 24302 32376 24308 32388
rect 24360 32376 24366 32428
rect 28353 32419 28411 32425
rect 28353 32385 28365 32419
rect 28399 32385 28411 32419
rect 28534 32416 28540 32428
rect 28495 32388 28540 32416
rect 28353 32379 28411 32385
rect 18693 32351 18751 32357
rect 18693 32317 18705 32351
rect 18739 32317 18751 32351
rect 18693 32311 18751 32317
rect 17954 32280 17960 32292
rect 5828 32252 12434 32280
rect 17880 32252 17960 32280
rect 3602 32212 3608 32224
rect 3563 32184 3608 32212
rect 3602 32172 3608 32184
rect 3660 32172 3666 32224
rect 6822 32172 6828 32224
rect 6880 32212 6886 32224
rect 7009 32215 7067 32221
rect 7009 32212 7021 32215
rect 6880 32184 7021 32212
rect 6880 32172 6886 32184
rect 7009 32181 7021 32184
rect 7055 32181 7067 32215
rect 10318 32212 10324 32224
rect 10279 32184 10324 32212
rect 7009 32175 7067 32181
rect 10318 32172 10324 32184
rect 10376 32172 10382 32224
rect 10410 32172 10416 32224
rect 10468 32212 10474 32224
rect 10686 32212 10692 32224
rect 10468 32184 10692 32212
rect 10468 32172 10474 32184
rect 10686 32172 10692 32184
rect 10744 32212 10750 32224
rect 10962 32212 10968 32224
rect 10744 32184 10968 32212
rect 10744 32172 10750 32184
rect 10962 32172 10968 32184
rect 11020 32172 11026 32224
rect 12406 32212 12434 32252
rect 17954 32240 17960 32252
rect 18012 32240 18018 32292
rect 13814 32212 13820 32224
rect 12406 32184 13820 32212
rect 13814 32172 13820 32184
rect 13872 32172 13878 32224
rect 17862 32172 17868 32224
rect 17920 32212 17926 32224
rect 18708 32212 18736 32311
rect 28166 32308 28172 32360
rect 28224 32348 28230 32360
rect 28368 32348 28396 32379
rect 28534 32376 28540 32388
rect 28592 32376 28598 32428
rect 28718 32416 28724 32428
rect 28679 32388 28724 32416
rect 28718 32376 28724 32388
rect 28776 32376 28782 32428
rect 30377 32419 30435 32425
rect 30377 32385 30389 32419
rect 30423 32416 30435 32419
rect 30834 32416 30840 32428
rect 30423 32388 30840 32416
rect 30423 32385 30435 32388
rect 30377 32379 30435 32385
rect 30834 32376 30840 32388
rect 30892 32376 30898 32428
rect 32217 32419 32275 32425
rect 32217 32385 32229 32419
rect 32263 32385 32275 32419
rect 32398 32416 32404 32428
rect 32359 32388 32404 32416
rect 32217 32379 32275 32385
rect 29362 32348 29368 32360
rect 28224 32320 29368 32348
rect 28224 32308 28230 32320
rect 29362 32308 29368 32320
rect 29420 32308 29426 32360
rect 32232 32348 32260 32379
rect 32398 32376 32404 32388
rect 32456 32376 32462 32428
rect 32508 32425 32536 32456
rect 32493 32419 32551 32425
rect 32493 32385 32505 32419
rect 32539 32385 32551 32419
rect 32493 32379 32551 32385
rect 32582 32376 32588 32428
rect 32640 32416 32646 32428
rect 32640 32388 32685 32416
rect 32640 32376 32646 32388
rect 36630 32376 36636 32428
rect 36688 32416 36694 32428
rect 38390 32419 38448 32425
rect 38390 32416 38402 32419
rect 36688 32388 38402 32416
rect 36688 32376 36694 32388
rect 38390 32385 38402 32388
rect 38436 32385 38448 32419
rect 38390 32379 38448 32385
rect 33502 32348 33508 32360
rect 32232 32320 33508 32348
rect 33502 32308 33508 32320
rect 33560 32308 33566 32360
rect 38657 32351 38715 32357
rect 38657 32317 38669 32351
rect 38703 32348 38715 32351
rect 38930 32348 38936 32360
rect 38703 32320 38936 32348
rect 38703 32317 38715 32320
rect 38657 32311 38715 32317
rect 38930 32308 38936 32320
rect 38988 32308 38994 32360
rect 23474 32240 23480 32292
rect 23532 32280 23538 32292
rect 24489 32283 24547 32289
rect 24489 32280 24501 32283
rect 23532 32252 24501 32280
rect 23532 32240 23538 32252
rect 24489 32249 24501 32252
rect 24535 32249 24547 32283
rect 24489 32243 24547 32249
rect 28718 32240 28724 32292
rect 28776 32280 28782 32292
rect 29638 32280 29644 32292
rect 28776 32252 29644 32280
rect 28776 32240 28782 32252
rect 29638 32240 29644 32252
rect 29696 32240 29702 32292
rect 17920 32184 18736 32212
rect 22373 32215 22431 32221
rect 17920 32172 17926 32184
rect 22373 32181 22385 32215
rect 22419 32212 22431 32215
rect 23750 32212 23756 32224
rect 22419 32184 23756 32212
rect 22419 32181 22431 32184
rect 22373 32175 22431 32181
rect 23750 32172 23756 32184
rect 23808 32212 23814 32224
rect 24394 32212 24400 32224
rect 23808 32184 24400 32212
rect 23808 32172 23814 32184
rect 24394 32172 24400 32184
rect 24452 32172 24458 32224
rect 26694 32172 26700 32224
rect 26752 32212 26758 32224
rect 28169 32215 28227 32221
rect 28169 32212 28181 32215
rect 26752 32184 28181 32212
rect 26752 32172 26758 32184
rect 28169 32181 28181 32184
rect 28215 32181 28227 32215
rect 37274 32212 37280 32224
rect 37235 32184 37280 32212
rect 28169 32175 28227 32181
rect 37274 32172 37280 32184
rect 37332 32172 37338 32224
rect 58158 32212 58164 32224
rect 58119 32184 58164 32212
rect 58158 32172 58164 32184
rect 58216 32172 58222 32224
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 2130 32008 2136 32020
rect 2091 31980 2136 32008
rect 2130 31968 2136 31980
rect 2188 31968 2194 32020
rect 6178 32008 6184 32020
rect 5276 31980 6184 32008
rect 5276 31952 5304 31980
rect 6178 31968 6184 31980
rect 6236 31968 6242 32020
rect 7006 31968 7012 32020
rect 7064 32008 7070 32020
rect 7193 32011 7251 32017
rect 7193 32008 7205 32011
rect 7064 31980 7205 32008
rect 7064 31968 7070 31980
rect 7193 31977 7205 31980
rect 7239 32008 7251 32011
rect 8202 32008 8208 32020
rect 7239 31980 8208 32008
rect 7239 31977 7251 31980
rect 7193 31971 7251 31977
rect 8202 31968 8208 31980
rect 8260 31968 8266 32020
rect 10873 32011 10931 32017
rect 10873 31977 10885 32011
rect 10919 32008 10931 32011
rect 11054 32008 11060 32020
rect 10919 31980 11060 32008
rect 10919 31977 10931 31980
rect 10873 31971 10931 31977
rect 11054 31968 11060 31980
rect 11112 31968 11118 32020
rect 13357 32011 13415 32017
rect 13357 31977 13369 32011
rect 13403 32008 13415 32011
rect 14550 32008 14556 32020
rect 13403 31980 14556 32008
rect 13403 31977 13415 31980
rect 13357 31971 13415 31977
rect 14550 31968 14556 31980
rect 14608 31968 14614 32020
rect 23750 31968 23756 32020
rect 23808 32008 23814 32020
rect 24118 32008 24124 32020
rect 23808 31980 24124 32008
rect 23808 31968 23814 31980
rect 24118 31968 24124 31980
rect 24176 31968 24182 32020
rect 27246 31968 27252 32020
rect 27304 32008 27310 32020
rect 27304 31980 28396 32008
rect 27304 31968 27310 31980
rect 5258 31900 5264 31952
rect 5316 31900 5322 31952
rect 5442 31900 5448 31952
rect 5500 31940 5506 31952
rect 8113 31943 8171 31949
rect 5500 31912 5580 31940
rect 5500 31900 5506 31912
rect 5276 31872 5304 31900
rect 5092 31844 5304 31872
rect 2314 31764 2320 31816
rect 2372 31813 2378 31816
rect 2372 31807 2421 31813
rect 2372 31773 2375 31807
rect 2409 31773 2421 31807
rect 2372 31767 2421 31773
rect 2482 31804 2540 31810
rect 2482 31770 2494 31804
rect 2528 31770 2540 31804
rect 2372 31764 2378 31767
rect 2482 31764 2540 31770
rect 2590 31764 2596 31816
rect 2648 31804 2654 31816
rect 2648 31776 2693 31804
rect 2648 31764 2654 31776
rect 2774 31764 2780 31816
rect 2832 31804 2838 31816
rect 4982 31804 4988 31816
rect 2832 31776 4988 31804
rect 2832 31764 2838 31776
rect 4982 31764 4988 31776
rect 5040 31764 5046 31816
rect 5092 31813 5120 31844
rect 5077 31807 5135 31813
rect 5077 31773 5089 31807
rect 5123 31773 5135 31807
rect 5077 31767 5135 31773
rect 5169 31807 5227 31813
rect 5169 31773 5181 31807
rect 5215 31773 5227 31807
rect 5169 31767 5227 31773
rect 2497 31736 2525 31764
rect 2682 31736 2688 31748
rect 2497 31708 2688 31736
rect 2682 31696 2688 31708
rect 2740 31696 2746 31748
rect 4890 31696 4896 31748
rect 4948 31736 4954 31748
rect 5184 31736 5212 31767
rect 5258 31764 5264 31816
rect 5316 31804 5322 31816
rect 5445 31807 5503 31813
rect 5316 31776 5361 31804
rect 5316 31764 5322 31776
rect 5445 31773 5457 31807
rect 5491 31804 5503 31807
rect 5552 31804 5580 31912
rect 8113 31909 8125 31943
rect 8159 31940 8171 31943
rect 8294 31940 8300 31952
rect 8159 31912 8300 31940
rect 8159 31909 8171 31912
rect 8113 31903 8171 31909
rect 5905 31807 5963 31813
rect 5491 31776 5593 31804
rect 5491 31773 5503 31776
rect 5445 31767 5503 31773
rect 5905 31773 5917 31807
rect 5951 31804 5963 31807
rect 8128 31804 8156 31903
rect 8294 31900 8300 31912
rect 8352 31900 8358 31952
rect 11330 31900 11336 31952
rect 11388 31940 11394 31952
rect 17218 31940 17224 31952
rect 11388 31912 17224 31940
rect 11388 31900 11394 31912
rect 17218 31900 17224 31912
rect 17276 31900 17282 31952
rect 27890 31900 27896 31952
rect 27948 31940 27954 31952
rect 28077 31943 28135 31949
rect 28077 31940 28089 31943
rect 27948 31912 28089 31940
rect 27948 31900 27954 31912
rect 28077 31909 28089 31912
rect 28123 31909 28135 31943
rect 28077 31903 28135 31909
rect 8202 31832 8208 31884
rect 8260 31872 8266 31884
rect 9493 31875 9551 31881
rect 9493 31872 9505 31875
rect 8260 31844 9505 31872
rect 8260 31832 8266 31844
rect 9493 31841 9505 31844
rect 9539 31841 9551 31875
rect 9493 31835 9551 31841
rect 12894 31832 12900 31884
rect 12952 31872 12958 31884
rect 12952 31844 13032 31872
rect 12952 31832 12958 31844
rect 5951 31776 8156 31804
rect 9760 31807 9818 31813
rect 5951 31773 5963 31776
rect 5905 31767 5963 31773
rect 9760 31773 9772 31807
rect 9806 31804 9818 31807
rect 10318 31804 10324 31816
rect 9806 31776 10324 31804
rect 9806 31773 9818 31776
rect 9760 31767 9818 31773
rect 4948 31708 5212 31736
rect 5460 31736 5488 31767
rect 10318 31764 10324 31776
rect 10376 31764 10382 31816
rect 13004 31813 13032 31844
rect 13446 31832 13452 31884
rect 13504 31872 13510 31884
rect 16301 31875 16359 31881
rect 13504 31844 14504 31872
rect 13504 31832 13510 31844
rect 14476 31813 14504 31844
rect 16301 31841 16313 31875
rect 16347 31872 16359 31875
rect 17954 31872 17960 31884
rect 16347 31844 17960 31872
rect 16347 31841 16359 31844
rect 16301 31835 16359 31841
rect 17954 31832 17960 31844
rect 18012 31832 18018 31884
rect 22833 31875 22891 31881
rect 22833 31872 22845 31875
rect 22066 31844 22845 31872
rect 12989 31807 13047 31813
rect 12989 31773 13001 31807
rect 13035 31773 13047 31807
rect 12989 31767 13047 31773
rect 14349 31807 14407 31813
rect 14349 31773 14361 31807
rect 14395 31804 14407 31807
rect 14458 31807 14516 31813
rect 14395 31773 14412 31804
rect 14349 31767 14412 31773
rect 14458 31773 14470 31807
rect 14504 31773 14516 31807
rect 14458 31767 14516 31773
rect 7374 31736 7380 31748
rect 5460 31708 7380 31736
rect 4948 31696 4954 31708
rect 4798 31668 4804 31680
rect 4759 31640 4804 31668
rect 4798 31628 4804 31640
rect 4856 31628 4862 31680
rect 5184 31668 5212 31708
rect 7374 31696 7380 31708
rect 7432 31696 7438 31748
rect 13078 31696 13084 31748
rect 13136 31736 13142 31748
rect 13173 31739 13231 31745
rect 13173 31736 13185 31739
rect 13136 31708 13185 31736
rect 13136 31696 13142 31708
rect 13173 31705 13185 31708
rect 13219 31705 13231 31739
rect 14384 31736 14412 31767
rect 14550 31764 14556 31816
rect 14608 31801 14614 31816
rect 14734 31804 14740 31816
rect 14608 31773 14650 31801
rect 14695 31776 14740 31804
rect 14608 31764 14614 31773
rect 14734 31764 14740 31776
rect 14792 31764 14798 31816
rect 16761 31807 16819 31813
rect 16761 31773 16773 31807
rect 16807 31804 16819 31807
rect 16850 31804 16856 31816
rect 16807 31776 16856 31804
rect 16807 31773 16819 31776
rect 16761 31767 16819 31773
rect 16850 31764 16856 31776
rect 16908 31764 16914 31816
rect 20438 31764 20444 31816
rect 20496 31804 20502 31816
rect 21453 31807 21511 31813
rect 21453 31804 21465 31807
rect 20496 31776 21465 31804
rect 20496 31764 20502 31776
rect 21453 31773 21465 31776
rect 21499 31804 21511 31807
rect 22066 31804 22094 31844
rect 22833 31841 22845 31844
rect 22879 31841 22891 31875
rect 22833 31835 22891 31841
rect 24670 31832 24676 31884
rect 24728 31872 24734 31884
rect 25041 31875 25099 31881
rect 25041 31872 25053 31875
rect 24728 31844 25053 31872
rect 24728 31832 24734 31844
rect 25041 31841 25053 31844
rect 25087 31841 25099 31875
rect 28368 31872 28396 31980
rect 28442 31968 28448 32020
rect 28500 32008 28506 32020
rect 30742 32008 30748 32020
rect 28500 31980 30748 32008
rect 28500 31968 28506 31980
rect 30742 31968 30748 31980
rect 30800 31968 30806 32020
rect 30929 32011 30987 32017
rect 30929 31977 30941 32011
rect 30975 32008 30987 32011
rect 31018 32008 31024 32020
rect 30975 31980 31024 32008
rect 30975 31977 30987 31980
rect 30929 31971 30987 31977
rect 31018 31968 31024 31980
rect 31076 32008 31082 32020
rect 31386 32008 31392 32020
rect 31076 31980 31392 32008
rect 31076 31968 31082 31980
rect 31386 31968 31392 31980
rect 31444 31968 31450 32020
rect 32125 32011 32183 32017
rect 32125 31977 32137 32011
rect 32171 32008 32183 32011
rect 32582 32008 32588 32020
rect 32171 31980 32588 32008
rect 32171 31977 32183 31980
rect 32125 31971 32183 31977
rect 32582 31968 32588 31980
rect 32640 31968 32646 32020
rect 36630 32008 36636 32020
rect 36591 31980 36636 32008
rect 36630 31968 36636 31980
rect 36688 31968 36694 32020
rect 33410 31900 33416 31952
rect 33468 31940 33474 31952
rect 35437 31943 35495 31949
rect 35437 31940 35449 31943
rect 33468 31912 35449 31940
rect 33468 31900 33474 31912
rect 35437 31909 35449 31912
rect 35483 31940 35495 31943
rect 35483 31912 36492 31940
rect 35483 31909 35495 31912
rect 35437 31903 35495 31909
rect 29549 31875 29607 31881
rect 29549 31872 29561 31875
rect 28368 31844 29561 31872
rect 25041 31835 25099 31841
rect 29549 31841 29561 31844
rect 29595 31841 29607 31875
rect 29549 31835 29607 31841
rect 22554 31804 22560 31816
rect 21499 31776 22094 31804
rect 22515 31776 22560 31804
rect 21499 31773 21511 31776
rect 21453 31767 21511 31773
rect 22554 31764 22560 31776
rect 22612 31764 22618 31816
rect 24765 31807 24823 31813
rect 24765 31773 24777 31807
rect 24811 31804 24823 31807
rect 24854 31804 24860 31816
rect 24811 31776 24860 31804
rect 24811 31773 24823 31776
rect 24765 31767 24823 31773
rect 24854 31764 24860 31776
rect 24912 31764 24918 31816
rect 28166 31764 28172 31816
rect 28224 31804 28230 31816
rect 28261 31807 28319 31813
rect 28261 31804 28273 31807
rect 28224 31776 28273 31804
rect 28224 31764 28230 31776
rect 28261 31773 28273 31776
rect 28307 31773 28319 31807
rect 28261 31767 28319 31773
rect 28350 31764 28356 31816
rect 28408 31804 28414 31816
rect 28626 31804 28632 31816
rect 28408 31776 28453 31804
rect 28587 31776 28632 31804
rect 28408 31764 28414 31776
rect 28626 31764 28632 31776
rect 28684 31764 28690 31816
rect 29816 31807 29874 31813
rect 29816 31773 29828 31807
rect 29862 31804 29874 31807
rect 30098 31804 30104 31816
rect 29862 31776 30104 31804
rect 29862 31773 29874 31776
rect 29816 31767 29874 31773
rect 30098 31764 30104 31776
rect 30156 31764 30162 31816
rect 30926 31764 30932 31816
rect 30984 31804 30990 31816
rect 35986 31804 35992 31816
rect 30984 31776 35992 31804
rect 30984 31764 30990 31776
rect 35986 31764 35992 31776
rect 36044 31764 36050 31816
rect 36170 31804 36176 31816
rect 36131 31776 36176 31804
rect 36170 31764 36176 31776
rect 36228 31764 36234 31816
rect 36377 31807 36435 31813
rect 36268 31801 36326 31807
rect 36268 31767 36280 31801
rect 36314 31767 36326 31801
rect 36377 31773 36389 31807
rect 36423 31804 36435 31807
rect 36464 31804 36492 31912
rect 36423 31776 36492 31804
rect 36423 31773 36435 31776
rect 36377 31767 36435 31773
rect 36268 31761 36326 31767
rect 14384 31708 15332 31736
rect 13173 31699 13231 31705
rect 6546 31668 6552 31680
rect 5184 31640 6552 31668
rect 6546 31628 6552 31640
rect 6604 31628 6610 31680
rect 14090 31668 14096 31680
rect 14051 31640 14096 31668
rect 14090 31628 14096 31640
rect 14148 31628 14154 31680
rect 15304 31677 15332 31708
rect 15562 31696 15568 31748
rect 15620 31736 15626 31748
rect 16117 31739 16175 31745
rect 16117 31736 16129 31739
rect 15620 31708 16129 31736
rect 15620 31696 15626 31708
rect 16117 31705 16129 31708
rect 16163 31705 16175 31739
rect 28442 31736 28448 31748
rect 28403 31708 28448 31736
rect 16117 31699 16175 31705
rect 28442 31696 28448 31708
rect 28500 31696 28506 31748
rect 36280 31680 36308 31761
rect 15289 31671 15347 31677
rect 15289 31637 15301 31671
rect 15335 31668 15347 31671
rect 15838 31668 15844 31680
rect 15335 31640 15844 31668
rect 15335 31637 15347 31640
rect 15289 31631 15347 31637
rect 15838 31628 15844 31640
rect 15896 31628 15902 31680
rect 17862 31628 17868 31680
rect 17920 31668 17926 31680
rect 18049 31671 18107 31677
rect 18049 31668 18061 31671
rect 17920 31640 18061 31668
rect 17920 31628 17926 31640
rect 18049 31637 18061 31640
rect 18095 31637 18107 31671
rect 26050 31668 26056 31680
rect 26011 31640 26056 31668
rect 18049 31631 18107 31637
rect 26050 31628 26056 31640
rect 26108 31628 26114 31680
rect 32398 31628 32404 31680
rect 32456 31668 32462 31680
rect 32585 31671 32643 31677
rect 32585 31668 32597 31671
rect 32456 31640 32597 31668
rect 32456 31628 32462 31640
rect 32585 31637 32597 31640
rect 32631 31637 32643 31671
rect 32585 31631 32643 31637
rect 36262 31628 36268 31680
rect 36320 31628 36326 31680
rect 37553 31671 37611 31677
rect 37553 31637 37565 31671
rect 37599 31668 37611 31671
rect 37642 31668 37648 31680
rect 37599 31640 37648 31668
rect 37599 31637 37611 31640
rect 37553 31631 37611 31637
rect 37642 31628 37648 31640
rect 37700 31628 37706 31680
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 2409 31467 2467 31473
rect 2409 31433 2421 31467
rect 2455 31464 2467 31467
rect 2590 31464 2596 31476
rect 2455 31436 2596 31464
rect 2455 31433 2467 31436
rect 2409 31427 2467 31433
rect 2590 31424 2596 31436
rect 2648 31424 2654 31476
rect 5258 31424 5264 31476
rect 5316 31464 5322 31476
rect 5445 31467 5503 31473
rect 5445 31464 5457 31467
rect 5316 31436 5457 31464
rect 5316 31424 5322 31436
rect 5445 31433 5457 31436
rect 5491 31433 5503 31467
rect 5445 31427 5503 31433
rect 8294 31424 8300 31476
rect 8352 31464 8358 31476
rect 12253 31467 12311 31473
rect 8352 31436 8397 31464
rect 8352 31424 8358 31436
rect 12253 31433 12265 31467
rect 12299 31464 12311 31467
rect 13078 31464 13084 31476
rect 12299 31436 13084 31464
rect 12299 31433 12311 31436
rect 12253 31427 12311 31433
rect 13078 31424 13084 31436
rect 13136 31424 13142 31476
rect 13538 31424 13544 31476
rect 13596 31464 13602 31476
rect 15378 31464 15384 31476
rect 13596 31436 15148 31464
rect 13596 31424 13602 31436
rect 5534 31356 5540 31408
rect 5592 31396 5598 31408
rect 5813 31399 5871 31405
rect 5813 31396 5825 31399
rect 5592 31368 5825 31396
rect 5592 31356 5598 31368
rect 5813 31365 5825 31368
rect 5859 31365 5871 31399
rect 5813 31359 5871 31365
rect 6546 31356 6552 31408
rect 6604 31396 6610 31408
rect 13388 31399 13446 31405
rect 6604 31368 6773 31396
rect 6604 31356 6610 31368
rect 6745 31340 6773 31368
rect 13388 31365 13400 31399
rect 13434 31396 13446 31399
rect 14090 31396 14096 31408
rect 13434 31368 14096 31396
rect 13434 31365 13446 31368
rect 13388 31359 13446 31365
rect 14090 31356 14096 31368
rect 14148 31356 14154 31408
rect 2593 31331 2651 31337
rect 2593 31297 2605 31331
rect 2639 31297 2651 31331
rect 2593 31291 2651 31297
rect 2777 31331 2835 31337
rect 2777 31297 2789 31331
rect 2823 31328 2835 31331
rect 2866 31328 2872 31340
rect 2823 31300 2872 31328
rect 2823 31297 2835 31300
rect 2777 31291 2835 31297
rect 2608 31260 2636 31291
rect 2866 31288 2872 31300
rect 2924 31328 2930 31340
rect 3326 31328 3332 31340
rect 2924 31300 3332 31328
rect 2924 31288 2930 31300
rect 3326 31288 3332 31300
rect 3384 31288 3390 31340
rect 5626 31328 5632 31340
rect 5587 31300 5632 31328
rect 5626 31288 5632 31300
rect 5684 31288 5690 31340
rect 6641 31331 6699 31337
rect 6641 31297 6653 31331
rect 6687 31297 6699 31331
rect 6641 31291 6699 31297
rect 6730 31334 6788 31340
rect 6730 31300 6742 31334
rect 6776 31300 6788 31334
rect 6730 31294 6788 31300
rect 3602 31260 3608 31272
rect 2608 31232 3608 31260
rect 3602 31220 3608 31232
rect 3660 31220 3666 31272
rect 6656 31260 6684 31291
rect 6822 31288 6828 31340
rect 6880 31337 6886 31340
rect 6880 31328 6888 31337
rect 7009 31331 7067 31337
rect 6880 31300 6925 31328
rect 6880 31291 6888 31300
rect 7009 31297 7021 31331
rect 7055 31328 7067 31331
rect 7374 31328 7380 31340
rect 7055 31300 7380 31328
rect 7055 31297 7067 31300
rect 7009 31291 7067 31297
rect 6880 31288 6886 31291
rect 7374 31288 7380 31300
rect 7432 31288 7438 31340
rect 9585 31331 9643 31337
rect 9585 31297 9597 31331
rect 9631 31328 9643 31331
rect 10134 31328 10140 31340
rect 9631 31300 10140 31328
rect 9631 31297 9643 31300
rect 9585 31291 9643 31297
rect 10134 31288 10140 31300
rect 10192 31288 10198 31340
rect 14918 31328 14924 31340
rect 14879 31300 14924 31328
rect 14918 31288 14924 31300
rect 14976 31288 14982 31340
rect 15014 31331 15072 31337
rect 15014 31297 15026 31331
rect 15060 31328 15072 31331
rect 15120 31328 15148 31436
rect 15212 31436 15384 31464
rect 15212 31405 15240 31436
rect 15378 31424 15384 31436
rect 15436 31464 15442 31476
rect 16022 31464 16028 31476
rect 15436 31436 16028 31464
rect 15436 31424 15442 31436
rect 16022 31424 16028 31436
rect 16080 31424 16086 31476
rect 16761 31467 16819 31473
rect 16761 31433 16773 31467
rect 16807 31464 16819 31467
rect 16850 31464 16856 31476
rect 16807 31436 16856 31464
rect 16807 31433 16819 31436
rect 16761 31427 16819 31433
rect 16850 31424 16856 31436
rect 16908 31424 16914 31476
rect 25225 31467 25283 31473
rect 25225 31433 25237 31467
rect 25271 31464 25283 31467
rect 25314 31464 25320 31476
rect 25271 31436 25320 31464
rect 25271 31433 25283 31436
rect 25225 31427 25283 31433
rect 25314 31424 25320 31436
rect 25372 31424 25378 31476
rect 25958 31424 25964 31476
rect 26016 31464 26022 31476
rect 26053 31467 26111 31473
rect 26053 31464 26065 31467
rect 26016 31436 26065 31464
rect 26016 31424 26022 31436
rect 26053 31433 26065 31436
rect 26099 31433 26111 31467
rect 32122 31464 32128 31476
rect 32083 31436 32128 31464
rect 26053 31427 26111 31433
rect 32122 31424 32128 31436
rect 32180 31464 32186 31476
rect 36170 31464 36176 31476
rect 32180 31436 32996 31464
rect 36131 31436 36176 31464
rect 32180 31424 32186 31436
rect 15197 31399 15255 31405
rect 15197 31365 15209 31399
rect 15243 31365 15255 31399
rect 15197 31359 15255 31365
rect 15289 31399 15347 31405
rect 15289 31365 15301 31399
rect 15335 31396 15347 31399
rect 15470 31396 15476 31408
rect 15335 31368 15476 31396
rect 15335 31365 15347 31368
rect 15289 31359 15347 31365
rect 15470 31356 15476 31368
rect 15528 31356 15534 31408
rect 28534 31396 28540 31408
rect 17595 31368 28540 31396
rect 15060 31300 15148 31328
rect 15386 31331 15444 31337
rect 15060 31297 15072 31300
rect 15014 31291 15072 31297
rect 15386 31297 15398 31331
rect 15432 31297 15444 31331
rect 16942 31328 16948 31340
rect 15386 31291 15444 31297
rect 16592 31300 16948 31328
rect 7926 31260 7932 31272
rect 6656 31232 7932 31260
rect 7926 31220 7932 31232
rect 7984 31220 7990 31272
rect 13633 31263 13691 31269
rect 13633 31229 13645 31263
rect 13679 31260 13691 31263
rect 15194 31260 15200 31272
rect 13679 31232 15200 31260
rect 13679 31229 13691 31232
rect 13633 31223 13691 31229
rect 15194 31220 15200 31232
rect 15252 31220 15258 31272
rect 15401 31260 15429 31291
rect 16592 31272 16620 31300
rect 16942 31288 16948 31300
rect 17000 31288 17006 31340
rect 16574 31260 16580 31272
rect 15401 31232 16580 31260
rect 13906 31152 13912 31204
rect 13964 31192 13970 31204
rect 14642 31192 14648 31204
rect 13964 31164 14648 31192
rect 13964 31152 13970 31164
rect 14642 31152 14648 31164
rect 14700 31192 14706 31204
rect 15401 31192 15429 31232
rect 16574 31220 16580 31232
rect 16632 31220 16638 31272
rect 16666 31220 16672 31272
rect 16724 31260 16730 31272
rect 17497 31263 17555 31269
rect 17497 31260 17509 31263
rect 16724 31232 17509 31260
rect 16724 31220 16730 31232
rect 17497 31229 17509 31232
rect 17543 31229 17555 31263
rect 17497 31223 17555 31229
rect 17595 31192 17623 31368
rect 28534 31356 28540 31368
rect 28592 31356 28598 31408
rect 31113 31399 31171 31405
rect 31113 31365 31125 31399
rect 31159 31396 31171 31399
rect 31570 31396 31576 31408
rect 31159 31368 31576 31396
rect 31159 31365 31171 31368
rect 31113 31359 31171 31365
rect 31570 31356 31576 31368
rect 31628 31356 31634 31408
rect 32968 31405 32996 31436
rect 36170 31424 36176 31436
rect 36228 31424 36234 31476
rect 32953 31399 33011 31405
rect 32953 31365 32965 31399
rect 32999 31365 33011 31399
rect 32953 31359 33011 31365
rect 17773 31331 17831 31337
rect 17773 31297 17785 31331
rect 17819 31328 17831 31331
rect 18690 31328 18696 31340
rect 17819 31300 18696 31328
rect 17819 31297 17831 31300
rect 17773 31291 17831 31297
rect 18690 31288 18696 31300
rect 18748 31288 18754 31340
rect 19696 31331 19754 31337
rect 19696 31297 19708 31331
rect 19742 31328 19754 31331
rect 19978 31328 19984 31340
rect 19742 31300 19984 31328
rect 19742 31297 19754 31300
rect 19696 31291 19754 31297
rect 19978 31288 19984 31300
rect 20036 31288 20042 31340
rect 20990 31288 20996 31340
rect 21048 31328 21054 31340
rect 21450 31328 21456 31340
rect 21048 31300 21456 31328
rect 21048 31288 21054 31300
rect 21450 31288 21456 31300
rect 21508 31328 21514 31340
rect 22465 31331 22523 31337
rect 22465 31328 22477 31331
rect 21508 31300 22477 31328
rect 21508 31288 21514 31300
rect 22465 31297 22477 31300
rect 22511 31297 22523 31331
rect 22465 31291 22523 31297
rect 22649 31331 22707 31337
rect 22649 31297 22661 31331
rect 22695 31328 22707 31331
rect 23382 31328 23388 31340
rect 22695 31300 23388 31328
rect 22695 31297 22707 31300
rect 22649 31291 22707 31297
rect 23382 31288 23388 31300
rect 23440 31288 23446 31340
rect 23842 31288 23848 31340
rect 23900 31328 23906 31340
rect 23937 31331 23995 31337
rect 23937 31328 23949 31331
rect 23900 31300 23949 31328
rect 23900 31288 23906 31300
rect 23937 31297 23949 31300
rect 23983 31297 23995 31331
rect 23937 31291 23995 31297
rect 24026 31288 24032 31340
rect 24084 31288 24090 31340
rect 25409 31331 25467 31337
rect 25409 31297 25421 31331
rect 25455 31297 25467 31331
rect 25409 31291 25467 31297
rect 17862 31220 17868 31272
rect 17920 31260 17926 31272
rect 19429 31263 19487 31269
rect 19429 31260 19441 31263
rect 17920 31232 19441 31260
rect 17920 31220 17926 31232
rect 19429 31229 19441 31232
rect 19475 31229 19487 31263
rect 19429 31223 19487 31229
rect 23293 31263 23351 31269
rect 23293 31229 23305 31263
rect 23339 31260 23351 31263
rect 23860 31260 23888 31288
rect 23339 31232 23888 31260
rect 24044 31260 24072 31288
rect 24673 31263 24731 31269
rect 24673 31260 24685 31263
rect 24044 31232 24685 31260
rect 23339 31229 23351 31232
rect 23293 31223 23351 31229
rect 24673 31229 24685 31232
rect 24719 31260 24731 31263
rect 25424 31260 25452 31291
rect 25498 31288 25504 31340
rect 25556 31328 25562 31340
rect 25869 31331 25927 31337
rect 25869 31328 25881 31331
rect 25556 31300 25881 31328
rect 25556 31288 25562 31300
rect 25869 31297 25881 31300
rect 25915 31328 25927 31331
rect 26050 31328 26056 31340
rect 25915 31300 26056 31328
rect 25915 31297 25927 31300
rect 25869 31291 25927 31297
rect 26050 31288 26056 31300
rect 26108 31288 26114 31340
rect 28074 31288 28080 31340
rect 28132 31328 28138 31340
rect 30377 31331 30435 31337
rect 30377 31328 30389 31331
rect 28132 31300 30389 31328
rect 28132 31288 28138 31300
rect 30377 31297 30389 31300
rect 30423 31297 30435 31331
rect 30377 31291 30435 31297
rect 30926 31288 30932 31340
rect 30984 31328 30990 31340
rect 31021 31331 31079 31337
rect 31021 31328 31033 31331
rect 30984 31300 31033 31328
rect 30984 31288 30990 31300
rect 31021 31297 31033 31300
rect 31067 31297 31079 31331
rect 31202 31328 31208 31340
rect 31163 31300 31208 31328
rect 31021 31291 31079 31297
rect 31202 31288 31208 31300
rect 31260 31288 31266 31340
rect 31389 31331 31447 31337
rect 31389 31297 31401 31331
rect 31435 31328 31447 31331
rect 31938 31328 31944 31340
rect 31435 31300 31944 31328
rect 31435 31297 31447 31300
rect 31389 31291 31447 31297
rect 31938 31288 31944 31300
rect 31996 31288 32002 31340
rect 32309 31331 32367 31337
rect 32309 31297 32321 31331
rect 32355 31297 32367 31331
rect 32309 31291 32367 31297
rect 28534 31260 28540 31272
rect 24719 31232 28540 31260
rect 24719 31229 24731 31232
rect 24673 31223 24731 31229
rect 28534 31220 28540 31232
rect 28592 31220 28598 31272
rect 30742 31220 30748 31272
rect 30800 31260 30806 31272
rect 32324 31260 32352 31291
rect 32398 31288 32404 31340
rect 32456 31328 32462 31340
rect 33137 31331 33195 31337
rect 32456 31300 32501 31328
rect 32456 31288 32462 31300
rect 33137 31297 33149 31331
rect 33183 31328 33195 31331
rect 33226 31328 33232 31340
rect 33183 31300 33232 31328
rect 33183 31297 33195 31300
rect 33137 31291 33195 31297
rect 33226 31288 33232 31300
rect 33284 31288 33290 31340
rect 35802 31328 35808 31340
rect 35763 31300 35808 31328
rect 35802 31288 35808 31300
rect 35860 31288 35866 31340
rect 35989 31331 36047 31337
rect 35989 31297 36001 31331
rect 36035 31328 36047 31331
rect 37274 31328 37280 31340
rect 36035 31300 37280 31328
rect 36035 31297 36047 31300
rect 35989 31291 36047 31297
rect 30800 31232 32352 31260
rect 30800 31220 30806 31232
rect 33502 31220 33508 31272
rect 33560 31260 33566 31272
rect 36004 31260 36032 31291
rect 37274 31288 37280 31300
rect 37332 31288 37338 31340
rect 37642 31328 37648 31340
rect 37603 31300 37648 31328
rect 37642 31288 37648 31300
rect 37700 31288 37706 31340
rect 33560 31232 36032 31260
rect 33560 31220 33566 31232
rect 14700 31164 15429 31192
rect 15488 31164 17623 31192
rect 14700 31152 14706 31164
rect 2314 31084 2320 31136
rect 2372 31124 2378 31136
rect 3329 31127 3387 31133
rect 3329 31124 3341 31127
rect 2372 31096 3341 31124
rect 2372 31084 2378 31096
rect 3329 31093 3341 31096
rect 3375 31124 3387 31127
rect 4062 31124 4068 31136
rect 3375 31096 4068 31124
rect 3375 31093 3387 31096
rect 3329 31087 3387 31093
rect 4062 31084 4068 31096
rect 4120 31084 4126 31136
rect 6365 31127 6423 31133
rect 6365 31093 6377 31127
rect 6411 31124 6423 31127
rect 6638 31124 6644 31136
rect 6411 31096 6644 31124
rect 6411 31093 6423 31096
rect 6365 31087 6423 31093
rect 6638 31084 6644 31096
rect 6696 31084 6702 31136
rect 10134 31124 10140 31136
rect 10095 31096 10140 31124
rect 10134 31084 10140 31096
rect 10192 31084 10198 31136
rect 12342 31084 12348 31136
rect 12400 31124 12406 31136
rect 15488 31124 15516 31164
rect 12400 31096 15516 31124
rect 15565 31127 15623 31133
rect 12400 31084 12406 31096
rect 15565 31093 15577 31127
rect 15611 31124 15623 31127
rect 16022 31124 16028 31136
rect 15611 31096 16028 31124
rect 15611 31093 15623 31096
rect 15565 31087 15623 31093
rect 16022 31084 16028 31096
rect 16080 31084 16086 31136
rect 20714 31084 20720 31136
rect 20772 31124 20778 31136
rect 20809 31127 20867 31133
rect 20809 31124 20821 31127
rect 20772 31096 20821 31124
rect 20772 31084 20778 31096
rect 20809 31093 20821 31096
rect 20855 31093 20867 31127
rect 20809 31087 20867 31093
rect 22738 31084 22744 31136
rect 22796 31124 22802 31136
rect 22833 31127 22891 31133
rect 22833 31124 22845 31127
rect 22796 31096 22845 31124
rect 22796 31084 22802 31096
rect 22833 31093 22845 31096
rect 22879 31093 22891 31127
rect 24026 31124 24032 31136
rect 23987 31096 24032 31124
rect 22833 31087 22891 31093
rect 24026 31084 24032 31096
rect 24084 31084 24090 31136
rect 28074 31124 28080 31136
rect 28035 31096 28080 31124
rect 28074 31084 28080 31096
rect 28132 31084 28138 31136
rect 28902 31084 28908 31136
rect 28960 31124 28966 31136
rect 29089 31127 29147 31133
rect 29089 31124 29101 31127
rect 28960 31096 29101 31124
rect 28960 31084 28966 31096
rect 29089 31093 29101 31096
rect 29135 31093 29147 31127
rect 29089 31087 29147 31093
rect 30558 31084 30564 31136
rect 30616 31124 30622 31136
rect 30837 31127 30895 31133
rect 30837 31124 30849 31127
rect 30616 31096 30849 31124
rect 30616 31084 30622 31096
rect 30837 31093 30849 31096
rect 30883 31093 30895 31127
rect 30837 31087 30895 31093
rect 32214 31084 32220 31136
rect 32272 31124 32278 31136
rect 33321 31127 33379 31133
rect 33321 31124 33333 31127
rect 32272 31096 33333 31124
rect 32272 31084 32278 31096
rect 33321 31093 33333 31096
rect 33367 31093 33379 31127
rect 38930 31124 38936 31136
rect 38891 31096 38936 31124
rect 33321 31087 33379 31093
rect 38930 31084 38936 31096
rect 38988 31084 38994 31136
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 7926 30880 7932 30932
rect 7984 30920 7990 30932
rect 8205 30923 8263 30929
rect 8205 30920 8217 30923
rect 7984 30892 8217 30920
rect 7984 30880 7990 30892
rect 8205 30889 8217 30892
rect 8251 30920 8263 30923
rect 12342 30920 12348 30932
rect 8251 30892 12348 30920
rect 8251 30889 8263 30892
rect 8205 30883 8263 30889
rect 12342 30880 12348 30892
rect 12400 30880 12406 30932
rect 13357 30923 13415 30929
rect 13357 30889 13369 30923
rect 13403 30920 13415 30923
rect 14918 30920 14924 30932
rect 13403 30892 14924 30920
rect 13403 30889 13415 30892
rect 13357 30883 13415 30889
rect 14918 30880 14924 30892
rect 14976 30880 14982 30932
rect 15105 30923 15163 30929
rect 15105 30889 15117 30923
rect 15151 30920 15163 30923
rect 15470 30920 15476 30932
rect 15151 30892 15476 30920
rect 15151 30889 15163 30892
rect 15105 30883 15163 30889
rect 1854 30784 1860 30796
rect 1815 30756 1860 30784
rect 1854 30744 1860 30756
rect 1912 30744 1918 30796
rect 1872 30716 1900 30744
rect 4525 30719 4583 30725
rect 4525 30716 4537 30719
rect 1872 30688 4537 30716
rect 4525 30685 4537 30688
rect 4571 30716 4583 30719
rect 6365 30719 6423 30725
rect 6365 30716 6377 30719
rect 4571 30688 6377 30716
rect 4571 30685 4583 30688
rect 4525 30679 4583 30685
rect 6365 30685 6377 30688
rect 6411 30716 6423 30719
rect 8202 30716 8208 30728
rect 6411 30688 8208 30716
rect 6411 30685 6423 30688
rect 6365 30679 6423 30685
rect 8202 30676 8208 30688
rect 8260 30676 8266 30728
rect 11054 30676 11060 30728
rect 11112 30716 11118 30728
rect 12805 30719 12863 30725
rect 12805 30716 12817 30719
rect 11112 30688 12817 30716
rect 11112 30676 11118 30688
rect 12805 30685 12817 30688
rect 12851 30685 12863 30719
rect 13078 30716 13084 30728
rect 13039 30688 13084 30716
rect 12805 30679 12863 30685
rect 13078 30676 13084 30688
rect 13136 30676 13142 30728
rect 13170 30676 13176 30728
rect 13228 30716 13234 30728
rect 13228 30688 13273 30716
rect 13228 30676 13234 30688
rect 13814 30676 13820 30728
rect 13872 30716 13878 30728
rect 14274 30716 14280 30728
rect 13872 30688 14280 30716
rect 13872 30676 13878 30688
rect 14274 30676 14280 30688
rect 14332 30676 14338 30728
rect 14461 30719 14519 30725
rect 14461 30685 14473 30719
rect 14507 30716 14519 30719
rect 15120 30716 15148 30883
rect 15470 30880 15476 30892
rect 15528 30880 15534 30932
rect 16758 30880 16764 30932
rect 16816 30920 16822 30932
rect 21729 30923 21787 30929
rect 21729 30920 21741 30923
rect 16816 30892 21741 30920
rect 16816 30880 16822 30892
rect 21729 30889 21741 30892
rect 21775 30889 21787 30923
rect 39301 30923 39359 30929
rect 39301 30920 39313 30923
rect 21729 30883 21787 30889
rect 35360 30892 39313 30920
rect 18693 30855 18751 30861
rect 18693 30821 18705 30855
rect 18739 30852 18751 30855
rect 20070 30852 20076 30864
rect 18739 30824 20076 30852
rect 18739 30821 18751 30824
rect 18693 30815 18751 30821
rect 20070 30812 20076 30824
rect 20128 30812 20134 30864
rect 14507 30688 15148 30716
rect 14507 30685 14519 30688
rect 14461 30679 14519 30685
rect 15194 30676 15200 30728
rect 15252 30716 15258 30728
rect 15746 30716 15752 30728
rect 15252 30688 15752 30716
rect 15252 30676 15258 30688
rect 15746 30676 15752 30688
rect 15804 30716 15810 30728
rect 16485 30719 16543 30725
rect 16485 30716 16497 30719
rect 15804 30688 16497 30716
rect 15804 30676 15810 30688
rect 16485 30685 16497 30688
rect 16531 30716 16543 30719
rect 17313 30719 17371 30725
rect 17313 30716 17325 30719
rect 16531 30688 17325 30716
rect 16531 30685 16543 30688
rect 16485 30679 16543 30685
rect 17313 30685 17325 30688
rect 17359 30716 17371 30719
rect 17862 30716 17868 30728
rect 17359 30688 17868 30716
rect 17359 30685 17371 30688
rect 17313 30679 17371 30685
rect 17862 30676 17868 30688
rect 17920 30676 17926 30728
rect 21744 30716 21772 30883
rect 22554 30812 22560 30864
rect 22612 30852 22618 30864
rect 28537 30855 28595 30861
rect 22612 30824 22968 30852
rect 22612 30812 22618 30824
rect 22462 30744 22468 30796
rect 22520 30784 22526 30796
rect 22520 30756 22692 30784
rect 22520 30744 22526 30756
rect 22664 30725 22692 30756
rect 22557 30719 22615 30725
rect 22557 30716 22569 30719
rect 21744 30688 22569 30716
rect 22557 30685 22569 30688
rect 22603 30685 22615 30719
rect 22557 30679 22615 30685
rect 22649 30719 22707 30725
rect 22649 30685 22661 30719
rect 22695 30685 22707 30719
rect 22649 30679 22707 30685
rect 2130 30657 2136 30660
rect 2124 30611 2136 30657
rect 2188 30648 2194 30660
rect 4798 30657 4804 30660
rect 4792 30648 4804 30657
rect 2188 30620 2224 30648
rect 4759 30620 4804 30648
rect 2130 30608 2136 30611
rect 2188 30608 2194 30620
rect 4792 30611 4804 30620
rect 4798 30608 4804 30611
rect 4856 30608 4862 30660
rect 6638 30657 6644 30660
rect 6632 30648 6644 30657
rect 6599 30620 6644 30648
rect 6632 30611 6644 30620
rect 6638 30608 6644 30611
rect 6696 30608 6702 30660
rect 12989 30651 13047 30657
rect 12989 30617 13001 30651
rect 13035 30648 13047 30651
rect 13262 30648 13268 30660
rect 13035 30620 13268 30648
rect 13035 30617 13047 30620
rect 12989 30611 13047 30617
rect 13262 30608 13268 30620
rect 13320 30608 13326 30660
rect 15654 30608 15660 30660
rect 15712 30648 15718 30660
rect 16218 30651 16276 30657
rect 16218 30648 16230 30651
rect 15712 30620 16230 30648
rect 15712 30608 15718 30620
rect 16218 30617 16230 30620
rect 16264 30617 16276 30651
rect 16218 30611 16276 30617
rect 17580 30651 17638 30657
rect 17580 30617 17592 30651
rect 17626 30648 17638 30651
rect 18046 30648 18052 30660
rect 17626 30620 18052 30648
rect 17626 30617 17638 30620
rect 17580 30611 17638 30617
rect 18046 30608 18052 30620
rect 18104 30608 18110 30660
rect 22572 30648 22600 30679
rect 22738 30676 22744 30728
rect 22796 30716 22802 30728
rect 22940 30725 22968 30824
rect 28537 30821 28549 30855
rect 28583 30821 28595 30855
rect 28537 30815 28595 30821
rect 26789 30787 26847 30793
rect 26789 30753 26801 30787
rect 26835 30784 26847 30787
rect 27246 30784 27252 30796
rect 26835 30756 27252 30784
rect 26835 30753 26847 30756
rect 26789 30747 26847 30753
rect 27246 30744 27252 30756
rect 27304 30784 27310 30796
rect 28552 30784 28580 30815
rect 32306 30812 32312 30864
rect 32364 30812 32370 30864
rect 33229 30855 33287 30861
rect 33229 30821 33241 30855
rect 33275 30852 33287 30855
rect 34054 30852 34060 30864
rect 33275 30824 34060 30852
rect 33275 30821 33287 30824
rect 33229 30815 33287 30821
rect 34054 30812 34060 30824
rect 34112 30812 34118 30864
rect 27304 30756 28580 30784
rect 27304 30744 27310 30756
rect 30282 30744 30288 30796
rect 30340 30784 30346 30796
rect 30377 30787 30435 30793
rect 30377 30784 30389 30787
rect 30340 30756 30389 30784
rect 30340 30744 30346 30756
rect 30377 30753 30389 30756
rect 30423 30753 30435 30787
rect 30377 30747 30435 30753
rect 22925 30719 22983 30725
rect 22796 30688 22841 30716
rect 22796 30676 22802 30688
rect 22925 30685 22937 30719
rect 22971 30685 22983 30719
rect 22925 30679 22983 30685
rect 24302 30676 24308 30728
rect 24360 30716 24366 30728
rect 24489 30719 24547 30725
rect 24489 30716 24501 30719
rect 24360 30688 24501 30716
rect 24360 30676 24366 30688
rect 24489 30685 24501 30688
rect 24535 30716 24547 30719
rect 24578 30716 24584 30728
rect 24535 30688 24584 30716
rect 24535 30685 24547 30688
rect 24489 30679 24547 30685
rect 24578 30676 24584 30688
rect 24636 30676 24642 30728
rect 30098 30716 30104 30728
rect 30059 30688 30104 30716
rect 30098 30676 30104 30688
rect 30156 30676 30162 30728
rect 30190 30676 30196 30728
rect 30248 30716 30254 30728
rect 30466 30716 30472 30728
rect 30248 30688 30472 30716
rect 30248 30676 30254 30688
rect 30466 30676 30472 30688
rect 30524 30716 30530 30728
rect 31481 30719 31539 30725
rect 31481 30716 31493 30719
rect 30524 30688 31493 30716
rect 30524 30676 30530 30688
rect 31481 30685 31493 30688
rect 31527 30716 31539 30719
rect 32033 30719 32091 30725
rect 32033 30716 32045 30719
rect 31527 30688 32045 30716
rect 31527 30685 31539 30688
rect 31481 30679 31539 30685
rect 32033 30685 32045 30688
rect 32079 30685 32091 30719
rect 32214 30716 32220 30728
rect 32175 30688 32220 30716
rect 32033 30679 32091 30685
rect 32214 30676 32220 30688
rect 32272 30676 32278 30728
rect 32324 30725 32352 30812
rect 33318 30784 33324 30796
rect 32416 30756 33324 30784
rect 32416 30725 32444 30756
rect 33318 30744 33324 30756
rect 33376 30744 33382 30796
rect 35360 30728 35388 30892
rect 39301 30889 39313 30892
rect 39347 30889 39359 30923
rect 39301 30883 39359 30889
rect 36262 30812 36268 30864
rect 36320 30812 36326 30864
rect 32309 30719 32367 30725
rect 32309 30685 32321 30719
rect 32355 30685 32367 30719
rect 32309 30679 32367 30685
rect 32401 30719 32459 30725
rect 32401 30685 32413 30719
rect 32447 30685 32459 30719
rect 33410 30716 33416 30728
rect 33371 30688 33416 30716
rect 32401 30679 32459 30685
rect 33410 30676 33416 30688
rect 33468 30676 33474 30728
rect 33502 30676 33508 30728
rect 33560 30716 33566 30728
rect 33778 30716 33784 30728
rect 33560 30688 33605 30716
rect 33739 30688 33784 30716
rect 33560 30676 33566 30688
rect 33778 30676 33784 30688
rect 33836 30676 33842 30728
rect 35342 30716 35348 30728
rect 35255 30688 35348 30716
rect 35342 30676 35348 30688
rect 35400 30676 35406 30728
rect 35986 30716 35992 30728
rect 35947 30688 35992 30716
rect 35986 30676 35992 30688
rect 36044 30676 36050 30728
rect 36280 30725 36308 30812
rect 36173 30719 36231 30725
rect 36173 30685 36185 30719
rect 36219 30685 36231 30719
rect 36173 30679 36231 30685
rect 36268 30719 36326 30725
rect 36268 30685 36280 30719
rect 36314 30685 36326 30719
rect 36268 30679 36326 30685
rect 36357 30719 36415 30725
rect 36357 30685 36369 30719
rect 36403 30716 36415 30719
rect 37093 30719 37151 30725
rect 37093 30716 37105 30719
rect 36403 30688 37105 30716
rect 36403 30685 36415 30688
rect 36357 30679 36415 30685
rect 37093 30685 37105 30688
rect 37139 30685 37151 30719
rect 37918 30716 37924 30728
rect 37879 30688 37924 30716
rect 37093 30679 37151 30685
rect 24118 30648 24124 30660
rect 22572 30620 24124 30648
rect 24118 30608 24124 30620
rect 24176 30608 24182 30660
rect 24670 30648 24676 30660
rect 24631 30620 24676 30648
rect 24670 30608 24676 30620
rect 24728 30648 24734 30660
rect 24728 30620 25452 30648
rect 24728 30608 24734 30620
rect 3237 30583 3295 30589
rect 3237 30549 3249 30583
rect 3283 30580 3295 30583
rect 3418 30580 3424 30592
rect 3283 30552 3424 30580
rect 3283 30549 3295 30552
rect 3237 30543 3295 30549
rect 3418 30540 3424 30552
rect 3476 30540 3482 30592
rect 5626 30540 5632 30592
rect 5684 30580 5690 30592
rect 5905 30583 5963 30589
rect 5905 30580 5917 30583
rect 5684 30552 5917 30580
rect 5684 30540 5690 30552
rect 5905 30549 5917 30552
rect 5951 30580 5963 30583
rect 6730 30580 6736 30592
rect 5951 30552 6736 30580
rect 5951 30549 5963 30552
rect 5905 30543 5963 30549
rect 6730 30540 6736 30552
rect 6788 30540 6794 30592
rect 7006 30540 7012 30592
rect 7064 30580 7070 30592
rect 7745 30583 7803 30589
rect 7745 30580 7757 30583
rect 7064 30552 7757 30580
rect 7064 30540 7070 30552
rect 7745 30549 7757 30552
rect 7791 30549 7803 30583
rect 7745 30543 7803 30549
rect 9953 30583 10011 30589
rect 9953 30549 9965 30583
rect 9999 30580 10011 30583
rect 10042 30580 10048 30592
rect 9999 30552 10048 30580
rect 9999 30549 10011 30552
rect 9953 30543 10011 30549
rect 10042 30540 10048 30552
rect 10100 30540 10106 30592
rect 14645 30583 14703 30589
rect 14645 30549 14657 30583
rect 14691 30580 14703 30583
rect 15194 30580 15200 30592
rect 14691 30552 15200 30580
rect 14691 30549 14703 30552
rect 14645 30543 14703 30549
rect 15194 30540 15200 30552
rect 15252 30540 15258 30592
rect 19334 30580 19340 30592
rect 19295 30552 19340 30580
rect 19334 30540 19340 30552
rect 19392 30540 19398 30592
rect 20254 30580 20260 30592
rect 20215 30552 20260 30580
rect 20254 30540 20260 30552
rect 20312 30540 20318 30592
rect 22281 30583 22339 30589
rect 22281 30549 22293 30583
rect 22327 30580 22339 30583
rect 22370 30580 22376 30592
rect 22327 30552 22376 30580
rect 22327 30549 22339 30552
rect 22281 30543 22339 30549
rect 22370 30540 22376 30552
rect 22428 30540 22434 30592
rect 24857 30583 24915 30589
rect 24857 30549 24869 30583
rect 24903 30580 24915 30583
rect 25314 30580 25320 30592
rect 24903 30552 25320 30580
rect 24903 30549 24915 30552
rect 24857 30543 24915 30549
rect 25314 30540 25320 30552
rect 25372 30540 25378 30592
rect 25424 30589 25452 30620
rect 26234 30608 26240 30660
rect 26292 30648 26298 30660
rect 26522 30651 26580 30657
rect 26522 30648 26534 30651
rect 26292 30620 26534 30648
rect 26292 30608 26298 30620
rect 26522 30617 26534 30620
rect 26568 30617 26580 30651
rect 26522 30611 26580 30617
rect 27249 30651 27307 30657
rect 27249 30617 27261 30651
rect 27295 30617 27307 30651
rect 27249 30611 27307 30617
rect 25409 30583 25467 30589
rect 25409 30549 25421 30583
rect 25455 30549 25467 30583
rect 27264 30580 27292 30611
rect 31202 30608 31208 30660
rect 31260 30648 31266 30660
rect 33594 30648 33600 30660
rect 31260 30620 33600 30648
rect 31260 30608 31266 30620
rect 33594 30608 33600 30620
rect 33652 30608 33658 30660
rect 35158 30648 35164 30660
rect 35119 30620 35164 30648
rect 35158 30608 35164 30620
rect 35216 30608 35222 30660
rect 35529 30651 35587 30657
rect 35529 30617 35541 30651
rect 35575 30648 35587 30651
rect 36188 30648 36216 30679
rect 35575 30620 36216 30648
rect 35575 30617 35587 30620
rect 35529 30611 35587 30617
rect 28902 30580 28908 30592
rect 27264 30552 28908 30580
rect 25409 30543 25467 30549
rect 28902 30540 28908 30552
rect 28960 30580 28966 30592
rect 29641 30583 29699 30589
rect 29641 30580 29653 30583
rect 28960 30552 29653 30580
rect 28960 30540 28966 30552
rect 29641 30549 29653 30552
rect 29687 30580 29699 30583
rect 30374 30580 30380 30592
rect 29687 30552 30380 30580
rect 29687 30549 29699 30552
rect 29641 30543 29699 30549
rect 30374 30540 30380 30552
rect 30432 30540 30438 30592
rect 32677 30583 32735 30589
rect 32677 30549 32689 30583
rect 32723 30580 32735 30583
rect 33134 30580 33140 30592
rect 32723 30552 33140 30580
rect 32723 30549 32735 30552
rect 32677 30543 32735 30549
rect 33134 30540 33140 30552
rect 33192 30540 33198 30592
rect 33870 30540 33876 30592
rect 33928 30580 33934 30592
rect 36372 30580 36400 30679
rect 37918 30676 37924 30688
rect 37976 30716 37982 30728
rect 38562 30716 38568 30728
rect 37976 30688 38568 30716
rect 37976 30676 37982 30688
rect 38562 30676 38568 30688
rect 38620 30716 38626 30728
rect 38930 30716 38936 30728
rect 38620 30688 38936 30716
rect 38620 30676 38626 30688
rect 38930 30676 38936 30688
rect 38988 30676 38994 30728
rect 58158 30716 58164 30728
rect 58119 30688 58164 30716
rect 58158 30676 58164 30688
rect 58216 30676 58222 30728
rect 36633 30651 36691 30657
rect 36633 30617 36645 30651
rect 36679 30648 36691 30651
rect 38166 30651 38224 30657
rect 38166 30648 38178 30651
rect 36679 30620 38178 30648
rect 36679 30617 36691 30620
rect 36633 30611 36691 30617
rect 38166 30617 38178 30620
rect 38212 30617 38224 30651
rect 38166 30611 38224 30617
rect 33928 30552 36400 30580
rect 33928 30540 33934 30552
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 2130 30376 2136 30388
rect 2091 30348 2136 30376
rect 2130 30336 2136 30348
rect 2188 30336 2194 30388
rect 7374 30376 7380 30388
rect 7287 30348 7380 30376
rect 7374 30336 7380 30348
rect 7432 30376 7438 30388
rect 30190 30376 30196 30388
rect 7432 30348 30196 30376
rect 7432 30336 7438 30348
rect 30190 30336 30196 30348
rect 30248 30336 30254 30388
rect 30374 30336 30380 30388
rect 30432 30376 30438 30388
rect 37642 30376 37648 30388
rect 30432 30348 37648 30376
rect 30432 30336 30438 30348
rect 37642 30336 37648 30348
rect 37700 30336 37706 30388
rect 2866 30308 2872 30320
rect 2424 30280 2872 30308
rect 2424 30249 2452 30280
rect 2866 30268 2872 30280
rect 2924 30268 2930 30320
rect 3326 30268 3332 30320
rect 3384 30308 3390 30320
rect 3605 30311 3663 30317
rect 3605 30308 3617 30311
rect 3384 30280 3617 30308
rect 3384 30268 3390 30280
rect 3605 30277 3617 30280
rect 3651 30277 3663 30311
rect 3605 30271 3663 30277
rect 7558 30268 7564 30320
rect 7616 30308 7622 30320
rect 7929 30311 7987 30317
rect 7929 30308 7941 30311
rect 7616 30280 7941 30308
rect 7616 30268 7622 30280
rect 7929 30277 7941 30280
rect 7975 30277 7987 30311
rect 7929 30271 7987 30277
rect 8113 30311 8171 30317
rect 8113 30277 8125 30311
rect 8159 30308 8171 30311
rect 8386 30308 8392 30320
rect 8159 30280 8392 30308
rect 8159 30277 8171 30280
rect 8113 30271 8171 30277
rect 8386 30268 8392 30280
rect 8444 30308 8450 30320
rect 10229 30311 10287 30317
rect 10229 30308 10241 30311
rect 8444 30280 9536 30308
rect 8444 30268 8450 30280
rect 2389 30243 2452 30249
rect 2389 30209 2401 30243
rect 2435 30212 2452 30243
rect 2482 30243 2540 30249
rect 2435 30209 2447 30212
rect 2389 30203 2447 30209
rect 2482 30209 2494 30243
rect 2528 30209 2540 30243
rect 2482 30203 2540 30209
rect 2593 30243 2651 30249
rect 2593 30209 2605 30243
rect 2639 30209 2651 30243
rect 2593 30203 2651 30209
rect 2497 30104 2525 30203
rect 2608 30172 2636 30203
rect 2774 30200 2780 30252
rect 2832 30240 2838 30252
rect 3142 30240 3148 30252
rect 2832 30212 3148 30240
rect 2832 30200 2838 30212
rect 3142 30200 3148 30212
rect 3200 30200 3206 30252
rect 3418 30240 3424 30252
rect 3379 30212 3424 30240
rect 3418 30200 3424 30212
rect 3476 30200 3482 30252
rect 9508 30249 9536 30280
rect 9600 30280 10241 30308
rect 9600 30249 9628 30280
rect 10229 30277 10241 30280
rect 10275 30277 10287 30311
rect 10229 30271 10287 30277
rect 10597 30311 10655 30317
rect 10597 30277 10609 30311
rect 10643 30308 10655 30311
rect 10962 30308 10968 30320
rect 10643 30280 10968 30308
rect 10643 30277 10655 30280
rect 10597 30271 10655 30277
rect 10962 30268 10968 30280
rect 11020 30308 11026 30320
rect 11609 30311 11667 30317
rect 11609 30308 11621 30311
rect 11020 30280 11621 30308
rect 11020 30268 11026 30280
rect 11609 30277 11621 30280
rect 11655 30277 11667 30311
rect 15654 30308 15660 30320
rect 15615 30280 15660 30308
rect 11609 30271 11667 30277
rect 15654 30268 15660 30280
rect 15712 30268 15718 30320
rect 16114 30268 16120 30320
rect 16172 30308 16178 30320
rect 18046 30308 18052 30320
rect 16172 30280 17448 30308
rect 18007 30280 18052 30308
rect 16172 30268 16178 30280
rect 17420 30252 17448 30280
rect 18046 30268 18052 30280
rect 18104 30268 18110 30320
rect 19242 30308 19248 30320
rect 18432 30280 19248 30308
rect 9401 30243 9459 30249
rect 9401 30209 9413 30243
rect 9447 30209 9459 30243
rect 9401 30203 9459 30209
rect 9493 30243 9551 30249
rect 9493 30209 9505 30243
rect 9539 30209 9551 30243
rect 9493 30203 9551 30209
rect 9585 30243 9643 30249
rect 9585 30209 9597 30243
rect 9631 30209 9643 30243
rect 9585 30203 9643 30209
rect 9769 30243 9827 30249
rect 9769 30209 9781 30243
rect 9815 30240 9827 30243
rect 9858 30240 9864 30252
rect 9815 30212 9864 30240
rect 9815 30209 9827 30212
rect 9769 30203 9827 30209
rect 3237 30175 3295 30181
rect 3237 30172 3249 30175
rect 2608 30144 3249 30172
rect 3237 30141 3249 30144
rect 3283 30141 3295 30175
rect 9416 30172 9444 30203
rect 9858 30200 9864 30212
rect 9916 30200 9922 30252
rect 10413 30243 10471 30249
rect 10413 30209 10425 30243
rect 10459 30240 10471 30243
rect 11054 30240 11060 30252
rect 10459 30212 11060 30240
rect 10459 30209 10471 30212
rect 10413 30203 10471 30209
rect 11054 30200 11060 30212
rect 11112 30200 11118 30252
rect 11698 30200 11704 30252
rect 11756 30240 11762 30252
rect 11793 30243 11851 30249
rect 11793 30240 11805 30243
rect 11756 30212 11805 30240
rect 11756 30200 11762 30212
rect 11793 30209 11805 30212
rect 11839 30209 11851 30243
rect 11793 30203 11851 30209
rect 14550 30200 14556 30252
rect 14608 30240 14614 30252
rect 15010 30240 15016 30252
rect 14608 30212 15016 30240
rect 14608 30200 14614 30212
rect 15010 30200 15016 30212
rect 15068 30200 15074 30252
rect 15194 30240 15200 30252
rect 15155 30212 15200 30240
rect 15194 30200 15200 30212
rect 15252 30200 15258 30252
rect 15292 30243 15350 30249
rect 15292 30209 15304 30243
rect 15338 30209 15350 30243
rect 15292 30203 15350 30209
rect 15381 30243 15439 30249
rect 15381 30209 15393 30243
rect 15427 30240 15439 30243
rect 15838 30240 15844 30252
rect 15427 30212 15844 30240
rect 15427 30209 15439 30212
rect 15381 30203 15439 30209
rect 10042 30172 10048 30184
rect 9416 30144 10048 30172
rect 3237 30135 3295 30141
rect 10042 30132 10048 30144
rect 10100 30132 10106 30184
rect 11882 30132 11888 30184
rect 11940 30172 11946 30184
rect 11977 30175 12035 30181
rect 11977 30172 11989 30175
rect 11940 30144 11989 30172
rect 11940 30132 11946 30144
rect 11977 30141 11989 30144
rect 12023 30172 12035 30175
rect 12023 30144 12434 30172
rect 12023 30141 12035 30144
rect 11977 30135 12035 30141
rect 2682 30104 2688 30116
rect 2497 30076 2688 30104
rect 2682 30064 2688 30076
rect 2740 30064 2746 30116
rect 9125 30039 9183 30045
rect 9125 30005 9137 30039
rect 9171 30036 9183 30039
rect 9214 30036 9220 30048
rect 9171 30008 9220 30036
rect 9171 30005 9183 30008
rect 9125 29999 9183 30005
rect 9214 29996 9220 30008
rect 9272 29996 9278 30048
rect 12406 30036 12434 30144
rect 14274 30064 14280 30116
rect 14332 30104 14338 30116
rect 15304 30104 15332 30203
rect 15838 30200 15844 30212
rect 15896 30200 15902 30252
rect 16574 30200 16580 30252
rect 16632 30240 16638 30252
rect 16853 30243 16911 30249
rect 16853 30240 16865 30243
rect 16632 30212 16865 30240
rect 16632 30200 16638 30212
rect 16853 30209 16865 30212
rect 16899 30209 16911 30243
rect 16853 30203 16911 30209
rect 17402 30200 17408 30252
rect 17460 30240 17466 30252
rect 18432 30249 18460 30280
rect 19242 30268 19248 30280
rect 19300 30308 19306 30320
rect 19702 30308 19708 30320
rect 19300 30280 19708 30308
rect 19300 30268 19306 30280
rect 18325 30243 18383 30249
rect 18325 30240 18337 30243
rect 17460 30212 18337 30240
rect 17460 30200 17466 30212
rect 18325 30209 18337 30212
rect 18371 30209 18383 30243
rect 18325 30203 18383 30209
rect 18417 30243 18475 30249
rect 18417 30209 18429 30243
rect 18463 30209 18475 30243
rect 18417 30203 18475 30209
rect 16758 30132 16764 30184
rect 16816 30172 16822 30184
rect 17037 30175 17095 30181
rect 17037 30172 17049 30175
rect 16816 30144 17049 30172
rect 16816 30132 16822 30144
rect 17037 30141 17049 30144
rect 17083 30141 17095 30175
rect 18432 30172 18460 30203
rect 18506 30200 18512 30252
rect 18564 30240 18570 30252
rect 18693 30243 18751 30249
rect 18564 30212 18609 30240
rect 18564 30200 18570 30212
rect 18693 30209 18705 30243
rect 18739 30240 18751 30243
rect 19153 30243 19211 30249
rect 19153 30240 19165 30243
rect 18739 30212 19165 30240
rect 18739 30209 18751 30212
rect 18693 30203 18751 30209
rect 19153 30209 19165 30212
rect 19199 30209 19211 30243
rect 19334 30240 19340 30252
rect 19295 30212 19340 30240
rect 19153 30203 19211 30209
rect 17037 30135 17095 30141
rect 17512 30144 18460 30172
rect 15562 30104 15568 30116
rect 14332 30076 15148 30104
rect 15304 30076 15568 30104
rect 14332 30064 14338 30076
rect 12529 30039 12587 30045
rect 12529 30036 12541 30039
rect 12406 30008 12541 30036
rect 12529 30005 12541 30008
rect 12575 30036 12587 30039
rect 14734 30036 14740 30048
rect 12575 30008 14740 30036
rect 12575 30005 12587 30008
rect 12529 29999 12587 30005
rect 14734 29996 14740 30008
rect 14792 29996 14798 30048
rect 15120 30036 15148 30076
rect 15562 30064 15568 30076
rect 15620 30064 15626 30116
rect 17512 30048 17540 30144
rect 18598 30132 18604 30184
rect 18656 30172 18662 30184
rect 18708 30172 18736 30203
rect 19334 30200 19340 30212
rect 19392 30200 19398 30252
rect 19444 30249 19472 30280
rect 19702 30268 19708 30280
rect 19760 30268 19766 30320
rect 19797 30311 19855 30317
rect 19797 30277 19809 30311
rect 19843 30308 19855 30311
rect 19978 30308 19984 30320
rect 19843 30280 19984 30308
rect 19843 30277 19855 30280
rect 19797 30271 19855 30277
rect 19978 30268 19984 30280
rect 20036 30268 20042 30320
rect 20438 30308 20444 30320
rect 20088 30280 20444 30308
rect 19429 30243 19487 30249
rect 19429 30209 19441 30243
rect 19475 30209 19487 30243
rect 19429 30203 19487 30209
rect 19521 30243 19579 30249
rect 19521 30209 19533 30243
rect 19567 30209 19579 30243
rect 19521 30203 19579 30209
rect 18656 30144 18736 30172
rect 18656 30132 18662 30144
rect 17954 30064 17960 30116
rect 18012 30104 18018 30116
rect 19536 30104 19564 30203
rect 19610 30132 19616 30184
rect 19668 30172 19674 30184
rect 20088 30172 20116 30280
rect 20438 30268 20444 30280
rect 20496 30268 20502 30320
rect 22554 30268 22560 30320
rect 22612 30308 22618 30320
rect 24210 30308 24216 30320
rect 22612 30280 22692 30308
rect 24171 30280 24216 30308
rect 22612 30268 22618 30280
rect 20990 30240 20996 30252
rect 20951 30212 20996 30240
rect 20990 30200 20996 30212
rect 21048 30200 21054 30252
rect 22370 30249 22376 30252
rect 22364 30240 22376 30249
rect 22331 30212 22376 30240
rect 22364 30203 22376 30212
rect 22370 30200 22376 30203
rect 22428 30200 22434 30252
rect 22664 30240 22692 30280
rect 24210 30268 24216 30280
rect 24268 30268 24274 30320
rect 25777 30311 25835 30317
rect 25777 30277 25789 30311
rect 25823 30308 25835 30311
rect 26234 30308 26240 30320
rect 25823 30280 26240 30308
rect 25823 30277 25835 30280
rect 25777 30271 25835 30277
rect 26234 30268 26240 30280
rect 26292 30268 26298 30320
rect 29270 30308 29276 30320
rect 29231 30280 29276 30308
rect 29270 30268 29276 30280
rect 29328 30268 29334 30320
rect 31018 30308 31024 30320
rect 30979 30280 31024 30308
rect 31018 30268 31024 30280
rect 31076 30268 31082 30320
rect 31113 30311 31171 30317
rect 31113 30277 31125 30311
rect 31159 30308 31171 30311
rect 31202 30308 31208 30320
rect 31159 30280 31208 30308
rect 31159 30277 31171 30280
rect 31113 30271 31171 30277
rect 31202 30268 31208 30280
rect 31260 30268 31266 30320
rect 33134 30268 33140 30320
rect 33192 30308 33198 30320
rect 33698 30311 33756 30317
rect 33698 30308 33710 30311
rect 33192 30280 33710 30308
rect 33192 30268 33198 30280
rect 33698 30277 33710 30280
rect 33744 30277 33756 30311
rect 33698 30271 33756 30277
rect 35437 30311 35495 30317
rect 35437 30277 35449 30311
rect 35483 30308 35495 30311
rect 36354 30308 36360 30320
rect 35483 30280 36103 30308
rect 35483 30277 35495 30280
rect 35437 30271 35495 30277
rect 24121 30243 24179 30249
rect 24121 30240 24133 30243
rect 22664 30212 24133 30240
rect 24121 30209 24133 30212
rect 24167 30209 24179 30243
rect 24121 30203 24179 30209
rect 24305 30243 24363 30249
rect 24305 30209 24317 30243
rect 24351 30209 24363 30243
rect 24486 30240 24492 30252
rect 24447 30212 24492 30240
rect 24305 30203 24363 30209
rect 19668 30144 20116 30172
rect 19668 30132 19674 30144
rect 20254 30132 20260 30184
rect 20312 30172 20318 30184
rect 21269 30175 21327 30181
rect 21269 30172 21281 30175
rect 20312 30144 21281 30172
rect 20312 30132 20318 30144
rect 21269 30141 21281 30144
rect 21315 30141 21327 30175
rect 21269 30135 21327 30141
rect 22094 30132 22100 30184
rect 22152 30172 22158 30184
rect 22152 30144 22197 30172
rect 22152 30132 22158 30144
rect 23198 30132 23204 30184
rect 23256 30172 23262 30184
rect 24320 30172 24348 30203
rect 24486 30200 24492 30212
rect 24544 30200 24550 30252
rect 24946 30200 24952 30252
rect 25004 30240 25010 30252
rect 25133 30243 25191 30249
rect 25133 30240 25145 30243
rect 25004 30212 25145 30240
rect 25004 30200 25010 30212
rect 25133 30209 25145 30212
rect 25179 30209 25191 30243
rect 25314 30240 25320 30252
rect 25275 30212 25320 30240
rect 25133 30203 25191 30209
rect 25314 30200 25320 30212
rect 25372 30200 25378 30252
rect 25409 30243 25467 30249
rect 25409 30209 25421 30243
rect 25455 30209 25467 30243
rect 25409 30203 25467 30209
rect 23256 30144 24348 30172
rect 23256 30132 23262 30144
rect 24854 30132 24860 30184
rect 24912 30172 24918 30184
rect 25424 30172 25452 30203
rect 25498 30200 25504 30252
rect 25556 30240 25562 30252
rect 29089 30243 29147 30249
rect 25556 30212 26372 30240
rect 25556 30200 25562 30212
rect 24912 30144 25452 30172
rect 24912 30132 24918 30144
rect 25332 30116 25360 30144
rect 18012 30076 19564 30104
rect 18012 30064 18018 30076
rect 19702 30064 19708 30116
rect 19760 30104 19766 30116
rect 20622 30104 20628 30116
rect 19760 30076 20628 30104
rect 19760 30064 19766 30076
rect 20622 30064 20628 30076
rect 20680 30064 20686 30116
rect 23382 30064 23388 30116
rect 23440 30104 23446 30116
rect 23477 30107 23535 30113
rect 23477 30104 23489 30107
rect 23440 30076 23489 30104
rect 23440 30064 23446 30076
rect 23477 30073 23489 30076
rect 23523 30073 23535 30107
rect 23477 30067 23535 30073
rect 23768 30076 25268 30104
rect 16666 30036 16672 30048
rect 15120 30008 16672 30036
rect 16666 29996 16672 30008
rect 16724 29996 16730 30048
rect 17494 30036 17500 30048
rect 17455 30008 17500 30036
rect 17494 29996 17500 30008
rect 17552 29996 17558 30048
rect 20162 29996 20168 30048
rect 20220 30036 20226 30048
rect 20438 30036 20444 30048
rect 20220 30008 20444 30036
rect 20220 29996 20226 30008
rect 20438 29996 20444 30008
rect 20496 29996 20502 30048
rect 20806 29996 20812 30048
rect 20864 30036 20870 30048
rect 23768 30036 23796 30076
rect 20864 30008 23796 30036
rect 20864 29996 20870 30008
rect 23842 29996 23848 30048
rect 23900 30036 23906 30048
rect 23937 30039 23995 30045
rect 23937 30036 23949 30039
rect 23900 30008 23949 30036
rect 23900 29996 23906 30008
rect 23937 30005 23949 30008
rect 23983 30005 23995 30039
rect 25240 30036 25268 30076
rect 25314 30064 25320 30116
rect 25372 30064 25378 30116
rect 26344 30113 26372 30212
rect 29089 30209 29101 30243
rect 29135 30240 29147 30243
rect 29546 30240 29552 30252
rect 29135 30212 29552 30240
rect 29135 30209 29147 30212
rect 29089 30203 29147 30209
rect 29546 30200 29552 30212
rect 29604 30200 29610 30252
rect 30926 30240 30932 30252
rect 30887 30212 30932 30240
rect 30926 30200 30932 30212
rect 30984 30200 30990 30252
rect 31297 30243 31355 30249
rect 31297 30209 31309 30243
rect 31343 30240 31355 30243
rect 32030 30240 32036 30252
rect 31343 30212 32036 30240
rect 31343 30209 31355 30212
rect 31297 30203 31355 30209
rect 32030 30200 32036 30212
rect 32088 30200 32094 30252
rect 33410 30240 33416 30252
rect 32968 30212 33416 30240
rect 30944 30172 30972 30200
rect 32968 30172 32996 30212
rect 33410 30200 33416 30212
rect 33468 30200 33474 30252
rect 35069 30243 35127 30249
rect 35069 30209 35081 30243
rect 35115 30209 35127 30243
rect 35069 30203 35127 30209
rect 35253 30243 35311 30249
rect 35253 30209 35265 30243
rect 35299 30240 35311 30243
rect 35526 30240 35532 30252
rect 35299 30212 35532 30240
rect 35299 30209 35311 30212
rect 35253 30203 35311 30209
rect 30944 30144 32996 30172
rect 33965 30175 34023 30181
rect 33965 30141 33977 30175
rect 34011 30141 34023 30175
rect 35084 30172 35112 30203
rect 35526 30200 35532 30212
rect 35584 30200 35590 30252
rect 35894 30240 35900 30252
rect 35855 30212 35900 30240
rect 35894 30200 35900 30212
rect 35952 30200 35958 30252
rect 36075 30249 36103 30280
rect 36188 30280 36360 30308
rect 36188 30249 36216 30280
rect 36354 30268 36360 30280
rect 36412 30268 36418 30320
rect 36060 30243 36118 30249
rect 36060 30209 36072 30243
rect 36106 30209 36118 30243
rect 36060 30203 36118 30209
rect 36173 30243 36231 30249
rect 36173 30209 36185 30243
rect 36219 30209 36231 30243
rect 36173 30203 36231 30209
rect 36265 30243 36323 30249
rect 36265 30209 36277 30243
rect 36311 30209 36323 30243
rect 37277 30243 37335 30249
rect 37277 30240 37289 30243
rect 36265 30203 36323 30209
rect 36464 30212 37289 30240
rect 35158 30172 35164 30184
rect 35071 30144 35164 30172
rect 33965 30135 34023 30141
rect 26329 30107 26387 30113
rect 26329 30073 26341 30107
rect 26375 30104 26387 30107
rect 31202 30104 31208 30116
rect 26375 30076 31208 30104
rect 26375 30073 26387 30076
rect 26329 30067 26387 30073
rect 31202 30064 31208 30076
rect 31260 30064 31266 30116
rect 27798 30036 27804 30048
rect 25240 30008 27804 30036
rect 23937 29999 23995 30005
rect 27798 29996 27804 30008
rect 27856 29996 27862 30048
rect 28810 29996 28816 30048
rect 28868 30036 28874 30048
rect 28905 30039 28963 30045
rect 28905 30036 28917 30039
rect 28868 30008 28917 30036
rect 28868 29996 28874 30008
rect 28905 30005 28917 30008
rect 28951 30005 28963 30039
rect 28905 29999 28963 30005
rect 30745 30039 30803 30045
rect 30745 30005 30757 30039
rect 30791 30036 30803 30039
rect 31386 30036 31392 30048
rect 30791 30008 31392 30036
rect 30791 30005 30803 30008
rect 30745 29999 30803 30005
rect 31386 29996 31392 30008
rect 31444 29996 31450 30048
rect 32585 30039 32643 30045
rect 32585 30005 32597 30039
rect 32631 30036 32643 30039
rect 33226 30036 33232 30048
rect 32631 30008 33232 30036
rect 32631 30005 32643 30008
rect 32585 29999 32643 30005
rect 33226 29996 33232 30008
rect 33284 29996 33290 30048
rect 33980 30036 34008 30135
rect 35158 30132 35164 30144
rect 35216 30172 35222 30184
rect 35802 30172 35808 30184
rect 35216 30144 35808 30172
rect 35216 30132 35222 30144
rect 35802 30132 35808 30144
rect 35860 30132 35866 30184
rect 34238 30064 34244 30116
rect 34296 30104 34302 30116
rect 36280 30104 36308 30203
rect 36464 30172 36492 30212
rect 37277 30209 37289 30212
rect 37323 30209 37335 30243
rect 37277 30203 37335 30209
rect 36391 30144 36492 30172
rect 36391 30104 36419 30144
rect 37918 30104 37924 30116
rect 34296 30076 36419 30104
rect 36464 30076 37924 30104
rect 34296 30064 34302 30076
rect 36464 30036 36492 30076
rect 37918 30064 37924 30076
rect 37976 30064 37982 30116
rect 33980 30008 36492 30036
rect 36538 29996 36544 30048
rect 36596 30036 36602 30048
rect 36596 30008 36641 30036
rect 36596 29996 36602 30008
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 2866 29832 2872 29844
rect 2827 29804 2872 29832
rect 2866 29792 2872 29804
rect 2924 29792 2930 29844
rect 7926 29792 7932 29844
rect 7984 29832 7990 29844
rect 8110 29832 8116 29844
rect 7984 29804 8116 29832
rect 7984 29792 7990 29804
rect 8110 29792 8116 29804
rect 8168 29832 8174 29844
rect 8168 29804 10180 29832
rect 8168 29792 8174 29804
rect 10152 29764 10180 29804
rect 10226 29792 10232 29844
rect 10284 29832 10290 29844
rect 10962 29832 10968 29844
rect 10284 29804 10968 29832
rect 10284 29792 10290 29804
rect 10962 29792 10968 29804
rect 11020 29792 11026 29844
rect 11882 29832 11888 29844
rect 11843 29804 11888 29832
rect 11882 29792 11888 29804
rect 11940 29792 11946 29844
rect 18506 29792 18512 29844
rect 18564 29832 18570 29844
rect 19245 29835 19303 29841
rect 19245 29832 19257 29835
rect 18564 29804 19257 29832
rect 18564 29792 18570 29804
rect 19245 29801 19257 29804
rect 19291 29801 19303 29835
rect 19245 29795 19303 29801
rect 19334 29792 19340 29844
rect 19392 29832 19398 29844
rect 20165 29835 20223 29841
rect 20165 29832 20177 29835
rect 19392 29804 20177 29832
rect 19392 29792 19398 29804
rect 20165 29801 20177 29804
rect 20211 29801 20223 29835
rect 25498 29832 25504 29844
rect 20165 29795 20223 29801
rect 20272 29804 25504 29832
rect 13446 29764 13452 29776
rect 10152 29736 13452 29764
rect 13446 29724 13452 29736
rect 13504 29724 13510 29776
rect 15838 29764 15844 29776
rect 15751 29736 15844 29764
rect 15838 29724 15844 29736
rect 15896 29764 15902 29776
rect 17126 29764 17132 29776
rect 15896 29736 17132 29764
rect 15896 29724 15902 29736
rect 17126 29724 17132 29736
rect 17184 29764 17190 29776
rect 20272 29764 20300 29804
rect 25498 29792 25504 29804
rect 25556 29792 25562 29844
rect 27798 29832 27804 29844
rect 27759 29804 27804 29832
rect 27798 29792 27804 29804
rect 27856 29792 27862 29844
rect 29546 29832 29552 29844
rect 29507 29804 29552 29832
rect 29546 29792 29552 29804
rect 29604 29792 29610 29844
rect 31110 29832 31116 29844
rect 30024 29804 31116 29832
rect 17184 29736 20300 29764
rect 21269 29767 21327 29773
rect 17184 29724 17190 29736
rect 21269 29733 21281 29767
rect 21315 29764 21327 29767
rect 22462 29764 22468 29776
rect 21315 29736 22468 29764
rect 21315 29733 21327 29736
rect 21269 29727 21327 29733
rect 22462 29724 22468 29736
rect 22520 29724 22526 29776
rect 25038 29764 25044 29776
rect 22664 29736 25044 29764
rect 3234 29656 3240 29708
rect 3292 29696 3298 29708
rect 3292 29668 4660 29696
rect 3292 29656 3298 29668
rect 3602 29588 3608 29640
rect 3660 29628 3666 29640
rect 4632 29637 4660 29668
rect 8202 29656 8208 29708
rect 8260 29696 8266 29708
rect 9125 29699 9183 29705
rect 9125 29696 9137 29699
rect 8260 29668 9137 29696
rect 8260 29656 8266 29668
rect 9125 29665 9137 29668
rect 9171 29665 9183 29699
rect 9125 29659 9183 29665
rect 11333 29699 11391 29705
rect 11333 29665 11345 29699
rect 11379 29696 11391 29699
rect 11882 29696 11888 29708
rect 11379 29668 11888 29696
rect 11379 29665 11391 29668
rect 11333 29659 11391 29665
rect 11882 29656 11888 29668
rect 11940 29656 11946 29708
rect 19610 29696 19616 29708
rect 18064 29668 19616 29696
rect 4341 29631 4399 29637
rect 4341 29628 4353 29631
rect 3660 29600 4353 29628
rect 3660 29588 3666 29600
rect 4341 29597 4353 29600
rect 4387 29597 4399 29631
rect 4341 29591 4399 29597
rect 4617 29631 4675 29637
rect 4617 29597 4629 29631
rect 4663 29597 4675 29631
rect 4617 29591 4675 29597
rect 4706 29588 4712 29640
rect 4764 29628 4770 29640
rect 4764 29600 4809 29628
rect 4764 29588 4770 29600
rect 9214 29588 9220 29640
rect 9272 29628 9278 29640
rect 9381 29631 9439 29637
rect 9381 29628 9393 29631
rect 9272 29600 9393 29628
rect 9272 29588 9278 29600
rect 9381 29597 9393 29600
rect 9427 29597 9439 29631
rect 9381 29591 9439 29597
rect 10778 29588 10784 29640
rect 10836 29628 10842 29640
rect 11149 29631 11207 29637
rect 11149 29628 11161 29631
rect 10836 29600 11161 29628
rect 10836 29588 10842 29600
rect 11149 29597 11161 29600
rect 11195 29597 11207 29631
rect 11149 29591 11207 29597
rect 12250 29588 12256 29640
rect 12308 29628 12314 29640
rect 17494 29628 17500 29640
rect 12308 29600 17500 29628
rect 12308 29588 12314 29600
rect 17494 29588 17500 29600
rect 17552 29588 17558 29640
rect 17862 29588 17868 29640
rect 17920 29628 17926 29640
rect 18064 29637 18092 29668
rect 19610 29656 19616 29668
rect 19668 29656 19674 29708
rect 20714 29696 20720 29708
rect 20364 29668 20720 29696
rect 18049 29631 18107 29637
rect 18049 29628 18061 29631
rect 17920 29600 18061 29628
rect 17920 29588 17926 29600
rect 18049 29597 18061 29600
rect 18095 29597 18107 29631
rect 18049 29591 18107 29597
rect 19429 29631 19487 29637
rect 19429 29597 19441 29631
rect 19475 29628 19487 29631
rect 20070 29628 20076 29640
rect 19475 29600 20076 29628
rect 19475 29597 19487 29600
rect 19429 29591 19487 29597
rect 20070 29588 20076 29600
rect 20128 29588 20134 29640
rect 20364 29637 20392 29668
rect 20714 29656 20720 29668
rect 20772 29696 20778 29708
rect 22370 29696 22376 29708
rect 20772 29668 22376 29696
rect 20772 29656 20778 29668
rect 22370 29656 22376 29668
rect 22428 29656 22434 29708
rect 20349 29631 20407 29637
rect 20349 29597 20361 29631
rect 20395 29597 20407 29631
rect 22554 29628 22560 29640
rect 22515 29600 22560 29628
rect 20349 29591 20407 29597
rect 22554 29588 22560 29600
rect 22612 29588 22618 29640
rect 22664 29637 22692 29736
rect 25038 29724 25044 29736
rect 25096 29724 25102 29776
rect 30024 29764 30052 29804
rect 31110 29792 31116 29804
rect 31168 29792 31174 29844
rect 35526 29792 35532 29844
rect 35584 29832 35590 29844
rect 39301 29835 39359 29841
rect 39301 29832 39313 29835
rect 35584 29804 39313 29832
rect 35584 29792 35590 29804
rect 39301 29801 39313 29804
rect 39347 29801 39359 29835
rect 39301 29795 39359 29801
rect 28736 29736 30052 29764
rect 24946 29696 24952 29708
rect 24872 29668 24952 29696
rect 22649 29631 22707 29637
rect 22649 29597 22661 29631
rect 22695 29597 22707 29631
rect 22649 29591 22707 29597
rect 22925 29631 22983 29637
rect 22925 29597 22937 29631
rect 22971 29628 22983 29631
rect 23382 29628 23388 29640
rect 22971 29600 23388 29628
rect 22971 29597 22983 29600
rect 22925 29591 22983 29597
rect 23382 29588 23388 29600
rect 23440 29588 23446 29640
rect 23474 29588 23480 29640
rect 23532 29628 23538 29640
rect 24872 29637 24900 29668
rect 24946 29656 24952 29668
rect 25004 29656 25010 29708
rect 25314 29696 25320 29708
rect 25148 29668 25320 29696
rect 23845 29631 23903 29637
rect 23845 29628 23857 29631
rect 23532 29600 23857 29628
rect 23532 29588 23538 29600
rect 23845 29597 23857 29600
rect 23891 29597 23903 29631
rect 23845 29591 23903 29597
rect 24857 29631 24915 29637
rect 24857 29597 24869 29631
rect 24903 29597 24915 29631
rect 25038 29628 25044 29640
rect 24999 29600 25044 29628
rect 24857 29591 24915 29597
rect 25038 29588 25044 29600
rect 25096 29588 25102 29640
rect 25148 29637 25176 29668
rect 25314 29656 25320 29668
rect 25372 29656 25378 29708
rect 25133 29631 25191 29637
rect 25133 29597 25145 29631
rect 25179 29597 25191 29631
rect 25133 29591 25191 29597
rect 25225 29631 25283 29637
rect 25225 29597 25237 29631
rect 25271 29628 25283 29631
rect 25271 29600 27200 29628
rect 25271 29597 25283 29600
rect 25225 29591 25283 29597
rect 4525 29563 4583 29569
rect 4525 29529 4537 29563
rect 4571 29560 4583 29563
rect 4798 29560 4804 29572
rect 4571 29532 4804 29560
rect 4571 29529 4583 29532
rect 4525 29523 4583 29529
rect 4798 29520 4804 29532
rect 4856 29520 4862 29572
rect 10042 29560 10048 29572
rect 9955 29532 10048 29560
rect 9968 29504 9996 29532
rect 10042 29520 10048 29532
rect 10100 29560 10106 29572
rect 17954 29560 17960 29572
rect 10100 29532 11192 29560
rect 10100 29520 10106 29532
rect 4893 29495 4951 29501
rect 4893 29461 4905 29495
rect 4939 29492 4951 29495
rect 4982 29492 4988 29504
rect 4939 29464 4988 29492
rect 4939 29461 4951 29464
rect 4893 29455 4951 29461
rect 4982 29452 4988 29464
rect 5040 29452 5046 29504
rect 9950 29452 9956 29504
rect 10008 29452 10014 29504
rect 10505 29495 10563 29501
rect 10505 29461 10517 29495
rect 10551 29492 10563 29495
rect 11054 29492 11060 29504
rect 10551 29464 11060 29492
rect 10551 29461 10563 29464
rect 10505 29455 10563 29461
rect 11054 29452 11060 29464
rect 11112 29452 11118 29504
rect 11164 29492 11192 29532
rect 12406 29532 17960 29560
rect 12406 29492 12434 29532
rect 17954 29520 17960 29532
rect 18012 29520 18018 29572
rect 18233 29563 18291 29569
rect 18233 29529 18245 29563
rect 18279 29560 18291 29563
rect 18598 29560 18604 29572
rect 18279 29532 18604 29560
rect 18279 29529 18291 29532
rect 18233 29523 18291 29529
rect 18598 29520 18604 29532
rect 18656 29520 18662 29572
rect 19334 29520 19340 29572
rect 19392 29560 19398 29572
rect 19613 29563 19671 29569
rect 19613 29560 19625 29563
rect 19392 29532 19625 29560
rect 19392 29520 19398 29532
rect 19613 29529 19625 29532
rect 19659 29560 19671 29563
rect 20254 29560 20260 29572
rect 19659 29532 20260 29560
rect 19659 29529 19671 29532
rect 19613 29523 19671 29529
rect 20254 29520 20260 29532
rect 20312 29560 20318 29572
rect 20533 29563 20591 29569
rect 20533 29560 20545 29563
rect 20312 29532 20545 29560
rect 20312 29520 20318 29532
rect 20533 29529 20545 29532
rect 20579 29529 20591 29563
rect 20533 29523 20591 29529
rect 11164 29464 12434 29492
rect 16758 29452 16764 29504
rect 16816 29492 16822 29504
rect 16853 29495 16911 29501
rect 16853 29492 16865 29495
rect 16816 29464 16865 29492
rect 16816 29452 16822 29464
rect 16853 29461 16865 29464
rect 16899 29461 16911 29495
rect 16853 29455 16911 29461
rect 17034 29452 17040 29504
rect 17092 29492 17098 29504
rect 17402 29492 17408 29504
rect 17092 29464 17408 29492
rect 17092 29452 17098 29464
rect 17402 29452 17408 29464
rect 17460 29452 17466 29504
rect 20548 29492 20576 29523
rect 20622 29520 20628 29572
rect 20680 29560 20686 29572
rect 20898 29560 20904 29572
rect 20680 29532 20904 29560
rect 20680 29520 20686 29532
rect 20898 29520 20904 29532
rect 20956 29560 20962 29572
rect 21085 29563 21143 29569
rect 21085 29560 21097 29563
rect 20956 29532 21097 29560
rect 20956 29520 20962 29532
rect 21085 29529 21097 29532
rect 21131 29529 21143 29563
rect 21085 29523 21143 29529
rect 22741 29563 22799 29569
rect 22741 29529 22753 29563
rect 22787 29560 22799 29563
rect 23198 29560 23204 29572
rect 22787 29532 23204 29560
rect 22787 29529 22799 29532
rect 22741 29523 22799 29529
rect 23198 29520 23204 29532
rect 23256 29520 23262 29572
rect 24394 29520 24400 29572
rect 24452 29560 24458 29572
rect 25240 29560 25268 29591
rect 24452 29532 25268 29560
rect 25501 29563 25559 29569
rect 24452 29520 24458 29532
rect 25501 29529 25513 29563
rect 25547 29560 25559 29563
rect 27074 29563 27132 29569
rect 27074 29560 27086 29563
rect 25547 29532 27086 29560
rect 25547 29529 25559 29532
rect 25501 29523 25559 29529
rect 27074 29529 27086 29532
rect 27120 29529 27132 29563
rect 27172 29560 27200 29600
rect 27246 29588 27252 29640
rect 27304 29628 27310 29640
rect 27341 29631 27399 29637
rect 27341 29628 27353 29631
rect 27304 29600 27353 29628
rect 27304 29588 27310 29600
rect 27341 29597 27353 29600
rect 27387 29597 27399 29631
rect 27341 29591 27399 29597
rect 27798 29588 27804 29640
rect 27856 29628 27862 29640
rect 28626 29628 28632 29640
rect 27856 29600 28632 29628
rect 27856 29588 27862 29600
rect 28626 29588 28632 29600
rect 28684 29588 28690 29640
rect 28736 29637 28764 29736
rect 35342 29696 35348 29708
rect 33796 29668 35348 29696
rect 28721 29631 28779 29637
rect 28721 29597 28733 29631
rect 28767 29597 28779 29631
rect 28721 29591 28779 29597
rect 28810 29588 28816 29640
rect 28868 29628 28874 29640
rect 28997 29631 29055 29637
rect 28868 29600 28913 29628
rect 28868 29588 28874 29600
rect 28997 29597 29009 29631
rect 29043 29628 29055 29631
rect 29822 29628 29828 29640
rect 29043 29600 29828 29628
rect 29043 29597 29055 29600
rect 28997 29591 29055 29597
rect 29822 29588 29828 29600
rect 29880 29588 29886 29640
rect 30926 29628 30932 29640
rect 30887 29600 30932 29628
rect 30926 29588 30932 29600
rect 30984 29588 30990 29640
rect 33410 29588 33416 29640
rect 33468 29628 33474 29640
rect 33796 29637 33824 29668
rect 35342 29656 35348 29668
rect 35400 29656 35406 29708
rect 37918 29656 37924 29708
rect 37976 29705 37982 29708
rect 37976 29696 37986 29705
rect 37976 29668 38021 29696
rect 37976 29659 37986 29668
rect 37976 29656 37982 29659
rect 33689 29631 33747 29637
rect 33689 29628 33701 29631
rect 33468 29600 33701 29628
rect 33468 29588 33474 29600
rect 33689 29597 33701 29600
rect 33735 29597 33747 29631
rect 33689 29591 33747 29597
rect 33781 29631 33839 29637
rect 33781 29597 33793 29631
rect 33827 29597 33839 29631
rect 33781 29591 33839 29597
rect 34057 29631 34115 29637
rect 34057 29597 34069 29631
rect 34103 29628 34115 29631
rect 34422 29628 34428 29640
rect 34103 29600 34428 29628
rect 34103 29597 34115 29600
rect 34057 29591 34115 29597
rect 34422 29588 34428 29600
rect 34480 29588 34486 29640
rect 36538 29588 36544 29640
rect 36596 29628 36602 29640
rect 38177 29631 38235 29637
rect 38177 29628 38189 29631
rect 36596 29600 38189 29628
rect 36596 29588 36602 29600
rect 38177 29597 38189 29600
rect 38223 29597 38235 29631
rect 58158 29628 58164 29640
rect 58119 29600 58164 29628
rect 38177 29591 38235 29597
rect 58158 29588 58164 29600
rect 58216 29588 58222 29640
rect 28353 29563 28411 29569
rect 27172 29532 27936 29560
rect 27074 29523 27132 29529
rect 21729 29495 21787 29501
rect 21729 29492 21741 29495
rect 20548 29464 21741 29492
rect 21729 29461 21741 29464
rect 21775 29461 21787 29495
rect 21729 29455 21787 29461
rect 22373 29495 22431 29501
rect 22373 29461 22385 29495
rect 22419 29492 22431 29495
rect 22462 29492 22468 29504
rect 22419 29464 22468 29492
rect 22419 29461 22431 29464
rect 22373 29455 22431 29461
rect 22462 29452 22468 29464
rect 22520 29452 22526 29504
rect 23658 29492 23664 29504
rect 23619 29464 23664 29492
rect 23658 29452 23664 29464
rect 23716 29452 23722 29504
rect 24486 29452 24492 29504
rect 24544 29492 24550 29504
rect 25961 29495 26019 29501
rect 25961 29492 25973 29495
rect 24544 29464 25973 29492
rect 24544 29452 24550 29464
rect 25961 29461 25973 29464
rect 26007 29461 26019 29495
rect 27908 29492 27936 29532
rect 28353 29529 28365 29563
rect 28399 29560 28411 29563
rect 30662 29563 30720 29569
rect 30662 29560 30674 29563
rect 28399 29532 30674 29560
rect 28399 29529 28411 29532
rect 28353 29523 28411 29529
rect 30662 29529 30674 29532
rect 30708 29529 30720 29563
rect 30662 29523 30720 29529
rect 33594 29520 33600 29572
rect 33652 29560 33658 29572
rect 33870 29560 33876 29572
rect 33652 29532 33876 29560
rect 33652 29520 33658 29532
rect 33870 29520 33876 29532
rect 33928 29520 33934 29572
rect 35802 29560 35808 29572
rect 35763 29532 35808 29560
rect 35802 29520 35808 29532
rect 35860 29520 35866 29572
rect 35894 29520 35900 29572
rect 35952 29560 35958 29572
rect 35989 29563 36047 29569
rect 35989 29560 36001 29563
rect 35952 29532 36001 29560
rect 35952 29520 35958 29532
rect 35989 29529 36001 29532
rect 36035 29560 36047 29563
rect 36630 29560 36636 29572
rect 36035 29532 36636 29560
rect 36035 29529 36047 29532
rect 35989 29523 36047 29529
rect 36630 29520 36636 29532
rect 36688 29520 36694 29572
rect 31941 29495 31999 29501
rect 31941 29492 31953 29495
rect 27908 29464 31953 29492
rect 25961 29455 26019 29461
rect 31941 29461 31953 29464
rect 31987 29492 31999 29495
rect 33318 29492 33324 29504
rect 31987 29464 33324 29492
rect 31987 29461 31999 29464
rect 31941 29455 31999 29461
rect 33318 29452 33324 29464
rect 33376 29452 33382 29504
rect 33505 29495 33563 29501
rect 33505 29461 33517 29495
rect 33551 29492 33563 29495
rect 34330 29492 34336 29504
rect 33551 29464 34336 29492
rect 33551 29461 33563 29464
rect 33505 29455 33563 29461
rect 34330 29452 34336 29464
rect 34388 29452 34394 29504
rect 36078 29452 36084 29504
rect 36136 29492 36142 29504
rect 36173 29495 36231 29501
rect 36173 29492 36185 29495
rect 36136 29464 36185 29492
rect 36136 29452 36142 29464
rect 36173 29461 36185 29464
rect 36219 29461 36231 29495
rect 36173 29455 36231 29461
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 3697 29291 3755 29297
rect 3697 29257 3709 29291
rect 3743 29288 3755 29291
rect 4614 29288 4620 29300
rect 3743 29260 4620 29288
rect 3743 29257 3755 29260
rect 3697 29251 3755 29257
rect 3712 29220 3740 29251
rect 4614 29248 4620 29260
rect 4672 29248 4678 29300
rect 11606 29288 11612 29300
rect 7760 29260 11612 29288
rect 2772 29192 3740 29220
rect 2772 29161 2800 29192
rect 3970 29180 3976 29232
rect 4028 29220 4034 29232
rect 4525 29223 4583 29229
rect 4525 29220 4537 29223
rect 4028 29192 4537 29220
rect 4028 29180 4034 29192
rect 4525 29189 4537 29192
rect 4571 29189 4583 29223
rect 4706 29220 4712 29232
rect 4525 29183 4583 29189
rect 4632 29192 4712 29220
rect 2772 29155 2835 29161
rect 2772 29127 2789 29155
rect 2777 29121 2789 29127
rect 2823 29121 2835 29155
rect 2777 29115 2835 29121
rect 2869 29155 2927 29161
rect 2869 29121 2881 29155
rect 2915 29121 2927 29155
rect 2869 29115 2927 29121
rect 2682 29044 2688 29096
rect 2740 29084 2746 29096
rect 2884 29084 2912 29115
rect 2958 29112 2964 29164
rect 3016 29152 3022 29164
rect 3016 29124 3061 29152
rect 3016 29112 3022 29124
rect 3142 29112 3148 29164
rect 3200 29152 3206 29164
rect 3200 29124 3245 29152
rect 3200 29112 3206 29124
rect 3418 29112 3424 29164
rect 3476 29152 3482 29164
rect 4632 29161 4660 29192
rect 4706 29180 4712 29192
rect 4764 29220 4770 29232
rect 4764 29192 5212 29220
rect 4764 29180 4770 29192
rect 5184 29164 5212 29192
rect 4249 29155 4307 29161
rect 4249 29152 4261 29155
rect 3476 29124 4261 29152
rect 3476 29112 3482 29124
rect 4249 29121 4261 29124
rect 4295 29121 4307 29155
rect 4249 29115 4307 29121
rect 4433 29155 4491 29161
rect 4433 29121 4445 29155
rect 4479 29121 4491 29155
rect 4433 29115 4491 29121
rect 4617 29155 4675 29161
rect 4617 29121 4629 29155
rect 4663 29121 4675 29155
rect 4617 29115 4675 29121
rect 2740 29056 2912 29084
rect 4448 29084 4476 29115
rect 4798 29112 4804 29164
rect 4856 29112 4862 29164
rect 5166 29112 5172 29164
rect 5224 29152 5230 29164
rect 7653 29155 7711 29161
rect 7653 29152 7665 29155
rect 5224 29124 7665 29152
rect 5224 29112 5230 29124
rect 7653 29121 7665 29124
rect 7699 29152 7711 29155
rect 7760 29152 7788 29260
rect 11606 29248 11612 29260
rect 11664 29248 11670 29300
rect 12802 29288 12808 29300
rect 12763 29260 12808 29288
rect 12802 29248 12808 29260
rect 12860 29248 12866 29300
rect 15657 29291 15715 29297
rect 15657 29257 15669 29291
rect 15703 29288 15715 29291
rect 15838 29288 15844 29300
rect 15703 29260 15844 29288
rect 15703 29257 15715 29260
rect 15657 29251 15715 29257
rect 15838 29248 15844 29260
rect 15896 29288 15902 29300
rect 19886 29288 19892 29300
rect 15896 29260 19892 29288
rect 15896 29248 15902 29260
rect 19886 29248 19892 29260
rect 19944 29248 19950 29300
rect 20254 29288 20260 29300
rect 20180 29260 20260 29288
rect 7926 29220 7932 29232
rect 7887 29192 7932 29220
rect 7926 29180 7932 29192
rect 7984 29180 7990 29232
rect 9398 29180 9404 29232
rect 9456 29220 9462 29232
rect 9456 29192 9901 29220
rect 9456 29180 9462 29192
rect 9873 29164 9901 29192
rect 10594 29180 10600 29232
rect 10652 29220 10658 29232
rect 10781 29223 10839 29229
rect 10781 29220 10793 29223
rect 10652 29192 10793 29220
rect 10652 29180 10658 29192
rect 10781 29189 10793 29192
rect 10827 29189 10839 29223
rect 10962 29220 10968 29232
rect 10923 29192 10968 29220
rect 10781 29183 10839 29189
rect 10962 29180 10968 29192
rect 11020 29180 11026 29232
rect 11054 29180 11060 29232
rect 11112 29220 11118 29232
rect 13725 29223 13783 29229
rect 11112 29192 12572 29220
rect 11112 29180 11118 29192
rect 7699 29124 7788 29152
rect 7837 29155 7895 29161
rect 7699 29121 7711 29124
rect 7653 29115 7711 29121
rect 7837 29121 7849 29155
rect 7883 29152 7895 29155
rect 8202 29152 8208 29164
rect 7883 29124 8208 29152
rect 7883 29121 7895 29124
rect 7837 29115 7895 29121
rect 8202 29112 8208 29124
rect 8260 29112 8266 29164
rect 9769 29155 9827 29161
rect 9769 29121 9781 29155
rect 9815 29121 9827 29155
rect 9769 29115 9827 29121
rect 9858 29158 9916 29164
rect 9858 29124 9870 29158
rect 9904 29124 9916 29158
rect 9858 29118 9916 29124
rect 9953 29155 10011 29161
rect 9953 29121 9965 29155
rect 9999 29121 10011 29155
rect 9953 29115 10011 29121
rect 10137 29155 10195 29161
rect 10137 29121 10149 29155
rect 10183 29152 10195 29155
rect 10870 29152 10876 29164
rect 10183 29124 10876 29152
rect 10183 29121 10195 29124
rect 10137 29115 10195 29121
rect 4816 29084 4844 29112
rect 4448 29056 4844 29084
rect 9033 29087 9091 29093
rect 2740 29044 2746 29056
rect 9033 29053 9045 29087
rect 9079 29084 9091 29087
rect 9784 29084 9812 29115
rect 9968 29084 9996 29115
rect 10870 29112 10876 29124
rect 10928 29152 10934 29164
rect 12544 29152 12572 29192
rect 12820 29192 13492 29220
rect 12820 29152 12848 29192
rect 13354 29152 13360 29164
rect 10928 29124 11008 29152
rect 12544 29124 12848 29152
rect 13315 29124 13360 29152
rect 10928 29112 10934 29124
rect 10597 29087 10655 29093
rect 10597 29084 10609 29087
rect 9079 29056 9904 29084
rect 9968 29056 10609 29084
rect 9079 29053 9091 29056
rect 9033 29047 9091 29053
rect 3510 28976 3516 29028
rect 3568 29016 3574 29028
rect 4706 29016 4712 29028
rect 3568 28988 4712 29016
rect 3568 28976 3574 28988
rect 4706 28976 4712 28988
rect 4764 28976 4770 29028
rect 4801 29019 4859 29025
rect 4801 28985 4813 29019
rect 4847 29016 4859 29019
rect 4890 29016 4896 29028
rect 4847 28988 4896 29016
rect 4847 28985 4859 28988
rect 4801 28979 4859 28985
rect 4890 28976 4896 28988
rect 4948 28976 4954 29028
rect 9876 29016 9904 29056
rect 10597 29053 10609 29056
rect 10643 29053 10655 29087
rect 10597 29047 10655 29053
rect 10980 29028 11008 29124
rect 13354 29112 13360 29124
rect 13412 29112 13418 29164
rect 13464 29161 13492 29192
rect 13725 29189 13737 29223
rect 13771 29220 13783 29223
rect 14366 29220 14372 29232
rect 13771 29192 14372 29220
rect 13771 29189 13783 29192
rect 13725 29183 13783 29189
rect 14366 29180 14372 29192
rect 14424 29220 14430 29232
rect 14829 29223 14887 29229
rect 14829 29220 14841 29223
rect 14424 29192 14841 29220
rect 14424 29180 14430 29192
rect 14829 29189 14841 29192
rect 14875 29189 14887 29223
rect 17862 29220 17868 29232
rect 17823 29192 17868 29220
rect 14829 29183 14887 29189
rect 17862 29180 17868 29192
rect 17920 29180 17926 29232
rect 17954 29180 17960 29232
rect 18012 29220 18018 29232
rect 18785 29223 18843 29229
rect 18785 29220 18797 29223
rect 18012 29192 18797 29220
rect 18012 29180 18018 29192
rect 18785 29189 18797 29192
rect 18831 29189 18843 29223
rect 20070 29220 20076 29232
rect 20031 29192 20076 29220
rect 18785 29183 18843 29189
rect 20070 29180 20076 29192
rect 20128 29180 20134 29232
rect 13450 29155 13508 29161
rect 13450 29121 13462 29155
rect 13496 29121 13508 29155
rect 13450 29115 13508 29121
rect 13633 29155 13691 29161
rect 13633 29121 13645 29155
rect 13679 29121 13691 29155
rect 13633 29115 13691 29121
rect 11698 29044 11704 29096
rect 11756 29084 11762 29096
rect 13648 29084 13676 29115
rect 13814 29112 13820 29164
rect 13872 29161 13878 29164
rect 13872 29152 13880 29161
rect 13872 29124 13917 29152
rect 13872 29115 13880 29124
rect 13872 29112 13878 29115
rect 14274 29112 14280 29164
rect 14332 29152 14338 29164
rect 14645 29155 14703 29161
rect 14645 29152 14657 29155
rect 14332 29124 14657 29152
rect 14332 29112 14338 29124
rect 14645 29121 14657 29124
rect 14691 29121 14703 29155
rect 14645 29115 14703 29121
rect 19889 29155 19947 29161
rect 19889 29121 19901 29155
rect 19935 29152 19947 29155
rect 19978 29152 19984 29164
rect 19935 29124 19984 29152
rect 19935 29121 19947 29124
rect 19889 29115 19947 29121
rect 19978 29112 19984 29124
rect 20036 29112 20042 29164
rect 20180 29161 20208 29260
rect 20254 29248 20260 29260
rect 20312 29248 20318 29300
rect 23750 29248 23756 29300
rect 23808 29288 23814 29300
rect 23845 29291 23903 29297
rect 23845 29288 23857 29291
rect 23808 29260 23857 29288
rect 23808 29248 23814 29260
rect 23845 29257 23857 29260
rect 23891 29288 23903 29291
rect 24394 29288 24400 29300
rect 23891 29260 24400 29288
rect 23891 29257 23903 29260
rect 23845 29251 23903 29257
rect 24394 29248 24400 29260
rect 24452 29248 24458 29300
rect 24673 29291 24731 29297
rect 24673 29257 24685 29291
rect 24719 29288 24731 29291
rect 25038 29288 25044 29300
rect 24719 29260 25044 29288
rect 24719 29257 24731 29260
rect 24673 29251 24731 29257
rect 25038 29248 25044 29260
rect 25096 29248 25102 29300
rect 25222 29248 25228 29300
rect 25280 29288 25286 29300
rect 25590 29288 25596 29300
rect 25280 29260 25596 29288
rect 25280 29248 25286 29260
rect 25590 29248 25596 29260
rect 25648 29248 25654 29300
rect 25866 29248 25872 29300
rect 25924 29288 25930 29300
rect 25961 29291 26019 29297
rect 25961 29288 25973 29291
rect 25924 29260 25973 29288
rect 25924 29248 25930 29260
rect 25961 29257 25973 29260
rect 26007 29257 26019 29291
rect 25961 29251 26019 29257
rect 29546 29248 29552 29300
rect 29604 29248 29610 29300
rect 30561 29291 30619 29297
rect 30561 29257 30573 29291
rect 30607 29288 30619 29291
rect 32306 29288 32312 29300
rect 30607 29260 32312 29288
rect 30607 29257 30619 29260
rect 30561 29251 30619 29257
rect 32306 29248 32312 29260
rect 32364 29248 32370 29300
rect 35526 29288 35532 29300
rect 33796 29260 35532 29288
rect 21910 29180 21916 29232
rect 21968 29220 21974 29232
rect 22097 29223 22155 29229
rect 22097 29220 22109 29223
rect 21968 29192 22109 29220
rect 21968 29180 21974 29192
rect 22097 29189 22109 29192
rect 22143 29189 22155 29223
rect 22097 29183 22155 29189
rect 22186 29180 22192 29232
rect 22244 29220 22250 29232
rect 24486 29220 24492 29232
rect 22244 29192 22968 29220
rect 24447 29192 24492 29220
rect 22244 29180 22250 29192
rect 20161 29155 20219 29161
rect 20161 29121 20173 29155
rect 20207 29121 20219 29155
rect 20161 29115 20219 29121
rect 20257 29155 20315 29161
rect 20257 29121 20269 29155
rect 20303 29121 20315 29155
rect 20257 29115 20315 29121
rect 22005 29155 22063 29161
rect 22005 29121 22017 29155
rect 22051 29121 22063 29155
rect 22370 29152 22376 29164
rect 22331 29124 22376 29152
rect 22005 29115 22063 29121
rect 15378 29084 15384 29096
rect 11756 29056 15384 29084
rect 11756 29044 11762 29056
rect 15378 29044 15384 29056
rect 15436 29044 15442 29096
rect 20272 29084 20300 29115
rect 22020 29084 22048 29115
rect 22370 29112 22376 29124
rect 22428 29112 22434 29164
rect 22940 29161 22968 29192
rect 24486 29180 24492 29192
rect 24544 29180 24550 29232
rect 29454 29220 29460 29232
rect 29415 29192 29460 29220
rect 29454 29180 29460 29192
rect 29512 29180 29518 29232
rect 29564 29220 29592 29248
rect 30742 29220 30748 29232
rect 29564 29192 29776 29220
rect 22925 29155 22983 29161
rect 22925 29121 22937 29155
rect 22971 29152 22983 29155
rect 23198 29152 23204 29164
rect 22971 29124 23204 29152
rect 22971 29121 22983 29124
rect 22925 29115 22983 29121
rect 23198 29112 23204 29124
rect 23256 29112 23262 29164
rect 24302 29152 24308 29164
rect 24263 29124 24308 29152
rect 24302 29112 24308 29124
rect 24360 29152 24366 29164
rect 24578 29152 24584 29164
rect 24360 29124 24584 29152
rect 24360 29112 24366 29124
rect 24578 29112 24584 29124
rect 24636 29112 24642 29164
rect 25406 29152 25412 29164
rect 25367 29124 25412 29152
rect 25406 29112 25412 29124
rect 25464 29112 25470 29164
rect 26142 29152 26148 29164
rect 26103 29124 26148 29152
rect 26142 29112 26148 29124
rect 26200 29152 26206 29164
rect 26973 29155 27031 29161
rect 26973 29152 26985 29155
rect 26200 29124 26985 29152
rect 26200 29112 26206 29124
rect 26973 29121 26985 29124
rect 27019 29152 27031 29155
rect 27338 29152 27344 29164
rect 27019 29124 27344 29152
rect 27019 29121 27031 29124
rect 26973 29115 27031 29121
rect 27338 29112 27344 29124
rect 27396 29112 27402 29164
rect 29362 29152 29368 29164
rect 29323 29124 29368 29152
rect 29362 29112 29368 29124
rect 29420 29112 29426 29164
rect 29748 29161 29776 29192
rect 30392 29192 30748 29220
rect 30392 29161 30420 29192
rect 30742 29180 30748 29192
rect 30800 29180 30806 29232
rect 33796 29229 33824 29260
rect 35526 29248 35532 29260
rect 35584 29248 35590 29300
rect 36446 29288 36452 29300
rect 36407 29260 36452 29288
rect 36446 29248 36452 29260
rect 36504 29248 36510 29300
rect 36630 29248 36636 29300
rect 36688 29288 36694 29300
rect 39301 29291 39359 29297
rect 39301 29288 39313 29291
rect 36688 29260 39313 29288
rect 36688 29248 36694 29260
rect 39301 29257 39313 29260
rect 39347 29257 39359 29291
rect 39301 29251 39359 29257
rect 33781 29223 33839 29229
rect 33781 29189 33793 29223
rect 33827 29189 33839 29223
rect 33781 29183 33839 29189
rect 33870 29180 33876 29232
rect 33928 29220 33934 29232
rect 34606 29220 34612 29232
rect 33928 29192 33973 29220
rect 34072 29192 34612 29220
rect 33928 29180 33934 29192
rect 29549 29155 29607 29161
rect 29549 29121 29561 29155
rect 29595 29121 29607 29155
rect 29549 29115 29607 29121
rect 29733 29155 29791 29161
rect 29733 29121 29745 29155
rect 29779 29121 29791 29155
rect 29733 29115 29791 29121
rect 30377 29155 30435 29161
rect 30377 29121 30389 29155
rect 30423 29121 30435 29155
rect 30377 29115 30435 29121
rect 22554 29084 22560 29096
rect 20272 29056 22560 29084
rect 20272 29028 20300 29056
rect 22554 29044 22560 29056
rect 22612 29044 22618 29096
rect 23658 29044 23664 29096
rect 23716 29084 23722 29096
rect 29564 29084 29592 29115
rect 30392 29084 30420 29115
rect 30466 29112 30472 29164
rect 30524 29152 30530 29164
rect 30561 29155 30619 29161
rect 30561 29152 30573 29155
rect 30524 29124 30573 29152
rect 30524 29112 30530 29124
rect 30561 29121 30573 29124
rect 30607 29152 30619 29155
rect 31021 29155 31079 29161
rect 31021 29152 31033 29155
rect 30607 29124 31033 29152
rect 30607 29121 30619 29124
rect 30561 29115 30619 29121
rect 31021 29121 31033 29124
rect 31067 29121 31079 29155
rect 31021 29115 31079 29121
rect 33410 29112 33416 29164
rect 33468 29152 33474 29164
rect 34072 29161 34100 29192
rect 34606 29180 34612 29192
rect 34664 29180 34670 29232
rect 38562 29180 38568 29232
rect 38620 29220 38626 29232
rect 38746 29220 38752 29232
rect 38620 29192 38752 29220
rect 38620 29180 38626 29192
rect 38746 29180 38752 29192
rect 38804 29180 38810 29232
rect 33689 29155 33747 29161
rect 33689 29152 33701 29155
rect 33468 29124 33701 29152
rect 33468 29112 33474 29124
rect 33689 29121 33701 29124
rect 33735 29121 33747 29155
rect 33689 29115 33747 29121
rect 34057 29155 34115 29161
rect 34057 29121 34069 29155
rect 34103 29121 34115 29155
rect 34514 29152 34520 29164
rect 34475 29124 34520 29152
rect 34057 29115 34115 29121
rect 34514 29112 34520 29124
rect 34572 29112 34578 29164
rect 38010 29112 38016 29164
rect 38068 29152 38074 29164
rect 38177 29155 38235 29161
rect 38177 29152 38189 29155
rect 38068 29124 38189 29152
rect 38068 29112 38074 29124
rect 38177 29121 38189 29124
rect 38223 29121 38235 29155
rect 38177 29115 38235 29121
rect 34238 29084 34244 29096
rect 23716 29056 29500 29084
rect 29564 29056 30420 29084
rect 30852 29056 34244 29084
rect 23716 29044 23722 29056
rect 9950 29016 9956 29028
rect 9876 28988 9956 29016
rect 9950 28976 9956 28988
rect 10008 28976 10014 29028
rect 10962 28976 10968 29028
rect 11020 29016 11026 29028
rect 11517 29019 11575 29025
rect 11517 29016 11529 29019
rect 11020 28988 11529 29016
rect 11020 28976 11026 28988
rect 11517 28985 11529 28988
rect 11563 28985 11575 29019
rect 11517 28979 11575 28985
rect 14001 29019 14059 29025
rect 14001 28985 14013 29019
rect 14047 29016 14059 29019
rect 14918 29016 14924 29028
rect 14047 28988 14924 29016
rect 14047 28985 14059 28988
rect 14001 28979 14059 28985
rect 14918 28976 14924 28988
rect 14976 28976 14982 29028
rect 16114 28976 16120 29028
rect 16172 29016 16178 29028
rect 19334 29016 19340 29028
rect 16172 28988 19340 29016
rect 16172 28976 16178 28988
rect 19334 28976 19340 28988
rect 19392 28976 19398 29028
rect 20254 28976 20260 29028
rect 20312 28976 20318 29028
rect 20441 29019 20499 29025
rect 20441 28985 20453 29019
rect 20487 29016 20499 29019
rect 20530 29016 20536 29028
rect 20487 28988 20536 29016
rect 20487 28985 20499 28988
rect 20441 28979 20499 28985
rect 20530 28976 20536 28988
rect 20588 28976 20594 29028
rect 23106 29016 23112 29028
rect 23067 28988 23112 29016
rect 23106 28976 23112 28988
rect 23164 28976 23170 29028
rect 29178 29016 29184 29028
rect 29139 28988 29184 29016
rect 29178 28976 29184 28988
rect 29236 28976 29242 29028
rect 29472 29016 29500 29056
rect 30852 29016 30880 29056
rect 34238 29044 34244 29056
rect 34296 29044 34302 29096
rect 35161 29087 35219 29093
rect 35161 29084 35173 29087
rect 34624 29056 35173 29084
rect 29472 28988 30880 29016
rect 30944 28988 31156 29016
rect 2498 28948 2504 28960
rect 2459 28920 2504 28948
rect 2498 28908 2504 28920
rect 2556 28908 2562 28960
rect 8202 28908 8208 28960
rect 8260 28948 8266 28960
rect 8389 28951 8447 28957
rect 8389 28948 8401 28951
rect 8260 28920 8401 28948
rect 8260 28908 8266 28920
rect 8389 28917 8401 28920
rect 8435 28917 8447 28951
rect 9490 28948 9496 28960
rect 9451 28920 9496 28948
rect 8389 28911 8447 28917
rect 9490 28908 9496 28920
rect 9548 28908 9554 28960
rect 14826 28908 14832 28960
rect 14884 28948 14890 28960
rect 15013 28951 15071 28957
rect 15013 28948 15025 28951
rect 14884 28920 15025 28948
rect 14884 28908 14890 28920
rect 15013 28917 15025 28920
rect 15059 28917 15071 28951
rect 20898 28948 20904 28960
rect 20859 28920 20904 28948
rect 15013 28911 15071 28917
rect 20898 28908 20904 28920
rect 20956 28908 20962 28960
rect 21818 28948 21824 28960
rect 21779 28920 21824 28948
rect 21818 28908 21824 28920
rect 21876 28908 21882 28960
rect 30098 28908 30104 28960
rect 30156 28948 30162 28960
rect 30944 28948 30972 28988
rect 30156 28920 30972 28948
rect 31128 28948 31156 28988
rect 31202 28976 31208 29028
rect 31260 29016 31266 29028
rect 32582 29016 32588 29028
rect 31260 28988 32588 29016
rect 31260 28976 31266 28988
rect 32582 28976 32588 28988
rect 32640 28976 32646 29028
rect 33502 29016 33508 29028
rect 33463 28988 33508 29016
rect 33502 28976 33508 28988
rect 33560 28976 33566 29028
rect 34624 29016 34652 29056
rect 35161 29053 35173 29056
rect 35207 29053 35219 29087
rect 35161 29047 35219 29053
rect 35437 29087 35495 29093
rect 35437 29053 35449 29087
rect 35483 29084 35495 29087
rect 36262 29084 36268 29096
rect 35483 29056 36268 29084
rect 35483 29053 35495 29056
rect 35437 29047 35495 29053
rect 36262 29044 36268 29056
rect 36320 29044 36326 29096
rect 37918 29084 37924 29096
rect 37879 29056 37924 29084
rect 37918 29044 37924 29056
rect 37976 29044 37982 29096
rect 34440 28988 34652 29016
rect 34701 29019 34759 29025
rect 34238 28948 34244 28960
rect 31128 28920 34244 28948
rect 30156 28908 30162 28920
rect 34238 28908 34244 28920
rect 34296 28948 34302 28960
rect 34440 28948 34468 28988
rect 34701 28985 34713 29019
rect 34747 29016 34759 29019
rect 35802 29016 35808 29028
rect 34747 28988 35808 29016
rect 34747 28985 34759 28988
rect 34701 28979 34759 28985
rect 35802 28976 35808 28988
rect 35860 28976 35866 29028
rect 34296 28920 34468 28948
rect 34296 28908 34302 28920
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 2958 28744 2964 28756
rect 2919 28716 2964 28744
rect 2958 28704 2964 28716
rect 3016 28704 3022 28756
rect 8570 28704 8576 28756
rect 8628 28744 8634 28756
rect 15562 28744 15568 28756
rect 8628 28716 15568 28744
rect 8628 28704 8634 28716
rect 12802 28636 12808 28688
rect 12860 28676 12866 28688
rect 12860 28648 13584 28676
rect 12860 28636 12866 28648
rect 12437 28611 12495 28617
rect 12437 28577 12449 28611
rect 12483 28608 12495 28611
rect 12483 28580 13400 28608
rect 12483 28577 12495 28580
rect 12437 28571 12495 28577
rect 2593 28543 2651 28549
rect 2593 28509 2605 28543
rect 2639 28540 2651 28543
rect 3326 28540 3332 28552
rect 2639 28512 3332 28540
rect 2639 28509 2651 28512
rect 2593 28503 2651 28509
rect 3326 28500 3332 28512
rect 3384 28500 3390 28552
rect 4617 28543 4675 28549
rect 4617 28509 4629 28543
rect 4663 28509 4675 28543
rect 4617 28503 4675 28509
rect 2777 28475 2835 28481
rect 2777 28441 2789 28475
rect 2823 28472 2835 28475
rect 3786 28472 3792 28484
rect 2823 28444 3792 28472
rect 2823 28441 2835 28444
rect 2777 28435 2835 28441
rect 3786 28432 3792 28444
rect 3844 28472 3850 28484
rect 4632 28472 4660 28503
rect 4706 28500 4712 28552
rect 4764 28540 4770 28552
rect 4893 28543 4951 28549
rect 4893 28540 4905 28543
rect 4764 28512 4905 28540
rect 4764 28500 4770 28512
rect 4893 28509 4905 28512
rect 4939 28509 4951 28543
rect 4893 28503 4951 28509
rect 4985 28543 5043 28549
rect 4985 28509 4997 28543
rect 5031 28540 5043 28543
rect 5166 28540 5172 28552
rect 5031 28512 5172 28540
rect 5031 28509 5043 28512
rect 4985 28503 5043 28509
rect 5166 28500 5172 28512
rect 5224 28500 5230 28552
rect 9217 28543 9275 28549
rect 9217 28509 9229 28543
rect 9263 28540 9275 28543
rect 9306 28540 9312 28552
rect 9263 28512 9312 28540
rect 9263 28509 9275 28512
rect 9217 28503 9275 28509
rect 9306 28500 9312 28512
rect 9364 28500 9370 28552
rect 9490 28549 9496 28552
rect 9484 28540 9496 28549
rect 9451 28512 9496 28540
rect 9484 28503 9496 28512
rect 9490 28500 9496 28503
rect 9548 28500 9554 28552
rect 12069 28543 12127 28549
rect 12069 28509 12081 28543
rect 12115 28540 12127 28543
rect 12526 28540 12532 28552
rect 12115 28512 12532 28540
rect 12115 28509 12127 28512
rect 12069 28503 12127 28509
rect 12526 28500 12532 28512
rect 12584 28540 12590 28552
rect 12986 28540 12992 28552
rect 12584 28512 12992 28540
rect 12584 28500 12590 28512
rect 12986 28500 12992 28512
rect 13044 28500 13050 28552
rect 13372 28549 13400 28580
rect 13556 28549 13584 28648
rect 13173 28543 13231 28549
rect 13173 28509 13185 28543
rect 13219 28509 13231 28543
rect 13173 28503 13231 28509
rect 13265 28543 13323 28549
rect 13265 28509 13277 28543
rect 13311 28509 13323 28543
rect 13265 28503 13323 28509
rect 13357 28543 13415 28549
rect 13357 28509 13369 28543
rect 13403 28509 13415 28543
rect 13357 28503 13415 28509
rect 13541 28543 13599 28549
rect 13541 28509 13553 28543
rect 13587 28509 13599 28543
rect 13541 28503 13599 28509
rect 3844 28444 4660 28472
rect 3844 28432 3850 28444
rect 4798 28432 4804 28484
rect 4856 28472 4862 28484
rect 9766 28472 9772 28484
rect 4856 28444 9772 28472
rect 4856 28432 4862 28444
rect 9766 28432 9772 28444
rect 9824 28432 9830 28484
rect 12253 28475 12311 28481
rect 12253 28441 12265 28475
rect 12299 28472 12311 28475
rect 12434 28472 12440 28484
rect 12299 28444 12440 28472
rect 12299 28441 12311 28444
rect 12253 28435 12311 28441
rect 12434 28432 12440 28444
rect 12492 28432 12498 28484
rect 5169 28407 5227 28413
rect 5169 28373 5181 28407
rect 5215 28404 5227 28407
rect 6362 28404 6368 28416
rect 5215 28376 6368 28404
rect 5215 28373 5227 28376
rect 5169 28367 5227 28373
rect 6362 28364 6368 28376
rect 6420 28364 6426 28416
rect 9674 28364 9680 28416
rect 9732 28404 9738 28416
rect 10042 28404 10048 28416
rect 9732 28376 10048 28404
rect 9732 28364 9738 28376
rect 10042 28364 10048 28376
rect 10100 28364 10106 28416
rect 10594 28404 10600 28416
rect 10555 28376 10600 28404
rect 10594 28364 10600 28376
rect 10652 28364 10658 28416
rect 12894 28404 12900 28416
rect 12855 28376 12900 28404
rect 12894 28364 12900 28376
rect 12952 28364 12958 28416
rect 13188 28404 13216 28503
rect 13280 28472 13308 28503
rect 14550 28500 14556 28552
rect 14608 28540 14614 28552
rect 14645 28543 14703 28549
rect 14645 28540 14657 28543
rect 14608 28512 14657 28540
rect 14608 28500 14614 28512
rect 14645 28509 14657 28512
rect 14691 28509 14703 28543
rect 14826 28540 14832 28552
rect 14787 28512 14832 28540
rect 14645 28503 14703 28509
rect 14826 28500 14832 28512
rect 14884 28500 14890 28552
rect 14936 28549 14964 28716
rect 15562 28704 15568 28716
rect 15620 28704 15626 28756
rect 26786 28704 26792 28756
rect 26844 28744 26850 28756
rect 26881 28747 26939 28753
rect 26881 28744 26893 28747
rect 26844 28716 26893 28744
rect 26844 28704 26850 28716
rect 26881 28713 26893 28716
rect 26927 28713 26939 28747
rect 26881 28707 26939 28713
rect 29641 28747 29699 28753
rect 29641 28713 29653 28747
rect 29687 28744 29699 28747
rect 30098 28744 30104 28756
rect 29687 28716 30104 28744
rect 29687 28713 29699 28716
rect 29641 28707 29699 28713
rect 30098 28704 30104 28716
rect 30156 28704 30162 28756
rect 35802 28704 35808 28756
rect 35860 28744 35866 28756
rect 36633 28747 36691 28753
rect 35860 28716 36387 28744
rect 35860 28704 35866 28716
rect 16025 28679 16083 28685
rect 16025 28645 16037 28679
rect 16071 28676 16083 28679
rect 16850 28676 16856 28688
rect 16071 28648 16856 28676
rect 16071 28645 16083 28648
rect 16025 28639 16083 28645
rect 16850 28636 16856 28648
rect 16908 28636 16914 28688
rect 24581 28679 24639 28685
rect 24581 28645 24593 28679
rect 24627 28676 24639 28679
rect 24762 28676 24768 28688
rect 24627 28648 24768 28676
rect 24627 28645 24639 28648
rect 24581 28639 24639 28645
rect 24762 28636 24768 28648
rect 24820 28676 24826 28688
rect 35526 28676 35532 28688
rect 24820 28648 35532 28676
rect 24820 28636 24826 28648
rect 35526 28636 35532 28648
rect 35584 28636 35590 28688
rect 36262 28636 36268 28688
rect 36320 28636 36326 28688
rect 36359 28676 36387 28716
rect 36633 28713 36645 28747
rect 36679 28744 36691 28747
rect 38010 28744 38016 28756
rect 36679 28716 38016 28744
rect 36679 28713 36691 28716
rect 36633 28707 36691 28713
rect 38010 28704 38016 28716
rect 38068 28704 38074 28756
rect 36359 28648 37136 28676
rect 23750 28608 23756 28620
rect 15028 28580 23756 28608
rect 15028 28549 15056 28580
rect 23750 28568 23756 28580
rect 23808 28568 23814 28620
rect 30742 28608 30748 28620
rect 30703 28580 30748 28608
rect 30742 28568 30748 28580
rect 30800 28568 30806 28620
rect 33410 28568 33416 28620
rect 33468 28608 33474 28620
rect 33505 28611 33563 28617
rect 33505 28608 33517 28611
rect 33468 28580 33517 28608
rect 33468 28568 33474 28580
rect 33505 28577 33517 28580
rect 33551 28577 33563 28611
rect 35894 28608 35900 28620
rect 33505 28571 33563 28577
rect 34992 28580 35900 28608
rect 14921 28543 14979 28549
rect 14921 28509 14933 28543
rect 14967 28509 14979 28543
rect 14921 28503 14979 28509
rect 15013 28543 15071 28549
rect 15013 28509 15025 28543
rect 15059 28509 15071 28543
rect 15838 28540 15844 28552
rect 15799 28512 15844 28540
rect 15013 28503 15071 28509
rect 13446 28472 13452 28484
rect 13280 28444 13452 28472
rect 13446 28432 13452 28444
rect 13504 28432 13510 28484
rect 13906 28432 13912 28484
rect 13964 28472 13970 28484
rect 14185 28475 14243 28481
rect 14185 28472 14197 28475
rect 13964 28444 14197 28472
rect 13964 28432 13970 28444
rect 14185 28441 14197 28444
rect 14231 28472 14243 28475
rect 15028 28472 15056 28503
rect 15838 28500 15844 28512
rect 15896 28500 15902 28552
rect 24397 28543 24455 28549
rect 24397 28509 24409 28543
rect 24443 28540 24455 28543
rect 24854 28540 24860 28552
rect 24443 28512 24860 28540
rect 24443 28509 24455 28512
rect 24397 28503 24455 28509
rect 24854 28500 24860 28512
rect 24912 28500 24918 28552
rect 26237 28543 26295 28549
rect 26237 28540 26249 28543
rect 25148 28512 26249 28540
rect 14231 28444 15056 28472
rect 14231 28441 14243 28444
rect 14185 28435 14243 28441
rect 15194 28432 15200 28484
rect 15252 28472 15258 28484
rect 17497 28475 17555 28481
rect 17497 28472 17509 28475
rect 15252 28444 17509 28472
rect 15252 28432 15258 28444
rect 17497 28441 17509 28444
rect 17543 28472 17555 28475
rect 18049 28475 18107 28481
rect 18049 28472 18061 28475
rect 17543 28444 18061 28472
rect 17543 28441 17555 28444
rect 17497 28435 17555 28441
rect 18049 28441 18061 28444
rect 18095 28472 18107 28475
rect 20714 28472 20720 28484
rect 18095 28444 20720 28472
rect 18095 28441 18107 28444
rect 18049 28435 18107 28441
rect 20714 28432 20720 28444
rect 20772 28432 20778 28484
rect 23474 28472 23480 28484
rect 23387 28444 23480 28472
rect 23474 28432 23480 28444
rect 23532 28472 23538 28484
rect 25148 28472 25176 28512
rect 26237 28509 26249 28512
rect 26283 28540 26295 28543
rect 26697 28543 26755 28549
rect 26697 28540 26709 28543
rect 26283 28512 26709 28540
rect 26283 28509 26295 28512
rect 26237 28503 26295 28509
rect 26697 28509 26709 28512
rect 26743 28540 26755 28543
rect 28902 28540 28908 28552
rect 26743 28512 28908 28540
rect 26743 28509 26755 28512
rect 26697 28503 26755 28509
rect 28902 28500 28908 28512
rect 28960 28500 28966 28552
rect 29362 28500 29368 28552
rect 29420 28540 29426 28552
rect 29549 28543 29607 28549
rect 29549 28540 29561 28543
rect 29420 28512 29561 28540
rect 29420 28500 29426 28512
rect 29549 28509 29561 28512
rect 29595 28509 29607 28543
rect 29549 28503 29607 28509
rect 29733 28543 29791 28549
rect 29733 28509 29745 28543
rect 29779 28540 29791 28543
rect 30466 28540 30472 28552
rect 29779 28512 30472 28540
rect 29779 28509 29791 28512
rect 29733 28503 29791 28509
rect 23532 28444 25176 28472
rect 25225 28475 25283 28481
rect 23532 28432 23538 28444
rect 25225 28441 25237 28475
rect 25271 28472 25283 28475
rect 25406 28472 25412 28484
rect 25271 28444 25412 28472
rect 25271 28441 25283 28444
rect 25225 28435 25283 28441
rect 25406 28432 25412 28444
rect 25464 28472 25470 28484
rect 27154 28472 27160 28484
rect 25464 28444 27160 28472
rect 25464 28432 25470 28444
rect 27154 28432 27160 28444
rect 27212 28432 27218 28484
rect 29748 28472 29776 28503
rect 30466 28500 30472 28512
rect 30524 28500 30530 28552
rect 31021 28543 31079 28549
rect 31021 28509 31033 28543
rect 31067 28540 31079 28543
rect 33778 28540 33784 28552
rect 31067 28512 31524 28540
rect 33739 28512 33784 28540
rect 31067 28509 31079 28512
rect 31021 28503 31079 28509
rect 29012 28444 29776 28472
rect 13924 28404 13952 28432
rect 29012 28416 29040 28444
rect 31496 28416 31524 28512
rect 33778 28500 33784 28512
rect 33836 28540 33842 28552
rect 34992 28549 35020 28580
rect 35894 28568 35900 28580
rect 35952 28568 35958 28620
rect 36078 28568 36084 28620
rect 36136 28608 36142 28620
rect 36136 28580 36216 28608
rect 36136 28568 36142 28580
rect 34885 28543 34943 28549
rect 34885 28540 34897 28543
rect 33836 28512 34897 28540
rect 33836 28500 33842 28512
rect 34885 28509 34897 28512
rect 34931 28509 34943 28543
rect 34885 28503 34943 28509
rect 34977 28543 35035 28549
rect 34977 28509 34989 28543
rect 35023 28509 35035 28543
rect 34977 28503 35035 28509
rect 35253 28543 35311 28549
rect 35253 28509 35265 28543
rect 35299 28540 35311 28543
rect 35434 28540 35440 28552
rect 35299 28512 35440 28540
rect 35299 28509 35311 28512
rect 35253 28503 35311 28509
rect 35434 28500 35440 28512
rect 35492 28500 35498 28552
rect 35986 28540 35992 28552
rect 35947 28512 35992 28540
rect 35986 28500 35992 28512
rect 36044 28500 36050 28552
rect 36188 28546 36216 28580
rect 36283 28549 36311 28636
rect 36446 28549 36452 28552
rect 36173 28540 36231 28546
rect 36173 28506 36185 28540
rect 36219 28506 36231 28540
rect 36173 28500 36231 28506
rect 36268 28543 36326 28549
rect 36268 28509 36280 28543
rect 36314 28509 36326 28543
rect 36268 28503 36326 28509
rect 36403 28543 36452 28549
rect 36403 28509 36415 28543
rect 36449 28509 36452 28543
rect 36403 28503 36452 28509
rect 36446 28500 36452 28503
rect 36504 28500 36510 28552
rect 37108 28549 37136 28648
rect 37093 28543 37151 28549
rect 37093 28509 37105 28543
rect 37139 28509 37151 28543
rect 37093 28503 37151 28509
rect 34422 28432 34428 28484
rect 34480 28472 34486 28484
rect 35069 28475 35127 28481
rect 35069 28472 35081 28475
rect 34480 28444 35081 28472
rect 34480 28432 34486 28444
rect 35069 28441 35081 28444
rect 35115 28441 35127 28475
rect 37274 28472 37280 28484
rect 37235 28444 37280 28472
rect 35069 28435 35127 28441
rect 37274 28432 37280 28444
rect 37332 28432 37338 28484
rect 15286 28404 15292 28416
rect 13188 28376 13952 28404
rect 15247 28376 15292 28404
rect 15286 28364 15292 28376
rect 15344 28364 15350 28416
rect 16942 28404 16948 28416
rect 16903 28376 16948 28404
rect 16942 28364 16948 28376
rect 17000 28364 17006 28416
rect 17954 28364 17960 28416
rect 18012 28404 18018 28416
rect 18141 28407 18199 28413
rect 18141 28404 18153 28407
rect 18012 28376 18153 28404
rect 18012 28364 18018 28376
rect 18141 28373 18153 28376
rect 18187 28373 18199 28407
rect 28994 28404 29000 28416
rect 28955 28376 29000 28404
rect 18141 28367 18199 28373
rect 28994 28364 29000 28376
rect 29052 28364 29058 28416
rect 31478 28404 31484 28416
rect 31439 28376 31484 28404
rect 31478 28364 31484 28376
rect 31536 28364 31542 28416
rect 34698 28404 34704 28416
rect 34659 28376 34704 28404
rect 34698 28364 34704 28376
rect 34756 28364 34762 28416
rect 37458 28404 37464 28416
rect 37419 28376 37464 28404
rect 37458 28364 37464 28376
rect 37516 28364 37522 28416
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 3786 28200 3792 28212
rect 3747 28172 3792 28200
rect 3786 28160 3792 28172
rect 3844 28160 3850 28212
rect 8570 28200 8576 28212
rect 6196 28172 6914 28200
rect 8531 28172 8576 28200
rect 2498 28092 2504 28144
rect 2556 28132 2562 28144
rect 2654 28135 2712 28141
rect 2654 28132 2666 28135
rect 2556 28104 2666 28132
rect 2556 28092 2562 28104
rect 2654 28101 2666 28104
rect 2700 28101 2712 28135
rect 5350 28132 5356 28144
rect 5311 28104 5356 28132
rect 2654 28095 2712 28101
rect 5350 28092 5356 28104
rect 5408 28092 5414 28144
rect 4982 28064 4988 28076
rect 4943 28036 4988 28064
rect 4982 28024 4988 28036
rect 5040 28024 5046 28076
rect 5078 28067 5136 28073
rect 5078 28033 5090 28067
rect 5124 28033 5136 28067
rect 5078 28027 5136 28033
rect 5261 28067 5319 28073
rect 5261 28033 5273 28067
rect 5307 28033 5319 28067
rect 5442 28064 5448 28076
rect 5401 28036 5448 28064
rect 5261 28027 5319 28033
rect 2406 27996 2412 28008
rect 2367 27968 2412 27996
rect 2406 27956 2412 27968
rect 2464 27956 2470 28008
rect 3602 27956 3608 28008
rect 3660 27996 3666 28008
rect 5092 27996 5120 28027
rect 3660 27968 5120 27996
rect 3660 27956 3666 27968
rect 5166 27956 5172 28008
rect 5224 27996 5230 28008
rect 5276 27996 5304 28027
rect 5442 28024 5448 28036
rect 5500 28073 5506 28076
rect 5500 28067 5549 28073
rect 5500 28033 5503 28067
rect 5537 28064 5549 28067
rect 6196 28064 6224 28172
rect 6730 28132 6736 28144
rect 6691 28104 6736 28132
rect 6730 28092 6736 28104
rect 6788 28092 6794 28144
rect 6362 28064 6368 28076
rect 5537 28036 6224 28064
rect 6323 28036 6368 28064
rect 5537 28033 5549 28036
rect 5500 28027 5549 28033
rect 5500 28024 5506 28027
rect 6362 28024 6368 28036
rect 6420 28024 6426 28076
rect 6546 28073 6552 28076
rect 6513 28067 6552 28073
rect 6513 28033 6525 28067
rect 6513 28027 6552 28033
rect 6546 28024 6552 28027
rect 6604 28024 6610 28076
rect 6886 28073 6914 28172
rect 8570 28160 8576 28172
rect 8628 28160 8634 28212
rect 9398 28200 9404 28212
rect 9359 28172 9404 28200
rect 9398 28160 9404 28172
rect 9456 28160 9462 28212
rect 11517 28203 11575 28209
rect 11517 28169 11529 28203
rect 11563 28200 11575 28203
rect 12526 28200 12532 28212
rect 11563 28172 12532 28200
rect 11563 28169 11575 28172
rect 11517 28163 11575 28169
rect 12526 28160 12532 28172
rect 12584 28160 12590 28212
rect 13081 28203 13139 28209
rect 13081 28169 13093 28203
rect 13127 28200 13139 28203
rect 13354 28200 13360 28212
rect 13127 28172 13360 28200
rect 13127 28169 13139 28172
rect 13081 28163 13139 28169
rect 13354 28160 13360 28172
rect 13412 28160 13418 28212
rect 13906 28200 13912 28212
rect 13867 28172 13912 28200
rect 13906 28160 13912 28172
rect 13964 28160 13970 28212
rect 14366 28200 14372 28212
rect 14327 28172 14372 28200
rect 14366 28160 14372 28172
rect 14424 28160 14430 28212
rect 17954 28160 17960 28212
rect 18012 28200 18018 28212
rect 28994 28200 29000 28212
rect 18012 28172 29000 28200
rect 18012 28160 18018 28172
rect 28994 28160 29000 28172
rect 29052 28160 29058 28212
rect 30285 28203 30343 28209
rect 30285 28169 30297 28203
rect 30331 28200 30343 28203
rect 30834 28200 30840 28212
rect 30331 28172 30840 28200
rect 30331 28169 30343 28172
rect 30285 28163 30343 28169
rect 30834 28160 30840 28172
rect 30892 28160 30898 28212
rect 34422 28160 34428 28212
rect 34480 28160 34486 28212
rect 35526 28200 35532 28212
rect 35487 28172 35532 28200
rect 35526 28160 35532 28172
rect 35584 28200 35590 28212
rect 35584 28172 36492 28200
rect 35584 28160 35590 28172
rect 9674 28132 9680 28144
rect 8404 28104 9680 28132
rect 6641 28067 6699 28073
rect 6641 28033 6653 28067
rect 6687 28033 6699 28067
rect 6641 28027 6699 28033
rect 6869 28067 6927 28073
rect 6869 28033 6881 28067
rect 6915 28064 6927 28067
rect 7098 28064 7104 28076
rect 6915 28036 7104 28064
rect 6915 28033 6927 28036
rect 6869 28027 6927 28033
rect 6656 27996 6684 28027
rect 7098 28024 7104 28036
rect 7156 28064 7162 28076
rect 8404 28073 8432 28104
rect 9674 28092 9680 28104
rect 9732 28092 9738 28144
rect 10594 28092 10600 28144
rect 10652 28132 10658 28144
rect 12710 28132 12716 28144
rect 10652 28104 12434 28132
rect 12623 28104 12716 28132
rect 10652 28092 10658 28104
rect 8389 28067 8447 28073
rect 8389 28064 8401 28067
rect 7156 28036 8401 28064
rect 7156 28024 7162 28036
rect 8389 28033 8401 28036
rect 8435 28033 8447 28067
rect 8389 28027 8447 28033
rect 8573 28067 8631 28073
rect 8573 28033 8585 28067
rect 8619 28033 8631 28067
rect 8573 28027 8631 28033
rect 9217 28067 9275 28073
rect 9217 28033 9229 28067
rect 9263 28033 9275 28067
rect 9217 28027 9275 28033
rect 9401 28067 9459 28073
rect 9401 28033 9413 28067
rect 9447 28064 9459 28067
rect 9490 28064 9496 28076
rect 9447 28036 9496 28064
rect 9447 28033 9459 28036
rect 9401 28027 9459 28033
rect 7929 27999 7987 28005
rect 5224 27968 6868 27996
rect 5224 27956 5230 27968
rect 6840 27940 6868 27968
rect 7929 27965 7941 27999
rect 7975 27996 7987 27999
rect 8202 27996 8208 28008
rect 7975 27968 8208 27996
rect 7975 27965 7987 27968
rect 7929 27959 7987 27965
rect 8202 27956 8208 27968
rect 8260 27996 8266 28008
rect 8588 27996 8616 28027
rect 8260 27968 8616 27996
rect 9232 27996 9260 28027
rect 9490 28024 9496 28036
rect 9548 28024 9554 28076
rect 11606 28024 11612 28076
rect 11664 28064 11670 28076
rect 11701 28067 11759 28073
rect 11701 28064 11713 28067
rect 11664 28036 11713 28064
rect 11664 28024 11670 28036
rect 11701 28033 11713 28036
rect 11747 28033 11759 28067
rect 11701 28027 11759 28033
rect 11790 28024 11796 28076
rect 11848 28064 11854 28076
rect 12406 28064 12434 28104
rect 12710 28092 12716 28104
rect 12768 28132 12774 28144
rect 13262 28132 13268 28144
rect 12768 28104 13268 28132
rect 12768 28092 12774 28104
rect 13262 28092 13268 28104
rect 13320 28092 13326 28144
rect 15286 28092 15292 28144
rect 15344 28132 15350 28144
rect 15482 28135 15540 28141
rect 15482 28132 15494 28135
rect 15344 28104 15494 28132
rect 15344 28092 15350 28104
rect 15482 28101 15494 28104
rect 15528 28101 15540 28135
rect 15482 28095 15540 28101
rect 22281 28135 22339 28141
rect 22281 28101 22293 28135
rect 22327 28132 22339 28135
rect 22554 28132 22560 28144
rect 22327 28104 22560 28132
rect 22327 28101 22339 28104
rect 22281 28095 22339 28101
rect 22554 28092 22560 28104
rect 22612 28092 22618 28144
rect 30742 28092 30748 28144
rect 30800 28132 30806 28144
rect 31478 28132 31484 28144
rect 30800 28104 31484 28132
rect 30800 28092 30806 28104
rect 31478 28092 31484 28104
rect 31536 28132 31542 28144
rect 34440 28132 34468 28160
rect 34517 28135 34575 28141
rect 34517 28132 34529 28135
rect 31536 28104 31754 28132
rect 31536 28092 31542 28104
rect 12529 28067 12587 28073
rect 12529 28064 12541 28067
rect 11848 28036 11893 28064
rect 12406 28036 12541 28064
rect 11848 28024 11854 28036
rect 12529 28033 12541 28036
rect 12575 28033 12587 28067
rect 12529 28027 12587 28033
rect 12618 28024 12624 28076
rect 12676 28064 12682 28076
rect 12805 28067 12863 28073
rect 12805 28064 12817 28067
rect 12676 28036 12817 28064
rect 12676 28024 12682 28036
rect 12805 28033 12817 28036
rect 12851 28033 12863 28067
rect 12805 28027 12863 28033
rect 12897 28067 12955 28073
rect 12897 28033 12909 28067
rect 12943 28064 12955 28067
rect 13170 28064 13176 28076
rect 12943 28036 13176 28064
rect 12943 28033 12955 28036
rect 12897 28027 12955 28033
rect 13170 28024 13176 28036
rect 13228 28024 13234 28076
rect 15194 28064 15200 28076
rect 14752 28036 15200 28064
rect 9766 27996 9772 28008
rect 9232 27968 9772 27996
rect 8260 27956 8266 27968
rect 6822 27888 6828 27940
rect 6880 27888 6886 27940
rect 8588 27928 8616 27968
rect 9766 27956 9772 27968
rect 9824 27996 9830 28008
rect 10870 27996 10876 28008
rect 9824 27968 10876 27996
rect 9824 27956 9830 27968
rect 10870 27956 10876 27968
rect 10928 27956 10934 28008
rect 11808 27996 11836 28024
rect 14752 27996 14780 28036
rect 15194 28024 15200 28036
rect 15252 28024 15258 28076
rect 15746 28064 15752 28076
rect 15707 28036 15752 28064
rect 15746 28024 15752 28036
rect 15804 28024 15810 28076
rect 16942 28024 16948 28076
rect 17000 28064 17006 28076
rect 17129 28067 17187 28073
rect 17129 28064 17141 28067
rect 17000 28036 17141 28064
rect 17000 28024 17006 28036
rect 17129 28033 17141 28036
rect 17175 28033 17187 28067
rect 17129 28027 17187 28033
rect 18509 28067 18567 28073
rect 18509 28033 18521 28067
rect 18555 28064 18567 28067
rect 20070 28064 20076 28076
rect 18555 28036 20076 28064
rect 18555 28033 18567 28036
rect 18509 28027 18567 28033
rect 11808 27968 14780 27996
rect 14734 27928 14740 27940
rect 8588 27900 14740 27928
rect 14734 27888 14740 27900
rect 14792 27888 14798 27940
rect 17144 27928 17172 28027
rect 20070 28024 20076 28036
rect 20128 28024 20134 28076
rect 29362 28024 29368 28076
rect 29420 28064 29426 28076
rect 30098 28064 30104 28076
rect 29420 28036 30104 28064
rect 29420 28024 29426 28036
rect 30098 28024 30104 28036
rect 30156 28024 30162 28076
rect 31297 28067 31355 28073
rect 31297 28033 31309 28067
rect 31343 28033 31355 28067
rect 31297 28027 31355 28033
rect 31573 28067 31631 28073
rect 31573 28033 31585 28067
rect 31619 28064 31631 28067
rect 31726 28064 31754 28104
rect 33704 28104 34529 28132
rect 33704 28073 33732 28104
rect 34517 28101 34529 28104
rect 34563 28101 34575 28135
rect 34517 28095 34575 28101
rect 36170 28092 36176 28144
rect 36228 28132 36234 28144
rect 36464 28132 36492 28172
rect 36725 28135 36783 28141
rect 36228 28104 36400 28132
rect 36464 28104 36512 28132
rect 36228 28092 36234 28104
rect 32125 28067 32183 28073
rect 32125 28064 32137 28067
rect 31619 28036 32137 28064
rect 31619 28033 31631 28036
rect 31573 28027 31631 28033
rect 32125 28033 32137 28036
rect 32171 28033 32183 28067
rect 33689 28067 33747 28073
rect 33689 28064 33701 28067
rect 32125 28027 32183 28033
rect 33336 28036 33701 28064
rect 18230 27996 18236 28008
rect 18191 27968 18236 27996
rect 18230 27956 18236 27968
rect 18288 27956 18294 28008
rect 19334 27956 19340 28008
rect 19392 27996 19398 28008
rect 19521 27999 19579 28005
rect 19521 27996 19533 27999
rect 19392 27968 19533 27996
rect 19392 27956 19398 27968
rect 19521 27965 19533 27968
rect 19567 27965 19579 27999
rect 19521 27959 19579 27965
rect 19797 27999 19855 28005
rect 19797 27965 19809 27999
rect 19843 27996 19855 27999
rect 20254 27996 20260 28008
rect 19843 27968 20260 27996
rect 19843 27965 19855 27968
rect 19797 27959 19855 27965
rect 20254 27956 20260 27968
rect 20312 27956 20318 28008
rect 29917 27999 29975 28005
rect 29917 27996 29929 27999
rect 29380 27968 29929 27996
rect 17144 27900 24348 27928
rect 5629 27863 5687 27869
rect 5629 27829 5641 27863
rect 5675 27860 5687 27863
rect 5810 27860 5816 27872
rect 5675 27832 5816 27860
rect 5675 27829 5687 27832
rect 5629 27823 5687 27829
rect 5810 27820 5816 27832
rect 5868 27820 5874 27872
rect 7009 27863 7067 27869
rect 7009 27829 7021 27863
rect 7055 27860 7067 27863
rect 7834 27860 7840 27872
rect 7055 27832 7840 27860
rect 7055 27829 7067 27832
rect 7009 27823 7067 27829
rect 7834 27820 7840 27832
rect 7892 27820 7898 27872
rect 9490 27820 9496 27872
rect 9548 27860 9554 27872
rect 9861 27863 9919 27869
rect 9861 27860 9873 27863
rect 9548 27832 9873 27860
rect 9548 27820 9554 27832
rect 9861 27829 9873 27832
rect 9907 27829 9919 27863
rect 9861 27823 9919 27829
rect 17221 27863 17279 27869
rect 17221 27829 17233 27863
rect 17267 27860 17279 27863
rect 17310 27860 17316 27872
rect 17267 27832 17316 27860
rect 17267 27829 17279 27832
rect 17221 27823 17279 27829
rect 17310 27820 17316 27832
rect 17368 27860 17374 27872
rect 17678 27860 17684 27872
rect 17368 27832 17684 27860
rect 17368 27820 17374 27832
rect 17678 27820 17684 27832
rect 17736 27820 17742 27872
rect 22278 27820 22284 27872
rect 22336 27860 22342 27872
rect 24320 27869 24348 27900
rect 22373 27863 22431 27869
rect 22373 27860 22385 27863
rect 22336 27832 22385 27860
rect 22336 27820 22342 27832
rect 22373 27829 22385 27832
rect 22419 27829 22431 27863
rect 22373 27823 22431 27829
rect 24305 27863 24363 27869
rect 24305 27829 24317 27863
rect 24351 27860 24363 27863
rect 24854 27860 24860 27872
rect 24351 27832 24860 27860
rect 24351 27829 24363 27832
rect 24305 27823 24363 27829
rect 24854 27820 24860 27832
rect 24912 27860 24918 27872
rect 25498 27860 25504 27872
rect 24912 27832 25504 27860
rect 24912 27820 24918 27832
rect 25498 27820 25504 27832
rect 25556 27820 25562 27872
rect 29270 27820 29276 27872
rect 29328 27860 29334 27872
rect 29380 27869 29408 27968
rect 29917 27965 29929 27968
rect 29963 27965 29975 27999
rect 31312 27996 31340 28027
rect 33134 27996 33140 28008
rect 31312 27968 33140 27996
rect 29917 27959 29975 27965
rect 29932 27928 29960 27959
rect 33134 27956 33140 27968
rect 33192 27996 33198 28008
rect 33336 27996 33364 28036
rect 33689 28033 33701 28036
rect 33735 28033 33747 28067
rect 33689 28027 33747 28033
rect 33778 28024 33784 28076
rect 33836 28064 33842 28076
rect 34333 28067 34391 28073
rect 34333 28064 34345 28067
rect 33836 28036 34345 28064
rect 33836 28024 33842 28036
rect 34333 28033 34345 28036
rect 34379 28033 34391 28067
rect 34333 28027 34391 28033
rect 34425 28067 34483 28073
rect 34425 28033 34437 28067
rect 34471 28033 34483 28067
rect 34425 28027 34483 28033
rect 34701 28067 34759 28073
rect 34701 28033 34713 28067
rect 34747 28064 34759 28067
rect 34790 28064 34796 28076
rect 34747 28036 34796 28064
rect 34747 28033 34759 28036
rect 34701 28027 34759 28033
rect 33192 27968 33364 27996
rect 33413 27999 33471 28005
rect 33192 27956 33198 27968
rect 33413 27965 33425 27999
rect 33459 27996 33471 27999
rect 33870 27996 33876 28008
rect 33459 27968 33876 27996
rect 33459 27965 33471 27968
rect 33413 27959 33471 27965
rect 33870 27956 33876 27968
rect 33928 27956 33934 28008
rect 32398 27928 32404 27940
rect 29932 27900 32404 27928
rect 32398 27888 32404 27900
rect 32456 27888 32462 27940
rect 34440 27928 34468 28027
rect 34790 28024 34796 28036
rect 34848 28024 34854 28076
rect 35986 28024 35992 28076
rect 36044 28064 36050 28076
rect 36372 28073 36400 28104
rect 36484 28073 36512 28104
rect 36725 28101 36737 28135
rect 36771 28132 36783 28135
rect 38482 28135 38540 28141
rect 38482 28132 38494 28135
rect 36771 28104 38494 28132
rect 36771 28101 36783 28104
rect 36725 28095 36783 28101
rect 38482 28101 38494 28104
rect 38528 28101 38540 28135
rect 38482 28095 38540 28101
rect 36081 28067 36139 28073
rect 36081 28064 36093 28067
rect 36044 28036 36093 28064
rect 36044 28024 36050 28036
rect 36081 28033 36093 28036
rect 36127 28033 36139 28067
rect 36081 28027 36139 28033
rect 36265 28067 36323 28073
rect 36265 28033 36277 28067
rect 36311 28033 36323 28067
rect 36265 28027 36323 28033
rect 36357 28067 36415 28073
rect 36357 28033 36369 28067
rect 36403 28033 36415 28067
rect 36484 28067 36553 28073
rect 36484 28036 36507 28067
rect 36357 28027 36415 28033
rect 36495 28033 36507 28036
rect 36541 28033 36553 28067
rect 38746 28064 38752 28076
rect 38707 28036 38752 28064
rect 36495 28027 36553 28033
rect 36280 27996 36308 28027
rect 38746 28024 38752 28036
rect 38804 28024 38810 28076
rect 37458 27996 37464 28008
rect 36280 27968 37464 27996
rect 37458 27956 37464 27968
rect 37516 27956 37522 28008
rect 37274 27928 37280 27940
rect 34440 27900 37280 27928
rect 37274 27888 37280 27900
rect 37332 27928 37338 27940
rect 37369 27931 37427 27937
rect 37369 27928 37381 27931
rect 37332 27900 37381 27928
rect 37332 27888 37338 27900
rect 37369 27897 37381 27900
rect 37415 27897 37427 27931
rect 58158 27928 58164 27940
rect 58119 27900 58164 27928
rect 37369 27891 37427 27897
rect 58158 27888 58164 27900
rect 58216 27888 58222 27940
rect 29365 27863 29423 27869
rect 29365 27860 29377 27863
rect 29328 27832 29377 27860
rect 29328 27820 29334 27832
rect 29365 27829 29377 27832
rect 29411 27829 29423 27863
rect 29365 27823 29423 27829
rect 32950 27820 32956 27872
rect 33008 27860 33014 27872
rect 34149 27863 34207 27869
rect 34149 27860 34161 27863
rect 33008 27832 34161 27860
rect 33008 27820 33014 27832
rect 34149 27829 34161 27832
rect 34195 27829 34207 27863
rect 34149 27823 34207 27829
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 11701 27659 11759 27665
rect 11701 27625 11713 27659
rect 11747 27656 11759 27659
rect 11790 27656 11796 27668
rect 11747 27628 11796 27656
rect 11747 27625 11759 27628
rect 11701 27619 11759 27625
rect 11790 27616 11796 27628
rect 11848 27616 11854 27668
rect 12434 27616 12440 27668
rect 12492 27656 12498 27668
rect 13541 27659 13599 27665
rect 13541 27656 13553 27659
rect 12492 27628 13553 27656
rect 12492 27616 12498 27628
rect 13541 27625 13553 27628
rect 13587 27625 13599 27659
rect 13541 27619 13599 27625
rect 5074 27548 5080 27600
rect 5132 27588 5138 27600
rect 5537 27591 5595 27597
rect 5132 27560 5304 27588
rect 5132 27548 5138 27560
rect 4890 27452 4896 27464
rect 4851 27424 4896 27452
rect 4890 27412 4896 27424
rect 4948 27412 4954 27464
rect 4986 27455 5044 27461
rect 4986 27421 4998 27455
rect 5032 27421 5044 27455
rect 5166 27452 5172 27464
rect 5127 27424 5172 27452
rect 4986 27415 5044 27421
rect 3050 27344 3056 27396
rect 3108 27384 3114 27396
rect 5000 27384 5028 27415
rect 5166 27412 5172 27424
rect 5224 27412 5230 27464
rect 5276 27461 5304 27560
rect 5537 27557 5549 27591
rect 5583 27588 5595 27591
rect 8478 27588 8484 27600
rect 5583 27560 8484 27588
rect 5583 27557 5595 27560
rect 5537 27551 5595 27557
rect 8478 27548 8484 27560
rect 8536 27548 8542 27600
rect 17129 27591 17187 27597
rect 17129 27588 17141 27591
rect 16408 27560 17141 27588
rect 6546 27480 6552 27532
rect 6604 27520 6610 27532
rect 6604 27492 7972 27520
rect 6604 27480 6610 27492
rect 5442 27461 5448 27464
rect 5261 27455 5319 27461
rect 5261 27421 5273 27455
rect 5307 27421 5319 27455
rect 5261 27415 5319 27421
rect 5399 27455 5448 27461
rect 5399 27421 5411 27455
rect 5445 27421 5448 27455
rect 5399 27415 5448 27421
rect 5442 27412 5448 27415
rect 5500 27412 5506 27464
rect 6454 27412 6460 27464
rect 6512 27452 6518 27464
rect 6641 27455 6699 27461
rect 6641 27452 6653 27455
rect 6512 27424 6653 27452
rect 6512 27412 6518 27424
rect 6641 27421 6653 27424
rect 6687 27421 6699 27455
rect 6641 27415 6699 27421
rect 6734 27455 6792 27461
rect 6734 27421 6746 27455
rect 6780 27421 6792 27455
rect 7006 27452 7012 27464
rect 6967 27424 7012 27452
rect 6734 27415 6792 27421
rect 3108 27356 5028 27384
rect 3108 27344 3114 27356
rect 5626 27344 5632 27396
rect 5684 27384 5690 27396
rect 6748 27384 6776 27415
rect 7006 27412 7012 27424
rect 7064 27412 7070 27464
rect 7098 27412 7104 27464
rect 7156 27461 7162 27464
rect 7944 27461 7972 27492
rect 8202 27480 8208 27532
rect 8260 27520 8266 27532
rect 9306 27520 9312 27532
rect 8260 27492 9312 27520
rect 8260 27480 8266 27492
rect 9306 27480 9312 27492
rect 9364 27520 9370 27532
rect 9364 27492 12204 27520
rect 9364 27480 9370 27492
rect 12176 27464 12204 27492
rect 7156 27452 7164 27461
rect 7929 27455 7987 27461
rect 7156 27424 7201 27452
rect 7300 27424 7880 27452
rect 7156 27415 7164 27424
rect 7156 27412 7162 27415
rect 5684 27356 6776 27384
rect 5684 27344 5690 27356
rect 6822 27344 6828 27396
rect 6880 27384 6886 27396
rect 6917 27387 6975 27393
rect 6917 27384 6929 27387
rect 6880 27356 6929 27384
rect 6880 27344 6886 27356
rect 6917 27353 6929 27356
rect 6963 27384 6975 27387
rect 7300 27384 7328 27424
rect 7742 27384 7748 27396
rect 6963 27356 7328 27384
rect 7703 27356 7748 27384
rect 6963 27353 6975 27356
rect 6917 27347 6975 27353
rect 7742 27344 7748 27356
rect 7800 27344 7806 27396
rect 7852 27384 7880 27424
rect 7929 27421 7941 27455
rect 7975 27421 7987 27455
rect 9214 27452 9220 27464
rect 9175 27424 9220 27452
rect 7929 27415 7987 27421
rect 9214 27412 9220 27424
rect 9272 27412 9278 27464
rect 9401 27455 9459 27461
rect 9401 27421 9413 27455
rect 9447 27452 9459 27455
rect 9490 27452 9496 27464
rect 9447 27424 9496 27452
rect 9447 27421 9459 27424
rect 9401 27415 9459 27421
rect 9490 27412 9496 27424
rect 9548 27412 9554 27464
rect 10870 27452 10876 27464
rect 10831 27424 10876 27452
rect 10870 27412 10876 27424
rect 10928 27412 10934 27464
rect 11146 27452 11152 27464
rect 11107 27424 11152 27452
rect 11146 27412 11152 27424
rect 11204 27412 11210 27464
rect 12158 27452 12164 27464
rect 12119 27424 12164 27452
rect 12158 27412 12164 27424
rect 12216 27412 12222 27464
rect 12428 27455 12486 27461
rect 12428 27421 12440 27455
rect 12474 27452 12486 27455
rect 12894 27452 12900 27464
rect 12474 27424 12900 27452
rect 12474 27421 12486 27424
rect 12428 27415 12486 27421
rect 12894 27412 12900 27424
rect 12952 27412 12958 27464
rect 14734 27412 14740 27464
rect 14792 27452 14798 27464
rect 16408 27452 16436 27560
rect 17129 27557 17141 27560
rect 17175 27588 17187 27591
rect 17954 27588 17960 27600
rect 17175 27560 17960 27588
rect 17175 27557 17187 27560
rect 17129 27551 17187 27557
rect 17954 27548 17960 27560
rect 18012 27548 18018 27600
rect 21085 27591 21143 27597
rect 21085 27557 21097 27591
rect 21131 27588 21143 27591
rect 22370 27588 22376 27600
rect 21131 27560 22376 27588
rect 21131 27557 21143 27560
rect 21085 27551 21143 27557
rect 22370 27548 22376 27560
rect 22428 27548 22434 27600
rect 25314 27520 25320 27532
rect 18156 27492 25320 27520
rect 16477 27455 16535 27461
rect 16477 27452 16489 27455
rect 14792 27424 16489 27452
rect 14792 27412 14798 27424
rect 16477 27421 16489 27424
rect 16523 27421 16535 27455
rect 16666 27452 16672 27464
rect 16627 27424 16672 27452
rect 16477 27415 16535 27421
rect 16666 27412 16672 27424
rect 16724 27412 16730 27464
rect 9232 27384 9260 27412
rect 16574 27384 16580 27396
rect 7852 27356 9260 27384
rect 16487 27356 16580 27384
rect 16574 27344 16580 27356
rect 16632 27384 16638 27396
rect 18156 27384 18184 27492
rect 25314 27480 25320 27492
rect 25372 27480 25378 27532
rect 30098 27480 30104 27532
rect 30156 27520 30162 27532
rect 30653 27523 30711 27529
rect 30653 27520 30665 27523
rect 30156 27492 30665 27520
rect 30156 27480 30162 27492
rect 30653 27489 30665 27492
rect 30699 27489 30711 27523
rect 30653 27483 30711 27489
rect 20441 27455 20499 27461
rect 20441 27421 20453 27455
rect 20487 27452 20499 27455
rect 20714 27452 20720 27464
rect 20487 27424 20720 27452
rect 20487 27421 20499 27424
rect 20441 27415 20499 27421
rect 20714 27412 20720 27424
rect 20772 27452 20778 27464
rect 20901 27455 20959 27461
rect 20901 27452 20913 27455
rect 20772 27424 20913 27452
rect 20772 27412 20778 27424
rect 20901 27421 20913 27424
rect 20947 27452 20959 27455
rect 21266 27452 21272 27464
rect 20947 27424 21272 27452
rect 20947 27421 20959 27424
rect 20901 27415 20959 27421
rect 21266 27412 21272 27424
rect 21324 27412 21330 27464
rect 26421 27455 26479 27461
rect 26421 27421 26433 27455
rect 26467 27452 26479 27455
rect 27246 27452 27252 27464
rect 26467 27424 27252 27452
rect 26467 27421 26479 27424
rect 26421 27415 26479 27421
rect 27246 27412 27252 27424
rect 27304 27412 27310 27464
rect 30377 27455 30435 27461
rect 30377 27452 30389 27455
rect 29932 27424 30389 27452
rect 16632 27356 18184 27384
rect 16632 27344 16638 27356
rect 20990 27344 20996 27396
rect 21048 27384 21054 27396
rect 21637 27387 21695 27393
rect 21637 27384 21649 27387
rect 21048 27356 21649 27384
rect 21048 27344 21054 27356
rect 21637 27353 21649 27356
rect 21683 27353 21695 27387
rect 21637 27347 21695 27353
rect 21821 27387 21879 27393
rect 21821 27353 21833 27387
rect 21867 27384 21879 27387
rect 22554 27384 22560 27396
rect 21867 27356 22560 27384
rect 21867 27353 21879 27356
rect 21821 27347 21879 27353
rect 22554 27344 22560 27356
rect 22612 27344 22618 27396
rect 25406 27344 25412 27396
rect 25464 27384 25470 27396
rect 26666 27387 26724 27393
rect 26666 27384 26678 27387
rect 25464 27356 26678 27384
rect 25464 27344 25470 27356
rect 26666 27353 26678 27356
rect 26712 27353 26724 27387
rect 26666 27347 26724 27353
rect 29932 27328 29960 27424
rect 30377 27421 30389 27424
rect 30423 27421 30435 27455
rect 30377 27415 30435 27421
rect 33137 27455 33195 27461
rect 33137 27421 33149 27455
rect 33183 27452 33195 27455
rect 33318 27452 33324 27464
rect 33183 27424 33324 27452
rect 33183 27421 33195 27424
rect 33137 27415 33195 27421
rect 33318 27412 33324 27424
rect 33376 27412 33382 27464
rect 30834 27344 30840 27396
rect 30892 27384 30898 27396
rect 32953 27387 33011 27393
rect 32953 27384 32965 27387
rect 30892 27356 32965 27384
rect 30892 27344 30898 27356
rect 32953 27353 32965 27356
rect 32999 27384 33011 27387
rect 34606 27384 34612 27396
rect 32999 27356 34612 27384
rect 32999 27353 33011 27356
rect 32953 27347 33011 27353
rect 34606 27344 34612 27356
rect 34664 27344 34670 27396
rect 7285 27319 7343 27325
rect 7285 27285 7297 27319
rect 7331 27316 7343 27319
rect 7926 27316 7932 27328
rect 7331 27288 7932 27316
rect 7331 27285 7343 27288
rect 7285 27279 7343 27285
rect 7926 27276 7932 27288
rect 7984 27276 7990 27328
rect 8110 27316 8116 27328
rect 8071 27288 8116 27316
rect 8110 27276 8116 27288
rect 8168 27276 8174 27328
rect 8386 27276 8392 27328
rect 8444 27316 8450 27328
rect 9309 27319 9367 27325
rect 9309 27316 9321 27319
rect 8444 27288 9321 27316
rect 8444 27276 8450 27288
rect 9309 27285 9321 27288
rect 9355 27285 9367 27319
rect 17678 27316 17684 27328
rect 17639 27288 17684 27316
rect 9309 27279 9367 27285
rect 17678 27276 17684 27288
rect 17736 27276 17742 27328
rect 21910 27276 21916 27328
rect 21968 27316 21974 27328
rect 22005 27319 22063 27325
rect 22005 27316 22017 27319
rect 21968 27288 22017 27316
rect 21968 27276 21974 27288
rect 22005 27285 22017 27288
rect 22051 27285 22063 27319
rect 22005 27279 22063 27285
rect 22738 27276 22744 27328
rect 22796 27316 22802 27328
rect 24397 27319 24455 27325
rect 24397 27316 24409 27319
rect 22796 27288 24409 27316
rect 22796 27276 22802 27288
rect 24397 27285 24409 27288
rect 24443 27316 24455 27319
rect 24762 27316 24768 27328
rect 24443 27288 24768 27316
rect 24443 27285 24455 27288
rect 24397 27279 24455 27285
rect 24762 27276 24768 27288
rect 24820 27276 24826 27328
rect 27801 27319 27859 27325
rect 27801 27285 27813 27319
rect 27847 27316 27859 27319
rect 28994 27316 29000 27328
rect 27847 27288 29000 27316
rect 27847 27285 27859 27288
rect 27801 27279 27859 27285
rect 28994 27276 29000 27288
rect 29052 27276 29058 27328
rect 29914 27316 29920 27328
rect 29875 27288 29920 27316
rect 29914 27276 29920 27288
rect 29972 27276 29978 27328
rect 33321 27319 33379 27325
rect 33321 27285 33333 27319
rect 33367 27316 33379 27319
rect 33686 27316 33692 27328
rect 33367 27288 33692 27316
rect 33367 27285 33379 27288
rect 33321 27279 33379 27285
rect 33686 27276 33692 27288
rect 33744 27276 33750 27328
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 6546 27072 6552 27124
rect 6604 27112 6610 27124
rect 6825 27115 6883 27121
rect 6825 27112 6837 27115
rect 6604 27084 6837 27112
rect 6604 27072 6610 27084
rect 6825 27081 6837 27084
rect 6871 27081 6883 27115
rect 6825 27075 6883 27081
rect 10502 27072 10508 27124
rect 10560 27112 10566 27124
rect 20806 27112 20812 27124
rect 10560 27084 20812 27112
rect 10560 27072 10566 27084
rect 20806 27072 20812 27084
rect 20864 27072 20870 27124
rect 25038 27112 25044 27124
rect 24943 27084 25044 27112
rect 3602 27044 3608 27056
rect 3563 27016 3608 27044
rect 3602 27004 3608 27016
rect 3660 27004 3666 27056
rect 18690 27044 18696 27056
rect 16960 27016 18696 27044
rect 3234 26936 3240 26988
rect 3292 26976 3298 26988
rect 3421 26979 3479 26985
rect 3421 26976 3433 26979
rect 3292 26948 3433 26976
rect 3292 26936 3298 26948
rect 3421 26945 3433 26948
rect 3467 26976 3479 26979
rect 5442 26976 5448 26988
rect 3467 26948 5448 26976
rect 3467 26945 3479 26948
rect 3421 26939 3479 26945
rect 5442 26936 5448 26948
rect 5500 26936 5506 26988
rect 7926 26976 7932 26988
rect 7984 26985 7990 26988
rect 7896 26948 7932 26976
rect 7926 26936 7932 26948
rect 7984 26939 7996 26985
rect 8202 26976 8208 26988
rect 8163 26948 8208 26976
rect 7984 26936 7990 26939
rect 8202 26936 8208 26948
rect 8260 26936 8266 26988
rect 9214 26936 9220 26988
rect 9272 26976 9278 26988
rect 10045 26979 10103 26985
rect 10045 26976 10057 26979
rect 9272 26948 10057 26976
rect 9272 26936 9278 26948
rect 10045 26945 10057 26948
rect 10091 26945 10103 26979
rect 10045 26939 10103 26945
rect 11885 26979 11943 26985
rect 11885 26945 11897 26979
rect 11931 26976 11943 26979
rect 12710 26976 12716 26988
rect 11931 26948 12716 26976
rect 11931 26945 11943 26948
rect 11885 26939 11943 26945
rect 12710 26936 12716 26948
rect 12768 26936 12774 26988
rect 13170 26976 13176 26988
rect 13131 26948 13176 26976
rect 13170 26936 13176 26948
rect 13228 26936 13234 26988
rect 16960 26985 16988 27016
rect 18690 27004 18696 27016
rect 18748 27044 18754 27056
rect 18748 27016 19196 27044
rect 18748 27004 18754 27016
rect 16945 26979 17003 26985
rect 16945 26945 16957 26979
rect 16991 26945 17003 26979
rect 16945 26939 17003 26945
rect 17212 26979 17270 26985
rect 17212 26945 17224 26979
rect 17258 26976 17270 26979
rect 17494 26976 17500 26988
rect 17258 26948 17500 26976
rect 17258 26945 17270 26948
rect 17212 26939 17270 26945
rect 17494 26936 17500 26948
rect 17552 26936 17558 26988
rect 19168 26985 19196 27016
rect 22094 27004 22100 27056
rect 22152 27044 22158 27056
rect 22922 27044 22928 27056
rect 22152 27016 22928 27044
rect 22152 27004 22158 27016
rect 22922 27004 22928 27016
rect 22980 27044 22986 27056
rect 22980 27016 23796 27044
rect 22980 27004 22986 27016
rect 19153 26979 19211 26985
rect 19153 26945 19165 26979
rect 19199 26945 19211 26979
rect 19153 26939 19211 26945
rect 19242 26936 19248 26988
rect 19300 26976 19306 26988
rect 19409 26979 19467 26985
rect 19409 26976 19421 26979
rect 19300 26948 19421 26976
rect 19300 26936 19306 26948
rect 19409 26945 19421 26948
rect 19455 26945 19467 26979
rect 23474 26976 23480 26988
rect 23532 26985 23538 26988
rect 23768 26985 23796 27016
rect 24943 26991 24971 27084
rect 25038 27072 25044 27084
rect 25096 27072 25102 27124
rect 25406 27112 25412 27124
rect 25367 27084 25412 27112
rect 25406 27072 25412 27084
rect 25464 27072 25470 27124
rect 29362 27112 29368 27124
rect 26068 27084 29368 27112
rect 26068 27053 26096 27084
rect 29362 27072 29368 27084
rect 29420 27072 29426 27124
rect 33778 27112 33784 27124
rect 32784 27084 33784 27112
rect 26053 27047 26111 27053
rect 26053 27013 26065 27047
rect 26099 27013 26111 27047
rect 30926 27044 30932 27056
rect 26053 27007 26111 27013
rect 27908 27016 30932 27044
rect 23444 26948 23480 26976
rect 19409 26939 19467 26945
rect 23474 26936 23480 26948
rect 23532 26939 23544 26985
rect 23753 26979 23811 26985
rect 23753 26945 23765 26979
rect 23799 26945 23811 26979
rect 24762 26976 24768 26988
rect 24723 26948 24768 26976
rect 23753 26939 23811 26945
rect 23532 26936 23538 26939
rect 9769 26911 9827 26917
rect 9769 26877 9781 26911
rect 9815 26908 9827 26911
rect 9950 26908 9956 26920
rect 9815 26880 9956 26908
rect 9815 26877 9827 26880
rect 9769 26871 9827 26877
rect 9950 26868 9956 26880
rect 10008 26868 10014 26920
rect 11146 26868 11152 26920
rect 11204 26908 11210 26920
rect 11609 26911 11667 26917
rect 11609 26908 11621 26911
rect 11204 26880 11621 26908
rect 11204 26868 11210 26880
rect 11609 26877 11621 26880
rect 11655 26877 11667 26911
rect 11609 26871 11667 26877
rect 12434 26868 12440 26920
rect 12492 26908 12498 26920
rect 12897 26911 12955 26917
rect 12897 26908 12909 26911
rect 12492 26880 12909 26908
rect 12492 26868 12498 26880
rect 12897 26877 12909 26880
rect 12943 26877 12955 26911
rect 12897 26871 12955 26877
rect 8294 26800 8300 26852
rect 8352 26840 8358 26852
rect 8757 26843 8815 26849
rect 8757 26840 8769 26843
rect 8352 26812 8769 26840
rect 8352 26800 8358 26812
rect 8757 26809 8769 26812
rect 8803 26840 8815 26843
rect 9306 26840 9312 26852
rect 8803 26812 9312 26840
rect 8803 26809 8815 26812
rect 8757 26803 8815 26809
rect 9306 26800 9312 26812
rect 9364 26800 9370 26852
rect 23768 26840 23796 26939
rect 24762 26936 24768 26948
rect 24820 26936 24826 26988
rect 24928 26985 24986 26991
rect 24928 26951 24940 26985
rect 24974 26951 24986 26985
rect 24928 26945 24986 26951
rect 25044 26979 25102 26985
rect 25044 26945 25056 26979
rect 25090 26945 25102 26979
rect 25044 26939 25102 26945
rect 25179 26979 25237 26985
rect 25179 26945 25191 26979
rect 25225 26976 25237 26979
rect 25314 26976 25320 26988
rect 25225 26948 25320 26976
rect 25225 26945 25237 26948
rect 25179 26939 25237 26945
rect 24578 26868 24584 26920
rect 24636 26908 24642 26920
rect 25056 26908 25084 26939
rect 25314 26936 25320 26948
rect 25372 26936 25378 26988
rect 26237 26979 26295 26985
rect 26237 26945 26249 26979
rect 26283 26976 26295 26979
rect 27430 26976 27436 26988
rect 26283 26948 27436 26976
rect 26283 26945 26295 26948
rect 26237 26939 26295 26945
rect 27430 26936 27436 26948
rect 27488 26936 27494 26988
rect 27908 26985 27936 27016
rect 30926 27004 30932 27016
rect 30984 27004 30990 27056
rect 27893 26979 27951 26985
rect 27893 26945 27905 26979
rect 27939 26945 27951 26979
rect 27893 26939 27951 26945
rect 27982 26936 27988 26988
rect 28040 26976 28046 26988
rect 32784 26985 32812 27084
rect 33778 27072 33784 27084
rect 33836 27072 33842 27124
rect 32861 27047 32919 27053
rect 32861 27013 32873 27047
rect 32907 27044 32919 27047
rect 33318 27044 33324 27056
rect 32907 27016 33324 27044
rect 32907 27013 32919 27016
rect 32861 27007 32919 27013
rect 33318 27004 33324 27016
rect 33376 27004 33382 27056
rect 28149 26979 28207 26985
rect 28149 26976 28161 26979
rect 28040 26948 28161 26976
rect 28040 26936 28046 26948
rect 28149 26945 28161 26948
rect 28195 26945 28207 26979
rect 28149 26939 28207 26945
rect 31021 26979 31079 26985
rect 31021 26945 31033 26979
rect 31067 26976 31079 26979
rect 32769 26979 32827 26985
rect 32769 26976 32781 26979
rect 31067 26948 32781 26976
rect 31067 26945 31079 26948
rect 31021 26939 31079 26945
rect 32769 26945 32781 26948
rect 32815 26945 32827 26979
rect 32769 26939 32827 26945
rect 32953 26979 33011 26985
rect 32953 26945 32965 26979
rect 32999 26976 33011 26979
rect 33042 26976 33048 26988
rect 32999 26948 33048 26976
rect 32999 26945 33011 26948
rect 32953 26939 33011 26945
rect 33042 26936 33048 26948
rect 33100 26936 33106 26988
rect 33137 26979 33195 26985
rect 33137 26945 33149 26979
rect 33183 26976 33195 26979
rect 33226 26976 33232 26988
rect 33183 26948 33232 26976
rect 33183 26945 33195 26948
rect 33137 26939 33195 26945
rect 33226 26936 33232 26948
rect 33284 26936 33290 26988
rect 33796 26985 33824 27072
rect 33873 27047 33931 27053
rect 33873 27013 33885 27047
rect 33919 27044 33931 27047
rect 34514 27044 34520 27056
rect 33919 27016 34520 27044
rect 33919 27013 33931 27016
rect 33873 27007 33931 27013
rect 34514 27004 34520 27016
rect 34572 27044 34578 27056
rect 34793 27047 34851 27053
rect 34793 27044 34805 27047
rect 34572 27016 34805 27044
rect 34572 27004 34578 27016
rect 34793 27013 34805 27016
rect 34839 27013 34851 27047
rect 34793 27007 34851 27013
rect 33781 26979 33839 26985
rect 33781 26945 33793 26979
rect 33827 26945 33839 26979
rect 33781 26939 33839 26945
rect 33965 26979 34023 26985
rect 33965 26945 33977 26979
rect 34011 26945 34023 26979
rect 34146 26976 34152 26988
rect 34107 26948 34152 26976
rect 33965 26939 34023 26945
rect 30745 26911 30803 26917
rect 30745 26908 30757 26911
rect 24636 26880 25084 26908
rect 30208 26880 30757 26908
rect 24636 26868 24642 26880
rect 25590 26840 25596 26852
rect 23768 26812 25596 26840
rect 25590 26800 25596 26812
rect 25648 26800 25654 26852
rect 29914 26840 29920 26852
rect 29196 26812 29920 26840
rect 3789 26775 3847 26781
rect 3789 26741 3801 26775
rect 3835 26772 3847 26775
rect 3970 26772 3976 26784
rect 3835 26744 3976 26772
rect 3835 26741 3847 26744
rect 3789 26735 3847 26741
rect 3970 26732 3976 26744
rect 4028 26732 4034 26784
rect 9214 26772 9220 26784
rect 9175 26744 9220 26772
rect 9214 26732 9220 26744
rect 9272 26772 9278 26784
rect 9490 26772 9496 26784
rect 9272 26744 9496 26772
rect 9272 26732 9278 26744
rect 9490 26732 9496 26744
rect 9548 26732 9554 26784
rect 18325 26775 18383 26781
rect 18325 26741 18337 26775
rect 18371 26772 18383 26775
rect 20070 26772 20076 26784
rect 18371 26744 20076 26772
rect 18371 26741 18383 26744
rect 18325 26735 18383 26741
rect 20070 26732 20076 26744
rect 20128 26732 20134 26784
rect 20533 26775 20591 26781
rect 20533 26741 20545 26775
rect 20579 26772 20591 26775
rect 20622 26772 20628 26784
rect 20579 26744 20628 26772
rect 20579 26741 20591 26744
rect 20533 26735 20591 26741
rect 20622 26732 20628 26744
rect 20680 26732 20686 26784
rect 22373 26775 22431 26781
rect 22373 26741 22385 26775
rect 22419 26772 22431 26775
rect 22554 26772 22560 26784
rect 22419 26744 22560 26772
rect 22419 26741 22431 26744
rect 22373 26735 22431 26741
rect 22554 26732 22560 26744
rect 22612 26732 22618 26784
rect 24118 26732 24124 26784
rect 24176 26772 24182 26784
rect 24213 26775 24271 26781
rect 24213 26772 24225 26775
rect 24176 26744 24225 26772
rect 24176 26732 24182 26744
rect 24213 26741 24225 26744
rect 24259 26772 24271 26775
rect 25314 26772 25320 26784
rect 24259 26744 25320 26772
rect 24259 26741 24271 26744
rect 24213 26735 24271 26741
rect 25314 26732 25320 26744
rect 25372 26732 25378 26784
rect 25682 26732 25688 26784
rect 25740 26772 25746 26784
rect 25869 26775 25927 26781
rect 25869 26772 25881 26775
rect 25740 26744 25881 26772
rect 25740 26732 25746 26744
rect 25869 26741 25881 26744
rect 25915 26741 25927 26775
rect 25869 26735 25927 26741
rect 26786 26732 26792 26784
rect 26844 26772 26850 26784
rect 29196 26772 29224 26812
rect 29914 26800 29920 26812
rect 29972 26840 29978 26852
rect 30208 26849 30236 26880
rect 30745 26877 30757 26880
rect 30791 26877 30803 26911
rect 33060 26908 33088 26936
rect 33980 26908 34008 26939
rect 34146 26936 34152 26948
rect 34204 26936 34210 26988
rect 34606 26976 34612 26988
rect 34567 26948 34612 26976
rect 34606 26936 34612 26948
rect 34664 26936 34670 26988
rect 39873 26979 39931 26985
rect 39873 26945 39885 26979
rect 39919 26976 39931 26979
rect 40586 26976 40592 26988
rect 39919 26948 40592 26976
rect 39919 26945 39931 26948
rect 39873 26939 39931 26945
rect 40586 26936 40592 26948
rect 40644 26936 40650 26988
rect 33060 26880 34008 26908
rect 40129 26911 40187 26917
rect 30745 26871 30803 26877
rect 40129 26877 40141 26911
rect 40175 26877 40187 26911
rect 40129 26871 40187 26877
rect 30193 26843 30251 26849
rect 30193 26840 30205 26843
rect 29972 26812 30205 26840
rect 29972 26800 29978 26812
rect 30193 26809 30205 26812
rect 30239 26809 30251 26843
rect 30193 26803 30251 26809
rect 26844 26744 29224 26772
rect 29273 26775 29331 26781
rect 26844 26732 26850 26744
rect 29273 26741 29285 26775
rect 29319 26772 29331 26775
rect 29362 26772 29368 26784
rect 29319 26744 29368 26772
rect 29319 26741 29331 26744
rect 29273 26735 29331 26741
rect 29362 26732 29368 26744
rect 29420 26772 29426 26784
rect 30282 26772 30288 26784
rect 29420 26744 30288 26772
rect 29420 26732 29426 26744
rect 30282 26732 30288 26744
rect 30340 26732 30346 26784
rect 30466 26732 30472 26784
rect 30524 26772 30530 26784
rect 32585 26775 32643 26781
rect 32585 26772 32597 26775
rect 30524 26744 32597 26772
rect 30524 26732 30530 26744
rect 32585 26741 32597 26744
rect 32631 26741 32643 26775
rect 32585 26735 32643 26741
rect 33597 26775 33655 26781
rect 33597 26741 33609 26775
rect 33643 26772 33655 26775
rect 33962 26772 33968 26784
rect 33643 26744 33968 26772
rect 33643 26741 33655 26744
rect 33597 26735 33655 26741
rect 33962 26732 33968 26744
rect 34020 26732 34026 26784
rect 34790 26732 34796 26784
rect 34848 26772 34854 26784
rect 34977 26775 35035 26781
rect 34977 26772 34989 26775
rect 34848 26744 34989 26772
rect 34848 26732 34854 26744
rect 34977 26741 34989 26744
rect 35023 26741 35035 26775
rect 34977 26735 35035 26741
rect 36262 26732 36268 26784
rect 36320 26772 36326 26784
rect 38746 26772 38752 26784
rect 36320 26744 38752 26772
rect 36320 26732 36326 26744
rect 38746 26732 38752 26744
rect 38804 26732 38810 26784
rect 39942 26732 39948 26784
rect 40000 26772 40006 26784
rect 40144 26772 40172 26871
rect 58158 26772 58164 26784
rect 40000 26744 40172 26772
rect 58119 26744 58164 26772
rect 40000 26732 40006 26744
rect 58158 26732 58164 26744
rect 58216 26732 58222 26784
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 4706 26528 4712 26580
rect 4764 26568 4770 26580
rect 7193 26571 7251 26577
rect 7193 26568 7205 26571
rect 4764 26540 7205 26568
rect 4764 26528 4770 26540
rect 7193 26537 7205 26540
rect 7239 26537 7251 26571
rect 7193 26531 7251 26537
rect 7745 26571 7803 26577
rect 7745 26537 7757 26571
rect 7791 26568 7803 26571
rect 7926 26568 7932 26580
rect 7791 26540 7932 26568
rect 7791 26537 7803 26540
rect 7745 26531 7803 26537
rect 2869 26503 2927 26509
rect 2869 26469 2881 26503
rect 2915 26500 2927 26503
rect 4614 26500 4620 26512
rect 2915 26472 4620 26500
rect 2915 26469 2927 26472
rect 2869 26463 2927 26469
rect 4614 26460 4620 26472
rect 4672 26460 4678 26512
rect 3878 26392 3884 26444
rect 3936 26432 3942 26444
rect 7208 26432 7236 26531
rect 7926 26528 7932 26540
rect 7984 26528 7990 26580
rect 11606 26528 11612 26580
rect 11664 26568 11670 26580
rect 11885 26571 11943 26577
rect 11885 26568 11897 26571
rect 11664 26540 11897 26568
rect 11664 26528 11670 26540
rect 11885 26537 11897 26540
rect 11931 26537 11943 26571
rect 11885 26531 11943 26537
rect 12713 26571 12771 26577
rect 12713 26537 12725 26571
rect 12759 26568 12771 26571
rect 13814 26568 13820 26580
rect 12759 26540 13820 26568
rect 12759 26537 12771 26540
rect 12713 26531 12771 26537
rect 13814 26528 13820 26540
rect 13872 26528 13878 26580
rect 18693 26571 18751 26577
rect 14476 26540 18460 26568
rect 8110 26460 8116 26512
rect 8168 26460 8174 26512
rect 14476 26500 14504 26540
rect 8404 26472 14504 26500
rect 18432 26500 18460 26540
rect 18693 26537 18705 26571
rect 18739 26568 18751 26571
rect 19242 26568 19248 26580
rect 18739 26540 19248 26568
rect 18739 26537 18751 26540
rect 18693 26531 18751 26537
rect 19242 26528 19248 26540
rect 19300 26528 19306 26580
rect 20806 26528 20812 26580
rect 20864 26568 20870 26580
rect 22094 26568 22100 26580
rect 20864 26540 22100 26568
rect 20864 26528 20870 26540
rect 22094 26528 22100 26540
rect 22152 26528 22158 26580
rect 22572 26540 24440 26568
rect 22186 26500 22192 26512
rect 18432 26472 22192 26500
rect 8128 26432 8156 26460
rect 3936 26404 6776 26432
rect 7208 26404 8064 26432
rect 8128 26404 8248 26432
rect 3936 26392 3942 26404
rect 3050 26364 3056 26376
rect 3011 26336 3056 26364
rect 3050 26324 3056 26336
rect 3108 26324 3114 26376
rect 3234 26364 3240 26376
rect 3195 26336 3240 26364
rect 3234 26324 3240 26336
rect 3292 26324 3298 26376
rect 4062 26364 4068 26376
rect 4023 26336 4068 26364
rect 4062 26324 4068 26336
rect 4120 26324 4126 26376
rect 4172 26373 4200 26404
rect 6748 26376 6776 26404
rect 4157 26367 4215 26373
rect 4157 26333 4169 26367
rect 4203 26333 4215 26367
rect 4157 26327 4215 26333
rect 4249 26367 4307 26373
rect 4249 26333 4261 26367
rect 4295 26364 4307 26367
rect 4433 26367 4491 26373
rect 4295 26336 4384 26364
rect 4295 26333 4307 26336
rect 4249 26327 4307 26333
rect 3970 26256 3976 26308
rect 4028 26296 4034 26308
rect 4356 26296 4384 26336
rect 4433 26333 4445 26367
rect 4479 26364 4491 26367
rect 4706 26364 4712 26376
rect 4479 26336 4712 26364
rect 4479 26333 4491 26336
rect 4433 26327 4491 26333
rect 4706 26324 4712 26336
rect 4764 26364 4770 26376
rect 4764 26336 5120 26364
rect 4764 26324 4770 26336
rect 4028 26268 4384 26296
rect 4028 26256 4034 26268
rect 3786 26228 3792 26240
rect 3747 26200 3792 26228
rect 3786 26188 3792 26200
rect 3844 26188 3850 26240
rect 4893 26231 4951 26237
rect 4893 26197 4905 26231
rect 4939 26228 4951 26231
rect 5092 26228 5120 26336
rect 6730 26324 6736 26376
rect 6788 26364 6794 26376
rect 7558 26364 7564 26376
rect 6788 26336 7564 26364
rect 6788 26324 6794 26336
rect 7558 26324 7564 26336
rect 7616 26364 7622 26376
rect 8036 26373 8064 26404
rect 8220 26373 8248 26404
rect 8404 26376 8432 26472
rect 22186 26460 22192 26472
rect 22244 26460 22250 26512
rect 11057 26435 11115 26441
rect 11057 26401 11069 26435
rect 11103 26432 11115 26435
rect 12158 26432 12164 26444
rect 11103 26404 12164 26432
rect 11103 26401 11115 26404
rect 11057 26395 11115 26401
rect 12158 26392 12164 26404
rect 12216 26392 12222 26444
rect 17129 26435 17187 26441
rect 17129 26401 17141 26435
rect 17175 26432 17187 26435
rect 17218 26432 17224 26444
rect 17175 26404 17224 26432
rect 17175 26401 17187 26404
rect 17129 26395 17187 26401
rect 17218 26392 17224 26404
rect 17276 26392 17282 26444
rect 17862 26392 17868 26444
rect 17920 26432 17926 26444
rect 17920 26404 18184 26432
rect 17920 26392 17926 26404
rect 8021 26367 8079 26373
rect 7616 26336 7981 26364
rect 7616 26324 7622 26336
rect 5442 26256 5448 26308
rect 5500 26296 5506 26308
rect 7742 26296 7748 26308
rect 5500 26268 7748 26296
rect 5500 26256 5506 26268
rect 7742 26256 7748 26268
rect 7800 26256 7806 26308
rect 7953 26296 7981 26336
rect 8021 26333 8033 26367
rect 8067 26333 8079 26367
rect 8021 26327 8079 26333
rect 8113 26367 8171 26373
rect 8113 26333 8125 26367
rect 8159 26333 8171 26367
rect 8113 26327 8171 26333
rect 8205 26367 8263 26373
rect 8205 26333 8217 26367
rect 8251 26333 8263 26367
rect 8205 26327 8263 26333
rect 8128 26296 8156 26327
rect 8386 26324 8392 26376
rect 8444 26364 8450 26376
rect 11977 26367 12035 26373
rect 8444 26336 8537 26364
rect 8444 26324 8450 26336
rect 11977 26333 11989 26367
rect 12023 26364 12035 26367
rect 12434 26364 12440 26376
rect 12023 26336 12440 26364
rect 12023 26333 12035 26336
rect 11977 26327 12035 26333
rect 12434 26324 12440 26336
rect 12492 26324 12498 26376
rect 16301 26367 16359 26373
rect 16301 26333 16313 26367
rect 16347 26364 16359 26367
rect 16758 26364 16764 26376
rect 16347 26336 16764 26364
rect 16347 26333 16359 26336
rect 16301 26327 16359 26333
rect 16758 26324 16764 26336
rect 16816 26324 16822 26376
rect 16945 26367 17003 26373
rect 16945 26333 16957 26367
rect 16991 26333 17003 26367
rect 16945 26327 17003 26333
rect 9306 26296 9312 26308
rect 7953 26268 8156 26296
rect 9267 26268 9312 26296
rect 9306 26256 9312 26268
rect 9364 26256 9370 26308
rect 12618 26296 12624 26308
rect 12579 26268 12624 26296
rect 12618 26256 12624 26268
rect 12676 26256 12682 26308
rect 7006 26228 7012 26240
rect 4939 26200 7012 26228
rect 4939 26197 4951 26200
rect 4893 26191 4951 26197
rect 7006 26188 7012 26200
rect 7064 26188 7070 26240
rect 13998 26188 14004 26240
rect 14056 26228 14062 26240
rect 16666 26228 16672 26240
rect 14056 26200 16672 26228
rect 14056 26188 14062 26200
rect 16666 26188 16672 26200
rect 16724 26228 16730 26240
rect 16960 26228 16988 26327
rect 17954 26324 17960 26376
rect 18012 26364 18018 26376
rect 18049 26367 18107 26373
rect 18049 26364 18061 26367
rect 18012 26336 18061 26364
rect 18012 26324 18018 26336
rect 18049 26333 18061 26336
rect 18095 26333 18107 26367
rect 18156 26364 18184 26404
rect 18874 26392 18880 26444
rect 18932 26432 18938 26444
rect 20898 26432 20904 26444
rect 18932 26404 20904 26432
rect 18932 26392 18938 26404
rect 20898 26392 20904 26404
rect 20956 26392 20962 26444
rect 22572 26432 22600 26540
rect 24302 26500 24308 26512
rect 21100 26404 22600 26432
rect 22664 26472 24308 26500
rect 18212 26367 18270 26373
rect 18212 26364 18224 26367
rect 18156 26336 18224 26364
rect 18049 26327 18107 26333
rect 18212 26333 18224 26336
rect 18258 26333 18270 26367
rect 18212 26327 18270 26333
rect 18322 26324 18328 26376
rect 18380 26364 18386 26376
rect 18463 26367 18521 26373
rect 18380 26336 18425 26364
rect 18380 26324 18386 26336
rect 18463 26333 18475 26367
rect 18509 26364 18521 26367
rect 18509 26336 18644 26364
rect 18509 26333 18521 26336
rect 18463 26327 18521 26333
rect 18616 26296 18644 26336
rect 18690 26324 18696 26376
rect 18748 26364 18754 26376
rect 20806 26364 20812 26376
rect 18748 26336 20812 26364
rect 18748 26324 18754 26336
rect 20806 26324 20812 26336
rect 20864 26364 20870 26376
rect 20993 26367 21051 26373
rect 20993 26364 21005 26367
rect 20864 26336 21005 26364
rect 20864 26324 20870 26336
rect 20993 26333 21005 26336
rect 21039 26333 21051 26367
rect 20993 26327 21051 26333
rect 19337 26299 19395 26305
rect 19337 26296 19349 26299
rect 18616 26268 19349 26296
rect 19337 26265 19349 26268
rect 19383 26296 19395 26299
rect 21100 26296 21128 26404
rect 22664 26364 22692 26472
rect 24302 26460 24308 26472
rect 24360 26460 24366 26512
rect 24412 26500 24440 26540
rect 25038 26528 25044 26580
rect 25096 26568 25102 26580
rect 27801 26571 27859 26577
rect 27801 26568 27813 26571
rect 25096 26540 27813 26568
rect 25096 26528 25102 26540
rect 27801 26537 27813 26540
rect 27847 26537 27859 26571
rect 27801 26531 27859 26537
rect 25222 26500 25228 26512
rect 24412 26472 25228 26500
rect 25222 26460 25228 26472
rect 25280 26460 25286 26512
rect 24578 26392 24584 26444
rect 24636 26432 24642 26444
rect 25590 26432 25596 26444
rect 24636 26404 24808 26432
rect 25551 26404 25596 26432
rect 24636 26392 24642 26404
rect 19383 26268 21128 26296
rect 21192 26336 22692 26364
rect 22741 26367 22799 26373
rect 19383 26265 19395 26268
rect 19337 26259 19395 26265
rect 16724 26200 16988 26228
rect 16724 26188 16730 26200
rect 20898 26188 20904 26240
rect 20956 26228 20962 26240
rect 21192 26228 21220 26336
rect 22741 26333 22753 26367
rect 22787 26364 22799 26367
rect 23201 26367 23259 26373
rect 23201 26364 23213 26367
rect 22787 26336 23213 26364
rect 22787 26333 22799 26336
rect 22741 26327 22799 26333
rect 23201 26333 23213 26336
rect 23247 26333 23259 26367
rect 24486 26364 24492 26376
rect 24447 26336 24492 26364
rect 23201 26327 23259 26333
rect 22186 26256 22192 26308
rect 22244 26296 22250 26308
rect 23216 26296 23244 26327
rect 24486 26324 24492 26336
rect 24544 26324 24550 26376
rect 24670 26364 24676 26376
rect 24631 26336 24676 26364
rect 24670 26324 24676 26336
rect 24728 26324 24734 26376
rect 24780 26373 24808 26404
rect 25590 26392 25596 26404
rect 25648 26392 25654 26444
rect 28997 26435 29055 26441
rect 28997 26401 29009 26435
rect 29043 26432 29055 26435
rect 29362 26432 29368 26444
rect 29043 26404 29368 26432
rect 29043 26401 29055 26404
rect 28997 26395 29055 26401
rect 29362 26392 29368 26404
rect 29420 26432 29426 26444
rect 29549 26435 29607 26441
rect 29549 26432 29561 26435
rect 29420 26404 29561 26432
rect 29420 26392 29426 26404
rect 29549 26401 29561 26404
rect 29595 26432 29607 26435
rect 29730 26432 29736 26444
rect 29595 26404 29736 26432
rect 29595 26401 29607 26404
rect 29549 26395 29607 26401
rect 29730 26392 29736 26404
rect 29788 26392 29794 26444
rect 29822 26392 29828 26444
rect 29880 26432 29886 26444
rect 35986 26432 35992 26444
rect 29880 26404 33916 26432
rect 29880 26392 29886 26404
rect 24765 26367 24823 26373
rect 24765 26333 24777 26367
rect 24811 26333 24823 26367
rect 24765 26327 24823 26333
rect 24857 26367 24915 26373
rect 24857 26333 24869 26367
rect 24903 26364 24915 26367
rect 25222 26364 25228 26376
rect 24903 26336 25228 26364
rect 24903 26333 24915 26336
rect 24857 26327 24915 26333
rect 25222 26324 25228 26336
rect 25280 26324 25286 26376
rect 25792 26336 29224 26364
rect 25792 26296 25820 26336
rect 22244 26268 22784 26296
rect 23216 26268 25820 26296
rect 25860 26299 25918 26305
rect 22244 26256 22250 26268
rect 22756 26240 22784 26268
rect 25860 26265 25872 26299
rect 25906 26265 25918 26299
rect 27430 26296 27436 26308
rect 27391 26268 27436 26296
rect 25860 26259 25918 26265
rect 20956 26200 21220 26228
rect 20956 26188 20962 26200
rect 22738 26188 22744 26240
rect 22796 26188 22802 26240
rect 25133 26231 25191 26237
rect 25133 26197 25145 26231
rect 25179 26228 25191 26231
rect 25884 26228 25912 26259
rect 27430 26256 27436 26268
rect 27488 26256 27494 26308
rect 27617 26299 27675 26305
rect 27617 26265 27629 26299
rect 27663 26296 27675 26299
rect 28994 26296 29000 26308
rect 27663 26268 29000 26296
rect 27663 26265 27675 26268
rect 27617 26259 27675 26265
rect 28994 26256 29000 26268
rect 29052 26296 29058 26308
rect 29196 26296 29224 26336
rect 32582 26324 32588 26376
rect 32640 26364 32646 26376
rect 32640 26336 33088 26364
rect 32640 26324 32646 26336
rect 30374 26296 30380 26308
rect 29052 26268 29132 26296
rect 29196 26268 30380 26296
rect 29052 26256 29058 26268
rect 26970 26228 26976 26240
rect 25179 26200 25912 26228
rect 26931 26200 26976 26228
rect 25179 26197 25191 26200
rect 25133 26191 25191 26197
rect 26970 26188 26976 26200
rect 27028 26188 27034 26240
rect 29104 26228 29132 26268
rect 30374 26256 30380 26268
rect 30432 26296 30438 26308
rect 30834 26296 30840 26308
rect 30432 26268 30840 26296
rect 30432 26256 30438 26268
rect 30834 26256 30840 26268
rect 30892 26296 30898 26308
rect 31021 26299 31079 26305
rect 31021 26296 31033 26299
rect 30892 26268 31033 26296
rect 30892 26256 30898 26268
rect 31021 26265 31033 26268
rect 31067 26265 31079 26299
rect 31021 26259 31079 26265
rect 32769 26299 32827 26305
rect 32769 26265 32781 26299
rect 32815 26265 32827 26299
rect 33060 26296 33088 26336
rect 33134 26324 33140 26376
rect 33192 26364 33198 26376
rect 33410 26364 33416 26376
rect 33192 26336 33416 26364
rect 33192 26324 33198 26336
rect 33410 26324 33416 26336
rect 33468 26373 33474 26376
rect 33468 26367 33517 26373
rect 33468 26333 33471 26367
rect 33505 26333 33517 26367
rect 33468 26327 33517 26333
rect 33597 26367 33655 26373
rect 33597 26333 33609 26367
rect 33643 26333 33655 26367
rect 33597 26327 33655 26333
rect 33468 26324 33474 26327
rect 33612 26296 33640 26327
rect 33686 26324 33692 26376
rect 33744 26364 33750 26376
rect 33888 26373 33916 26404
rect 34716 26404 35992 26432
rect 34716 26373 34744 26404
rect 35986 26392 35992 26404
rect 36044 26392 36050 26444
rect 33873 26367 33931 26373
rect 33744 26336 33789 26364
rect 33744 26324 33750 26336
rect 33873 26333 33885 26367
rect 33919 26364 33931 26367
rect 34701 26367 34759 26373
rect 34701 26364 34713 26367
rect 33919 26336 34713 26364
rect 33919 26333 33931 26336
rect 33873 26327 33931 26333
rect 34701 26333 34713 26336
rect 34747 26333 34759 26367
rect 34701 26327 34759 26333
rect 34790 26324 34796 26376
rect 34848 26364 34854 26376
rect 34885 26367 34943 26373
rect 34885 26364 34897 26367
rect 34848 26336 34897 26364
rect 34848 26324 34854 26336
rect 34885 26333 34897 26336
rect 34931 26333 34943 26367
rect 34885 26327 34943 26333
rect 34977 26367 35035 26373
rect 34977 26333 34989 26367
rect 35023 26333 35035 26367
rect 34977 26327 35035 26333
rect 35069 26367 35127 26373
rect 35069 26333 35081 26367
rect 35115 26364 35127 26367
rect 35805 26367 35863 26373
rect 35805 26364 35817 26367
rect 35115 26336 35817 26364
rect 35115 26333 35127 26336
rect 35069 26327 35127 26333
rect 35805 26333 35817 26336
rect 35851 26333 35863 26367
rect 35805 26327 35863 26333
rect 34238 26296 34244 26308
rect 33060 26268 33548 26296
rect 33612 26268 34244 26296
rect 32769 26259 32827 26265
rect 29638 26228 29644 26240
rect 29104 26200 29644 26228
rect 29638 26188 29644 26200
rect 29696 26188 29702 26240
rect 32784 26228 32812 26259
rect 33042 26228 33048 26240
rect 32784 26200 33048 26228
rect 33042 26188 33048 26200
rect 33100 26188 33106 26240
rect 33226 26228 33232 26240
rect 33187 26200 33232 26228
rect 33226 26188 33232 26200
rect 33284 26188 33290 26240
rect 33520 26228 33548 26268
rect 34238 26256 34244 26268
rect 34296 26296 34302 26308
rect 34992 26296 35020 26327
rect 34296 26268 35020 26296
rect 34296 26256 34302 26268
rect 35084 26228 35112 26327
rect 38746 26324 38752 26376
rect 38804 26364 38810 26376
rect 40221 26367 40279 26373
rect 40221 26364 40233 26367
rect 38804 26336 40233 26364
rect 38804 26324 38810 26336
rect 40221 26333 40233 26336
rect 40267 26333 40279 26367
rect 40221 26327 40279 26333
rect 35345 26299 35403 26305
rect 35345 26265 35357 26299
rect 35391 26296 35403 26299
rect 36078 26296 36084 26308
rect 35391 26268 36084 26296
rect 35391 26265 35403 26268
rect 35345 26259 35403 26265
rect 36078 26256 36084 26268
rect 36136 26256 36142 26308
rect 37550 26256 37556 26308
rect 37608 26296 37614 26308
rect 40037 26299 40095 26305
rect 40037 26296 40049 26299
rect 37608 26268 40049 26296
rect 37608 26256 37614 26268
rect 40037 26265 40049 26268
rect 40083 26296 40095 26299
rect 40865 26299 40923 26305
rect 40865 26296 40877 26299
rect 40083 26268 40877 26296
rect 40083 26265 40095 26268
rect 40037 26259 40095 26265
rect 40865 26265 40877 26268
rect 40911 26265 40923 26299
rect 41046 26296 41052 26308
rect 41007 26268 41052 26296
rect 40865 26259 40923 26265
rect 41046 26256 41052 26268
rect 41104 26256 41110 26308
rect 40402 26228 40408 26240
rect 33520 26200 35112 26228
rect 40363 26200 40408 26228
rect 40402 26188 40408 26200
rect 40460 26188 40466 26240
rect 40494 26188 40500 26240
rect 40552 26228 40558 26240
rect 41233 26231 41291 26237
rect 41233 26228 41245 26231
rect 40552 26200 41245 26228
rect 40552 26188 40558 26200
rect 41233 26197 41245 26200
rect 41279 26197 41291 26231
rect 41233 26191 41291 26197
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 3602 25984 3608 26036
rect 3660 26024 3666 26036
rect 3881 26027 3939 26033
rect 3881 26024 3893 26027
rect 3660 25996 3893 26024
rect 3660 25984 3666 25996
rect 3881 25993 3893 25996
rect 3927 25993 3939 26027
rect 7466 26024 7472 26036
rect 7427 25996 7472 26024
rect 3881 25987 3939 25993
rect 7466 25984 7472 25996
rect 7524 25984 7530 26036
rect 8386 26024 8392 26036
rect 8347 25996 8392 26024
rect 8386 25984 8392 25996
rect 8444 25984 8450 26036
rect 17494 26024 17500 26036
rect 17455 25996 17500 26024
rect 17494 25984 17500 25996
rect 17552 25984 17558 26036
rect 17862 25984 17868 26036
rect 17920 26024 17926 26036
rect 18877 26027 18935 26033
rect 18877 26024 18889 26027
rect 17920 25996 18889 26024
rect 17920 25984 17926 25996
rect 18877 25993 18889 25996
rect 18923 25993 18935 26027
rect 22094 26024 22100 26036
rect 18877 25987 18935 25993
rect 18964 25996 22100 26024
rect 2768 25959 2826 25965
rect 2768 25925 2780 25959
rect 2814 25956 2826 25959
rect 3786 25956 3792 25968
rect 2814 25928 3792 25956
rect 2814 25925 2826 25928
rect 2768 25919 2826 25925
rect 3786 25916 3792 25928
rect 3844 25916 3850 25968
rect 5442 25956 5448 25968
rect 5403 25928 5448 25956
rect 5442 25916 5448 25928
rect 5500 25916 5506 25968
rect 5626 25956 5632 25968
rect 5587 25928 5632 25956
rect 5626 25916 5632 25928
rect 5684 25916 5690 25968
rect 7484 25956 7512 25984
rect 8849 25959 8907 25965
rect 8849 25956 8861 25959
rect 7484 25928 8861 25956
rect 2406 25848 2412 25900
rect 2464 25888 2470 25900
rect 2501 25891 2559 25897
rect 2501 25888 2513 25891
rect 2464 25860 2513 25888
rect 2464 25848 2470 25860
rect 2501 25857 2513 25860
rect 2547 25857 2559 25891
rect 2501 25851 2559 25857
rect 6086 25848 6092 25900
rect 6144 25888 6150 25900
rect 6546 25888 6552 25900
rect 6144 25860 6552 25888
rect 6144 25848 6150 25860
rect 6546 25848 6552 25860
rect 6604 25897 6610 25900
rect 6604 25891 6653 25897
rect 6604 25857 6607 25891
rect 6641 25857 6653 25891
rect 6604 25851 6653 25857
rect 6699 25851 6705 25903
rect 6757 25900 6763 25903
rect 6757 25894 6772 25900
rect 6760 25860 6772 25894
rect 6757 25854 6772 25860
rect 6830 25891 6888 25897
rect 6830 25857 6842 25891
rect 6876 25857 6888 25891
rect 6757 25851 6763 25854
rect 6830 25851 6888 25857
rect 6604 25848 6610 25851
rect 5813 25823 5871 25829
rect 5813 25789 5825 25823
rect 5859 25820 5871 25823
rect 6840 25820 6868 25851
rect 7006 25848 7012 25900
rect 7064 25888 7070 25900
rect 7484 25888 7512 25928
rect 8849 25925 8861 25928
rect 8895 25925 8907 25959
rect 8849 25919 8907 25925
rect 9033 25959 9091 25965
rect 9033 25925 9045 25959
rect 9079 25956 9091 25959
rect 9766 25956 9772 25968
rect 9079 25928 9772 25956
rect 9079 25925 9091 25928
rect 9033 25919 9091 25925
rect 9766 25916 9772 25928
rect 9824 25956 9830 25968
rect 10042 25956 10048 25968
rect 9824 25928 10048 25956
rect 9824 25916 9830 25928
rect 10042 25916 10048 25928
rect 10100 25916 10106 25968
rect 13906 25916 13912 25968
rect 13964 25956 13970 25968
rect 14277 25959 14335 25965
rect 14277 25956 14289 25959
rect 13964 25928 14289 25956
rect 13964 25916 13970 25928
rect 14277 25925 14289 25928
rect 14323 25925 14335 25959
rect 18322 25956 18328 25968
rect 14277 25919 14335 25925
rect 17877 25928 18328 25956
rect 7064 25860 7512 25888
rect 7064 25848 7070 25860
rect 9674 25848 9680 25900
rect 9732 25888 9738 25900
rect 9861 25891 9919 25897
rect 9861 25888 9873 25891
rect 9732 25860 9873 25888
rect 9732 25848 9738 25860
rect 9861 25857 9873 25860
rect 9907 25857 9919 25891
rect 9861 25851 9919 25857
rect 5859 25792 6868 25820
rect 5859 25789 5871 25792
rect 5813 25783 5871 25789
rect 9490 25780 9496 25832
rect 9548 25820 9554 25832
rect 9585 25823 9643 25829
rect 9585 25820 9597 25823
rect 9548 25792 9597 25820
rect 9548 25780 9554 25792
rect 9585 25789 9597 25792
rect 9631 25789 9643 25823
rect 10060 25820 10088 25916
rect 17877 25900 17905 25928
rect 18322 25916 18328 25928
rect 18380 25956 18386 25968
rect 18964 25956 18992 25996
rect 22094 25984 22100 25996
rect 22152 25984 22158 26036
rect 25133 26027 25191 26033
rect 25133 25993 25145 26027
rect 25179 26024 25191 26027
rect 25222 26024 25228 26036
rect 25179 25996 25228 26024
rect 25179 25993 25191 25996
rect 25133 25987 25191 25993
rect 25222 25984 25228 25996
rect 25280 25984 25286 26036
rect 26237 26027 26295 26033
rect 26237 25993 26249 26027
rect 26283 26024 26295 26027
rect 27982 26024 27988 26036
rect 26283 25996 27988 26024
rect 26283 25993 26295 25996
rect 26237 25987 26295 25993
rect 27982 25984 27988 25996
rect 28040 25984 28046 26036
rect 30834 26024 30840 26036
rect 30795 25996 30840 26024
rect 30834 25984 30840 25996
rect 30892 25984 30898 26036
rect 32677 26027 32735 26033
rect 32677 25993 32689 26027
rect 32723 26024 32735 26027
rect 33134 26024 33140 26036
rect 32723 25996 33140 26024
rect 32723 25993 32735 25996
rect 32677 25987 32735 25993
rect 33134 25984 33140 25996
rect 33192 25984 33198 26036
rect 34514 25984 34520 26036
rect 34572 26024 34578 26036
rect 34977 26027 35035 26033
rect 34977 26024 34989 26027
rect 34572 25996 34989 26024
rect 34572 25984 34578 25996
rect 34977 25993 34989 25996
rect 35023 25993 35035 26027
rect 34977 25987 35035 25993
rect 39942 25984 39948 26036
rect 40000 25984 40006 26036
rect 40586 26024 40592 26036
rect 40547 25996 40592 26024
rect 40586 25984 40592 25996
rect 40644 25984 40650 26036
rect 18380 25928 18992 25956
rect 19061 25959 19119 25965
rect 18380 25916 18386 25928
rect 19061 25925 19073 25959
rect 19107 25956 19119 25959
rect 20622 25956 20628 25968
rect 19107 25928 20628 25956
rect 19107 25925 19119 25928
rect 19061 25919 19119 25925
rect 20622 25916 20628 25928
rect 20680 25916 20686 25968
rect 20901 25959 20959 25965
rect 20901 25925 20913 25959
rect 20947 25956 20959 25959
rect 20990 25956 20996 25968
rect 20947 25928 20996 25956
rect 20947 25925 20959 25928
rect 20901 25919 20959 25925
rect 11701 25891 11759 25897
rect 11701 25857 11713 25891
rect 11747 25888 11759 25891
rect 11747 25860 12434 25888
rect 11747 25857 11759 25860
rect 11701 25851 11759 25857
rect 11977 25823 12035 25829
rect 11977 25820 11989 25823
rect 10060 25792 11989 25820
rect 9585 25783 9643 25789
rect 11977 25789 11989 25792
rect 12023 25789 12035 25823
rect 12406 25820 12434 25860
rect 12986 25848 12992 25900
rect 13044 25888 13050 25900
rect 13817 25891 13875 25897
rect 13817 25888 13829 25891
rect 13044 25860 13829 25888
rect 13044 25848 13050 25860
rect 13817 25857 13829 25860
rect 13863 25888 13875 25891
rect 14461 25891 14519 25897
rect 14461 25888 14473 25891
rect 13863 25860 14473 25888
rect 13863 25857 13875 25860
rect 13817 25851 13875 25857
rect 14461 25857 14473 25860
rect 14507 25857 14519 25891
rect 14461 25851 14519 25857
rect 15841 25891 15899 25897
rect 15841 25857 15853 25891
rect 15887 25888 15899 25891
rect 16574 25888 16580 25900
rect 15887 25860 16580 25888
rect 15887 25857 15899 25860
rect 15841 25851 15899 25857
rect 16574 25848 16580 25860
rect 16632 25848 16638 25900
rect 16853 25891 16911 25897
rect 16853 25857 16865 25891
rect 16899 25888 16911 25891
rect 17218 25888 17224 25900
rect 16899 25860 17224 25888
rect 16899 25857 16911 25860
rect 16853 25851 16911 25857
rect 17218 25848 17224 25860
rect 17276 25848 17282 25900
rect 17678 25848 17684 25900
rect 17736 25888 17742 25900
rect 17773 25891 17831 25897
rect 17773 25888 17785 25891
rect 17736 25860 17785 25888
rect 17736 25848 17742 25860
rect 17773 25857 17785 25860
rect 17819 25857 17831 25891
rect 17773 25851 17831 25857
rect 17862 25894 17920 25900
rect 17862 25860 17874 25894
rect 17908 25860 17920 25894
rect 17862 25854 17920 25860
rect 17957 25891 18015 25897
rect 17957 25857 17969 25891
rect 18003 25857 18015 25891
rect 17957 25851 18015 25857
rect 18141 25891 18199 25897
rect 18141 25857 18153 25891
rect 18187 25888 18199 25891
rect 18874 25888 18880 25900
rect 18187 25860 18880 25888
rect 18187 25857 18199 25860
rect 18141 25851 18199 25857
rect 12406 25792 13124 25820
rect 11977 25783 12035 25789
rect 9600 25752 9628 25783
rect 12618 25752 12624 25764
rect 9600 25724 12624 25752
rect 12618 25712 12624 25724
rect 12676 25712 12682 25764
rect 4154 25644 4160 25696
rect 4212 25684 4218 25696
rect 4617 25687 4675 25693
rect 4617 25684 4629 25687
rect 4212 25656 4629 25684
rect 4212 25644 4218 25656
rect 4617 25653 4629 25656
rect 4663 25684 4675 25687
rect 4982 25684 4988 25696
rect 4663 25656 4988 25684
rect 4663 25653 4675 25656
rect 4617 25647 4675 25653
rect 4982 25644 4988 25656
rect 5040 25644 5046 25696
rect 6365 25687 6423 25693
rect 6365 25653 6377 25687
rect 6411 25684 6423 25687
rect 6454 25684 6460 25696
rect 6411 25656 6460 25684
rect 6411 25653 6423 25656
rect 6365 25647 6423 25653
rect 6454 25644 6460 25656
rect 6512 25644 6518 25696
rect 9030 25644 9036 25696
rect 9088 25684 9094 25696
rect 12986 25684 12992 25696
rect 9088 25656 12992 25684
rect 9088 25644 9094 25656
rect 12986 25644 12992 25656
rect 13044 25644 13050 25696
rect 13096 25693 13124 25792
rect 15102 25780 15108 25832
rect 15160 25820 15166 25832
rect 15565 25823 15623 25829
rect 15565 25820 15577 25823
rect 15160 25792 15577 25820
rect 15160 25780 15166 25792
rect 15565 25789 15577 25792
rect 15611 25789 15623 25823
rect 15565 25783 15623 25789
rect 13081 25687 13139 25693
rect 13081 25653 13093 25687
rect 13127 25684 13139 25687
rect 14182 25684 14188 25696
rect 13127 25656 14188 25684
rect 13127 25653 13139 25656
rect 13081 25647 13139 25653
rect 14182 25644 14188 25656
rect 14240 25644 14246 25696
rect 15286 25644 15292 25696
rect 15344 25684 15350 25696
rect 16669 25687 16727 25693
rect 16669 25684 16681 25687
rect 15344 25656 16681 25684
rect 15344 25644 15350 25656
rect 16669 25653 16681 25656
rect 16715 25653 16727 25687
rect 17788 25684 17816 25851
rect 17972 25820 18000 25851
rect 18874 25848 18880 25860
rect 18932 25848 18938 25900
rect 19150 25848 19156 25900
rect 19208 25888 19214 25900
rect 19245 25891 19303 25897
rect 19245 25888 19257 25891
rect 19208 25860 19257 25888
rect 19208 25848 19214 25860
rect 19245 25857 19257 25860
rect 19291 25888 19303 25891
rect 19889 25891 19947 25897
rect 19291 25860 19840 25888
rect 19291 25857 19303 25860
rect 19245 25851 19303 25857
rect 19705 25823 19763 25829
rect 19705 25820 19717 25823
rect 17972 25792 19717 25820
rect 19705 25789 19717 25792
rect 19751 25789 19763 25823
rect 19812 25820 19840 25860
rect 19889 25857 19901 25891
rect 19935 25888 19947 25891
rect 19978 25888 19984 25900
rect 19935 25860 19984 25888
rect 19935 25857 19947 25860
rect 19889 25851 19947 25857
rect 19978 25848 19984 25860
rect 20036 25848 20042 25900
rect 20073 25891 20131 25897
rect 20073 25857 20085 25891
rect 20119 25888 20131 25891
rect 20916 25888 20944 25919
rect 20990 25916 20996 25928
rect 21048 25916 21054 25968
rect 21269 25959 21327 25965
rect 21269 25925 21281 25959
rect 21315 25956 21327 25959
rect 21315 25928 22784 25956
rect 21315 25925 21327 25928
rect 21269 25919 21327 25925
rect 20119 25860 20944 25888
rect 21085 25891 21143 25897
rect 20119 25857 20131 25860
rect 20073 25851 20131 25857
rect 21085 25857 21097 25891
rect 21131 25888 21143 25891
rect 22186 25888 22192 25900
rect 21131 25860 22192 25888
rect 21131 25857 21143 25860
rect 21085 25851 21143 25857
rect 20088 25820 20116 25851
rect 22186 25848 22192 25860
rect 22244 25848 22250 25900
rect 22756 25897 22784 25928
rect 24578 25916 24584 25968
rect 24636 25956 24642 25968
rect 24636 25928 25912 25956
rect 24636 25916 24642 25928
rect 25884 25900 25912 25928
rect 26878 25916 26884 25968
rect 26936 25956 26942 25968
rect 26973 25959 27031 25965
rect 26973 25956 26985 25959
rect 26936 25928 26985 25956
rect 26936 25916 26942 25928
rect 26973 25925 26985 25928
rect 27019 25925 27031 25959
rect 26973 25919 27031 25925
rect 33226 25916 33232 25968
rect 33284 25956 33290 25968
rect 33382 25959 33440 25965
rect 33382 25956 33394 25959
rect 33284 25928 33394 25956
rect 33284 25916 33290 25928
rect 33382 25925 33394 25928
rect 33428 25925 33440 25959
rect 33382 25919 33440 25925
rect 36078 25916 36084 25968
rect 36136 25965 36142 25968
rect 36136 25956 36148 25965
rect 36136 25928 36181 25956
rect 36136 25919 36148 25928
rect 36136 25916 36142 25919
rect 38654 25916 38660 25968
rect 38712 25956 38718 25968
rect 39960 25956 39988 25984
rect 38712 25928 40172 25956
rect 38712 25916 38718 25928
rect 22557 25891 22615 25897
rect 22557 25857 22569 25891
rect 22603 25857 22615 25891
rect 22557 25851 22615 25857
rect 22741 25891 22799 25897
rect 22741 25857 22753 25891
rect 22787 25857 22799 25891
rect 22741 25851 22799 25857
rect 22833 25891 22891 25897
rect 22833 25857 22845 25891
rect 22879 25857 22891 25891
rect 22833 25851 22891 25857
rect 22925 25891 22983 25897
rect 22925 25857 22937 25891
rect 22971 25888 22983 25891
rect 23661 25891 23719 25897
rect 23661 25888 23673 25891
rect 22971 25860 23673 25888
rect 22971 25857 22983 25860
rect 22925 25851 22983 25857
rect 23661 25857 23673 25860
rect 23707 25857 23719 25891
rect 23661 25851 23719 25857
rect 22572 25820 22600 25851
rect 19812 25792 20116 25820
rect 22020 25792 22600 25820
rect 19705 25783 19763 25789
rect 18874 25712 18880 25764
rect 18932 25752 18938 25764
rect 21818 25752 21824 25764
rect 18932 25724 21824 25752
rect 18932 25712 18938 25724
rect 21818 25712 21824 25724
rect 21876 25752 21882 25764
rect 22020 25752 22048 25792
rect 21876 25724 22048 25752
rect 21876 25712 21882 25724
rect 22094 25712 22100 25764
rect 22152 25752 22158 25764
rect 22848 25752 22876 25851
rect 23676 25820 23704 25851
rect 24486 25848 24492 25900
rect 24544 25888 24550 25900
rect 25774 25897 25780 25900
rect 25593 25891 25651 25897
rect 25593 25888 25605 25891
rect 24544 25860 25605 25888
rect 24544 25848 24550 25860
rect 25593 25857 25605 25860
rect 25639 25857 25651 25891
rect 25772 25888 25780 25897
rect 25735 25860 25780 25888
rect 25593 25851 25651 25857
rect 25772 25851 25780 25860
rect 25774 25848 25780 25851
rect 25832 25848 25838 25900
rect 25866 25848 25872 25900
rect 25924 25888 25930 25900
rect 26007 25891 26065 25897
rect 25924 25860 25969 25888
rect 25924 25848 25930 25860
rect 26007 25857 26019 25891
rect 26053 25888 26065 25891
rect 26896 25888 26924 25916
rect 26053 25860 26924 25888
rect 26053 25857 26065 25860
rect 26007 25851 26065 25857
rect 26166 25820 26194 25860
rect 28994 25848 29000 25900
rect 29052 25888 29058 25900
rect 29282 25891 29340 25897
rect 29282 25888 29294 25891
rect 29052 25860 29294 25888
rect 29052 25848 29058 25860
rect 29282 25857 29294 25860
rect 29328 25857 29340 25891
rect 29282 25851 29340 25857
rect 29549 25891 29607 25897
rect 29549 25857 29561 25891
rect 29595 25888 29607 25891
rect 30926 25888 30932 25900
rect 29595 25860 30932 25888
rect 29595 25857 29607 25860
rect 29549 25851 29607 25857
rect 30926 25848 30932 25860
rect 30984 25848 30990 25900
rect 33042 25848 33048 25900
rect 33100 25888 33106 25900
rect 33137 25891 33195 25897
rect 33137 25888 33149 25891
rect 33100 25860 33149 25888
rect 33100 25848 33106 25860
rect 33137 25857 33149 25860
rect 33183 25857 33195 25891
rect 33137 25851 33195 25857
rect 39873 25891 39931 25897
rect 39873 25857 39885 25891
rect 39919 25888 39931 25891
rect 40034 25888 40040 25900
rect 39919 25860 40040 25888
rect 39919 25857 39931 25860
rect 39873 25851 39931 25857
rect 40034 25848 40040 25860
rect 40092 25848 40098 25900
rect 40144 25897 40172 25928
rect 40402 25916 40408 25968
rect 40460 25956 40466 25968
rect 40460 25928 41092 25956
rect 40460 25916 40466 25928
rect 40129 25891 40187 25897
rect 40129 25857 40141 25891
rect 40175 25857 40187 25891
rect 40862 25888 40868 25900
rect 40823 25860 40868 25888
rect 40129 25851 40187 25857
rect 40862 25848 40868 25860
rect 40920 25848 40926 25900
rect 41064 25897 41092 25928
rect 40957 25891 41015 25897
rect 40957 25857 40969 25891
rect 41003 25857 41015 25891
rect 40957 25851 41015 25857
rect 41049 25891 41107 25897
rect 41049 25857 41061 25891
rect 41095 25857 41107 25891
rect 41049 25851 41107 25857
rect 41233 25891 41291 25897
rect 41233 25857 41245 25891
rect 41279 25857 41291 25891
rect 41233 25851 41291 25857
rect 36354 25820 36360 25832
rect 23676 25792 26194 25820
rect 36315 25792 36360 25820
rect 36354 25780 36360 25792
rect 36412 25780 36418 25832
rect 40586 25780 40592 25832
rect 40644 25820 40650 25832
rect 40972 25820 41000 25851
rect 40644 25792 41000 25820
rect 40644 25780 40650 25792
rect 22152 25724 22876 25752
rect 22152 25712 22158 25724
rect 40954 25712 40960 25764
rect 41012 25752 41018 25764
rect 41248 25752 41276 25851
rect 41012 25724 41276 25752
rect 41012 25712 41018 25724
rect 20990 25684 20996 25696
rect 17788 25656 20996 25684
rect 16669 25647 16727 25653
rect 20990 25644 20996 25656
rect 21048 25644 21054 25696
rect 23198 25684 23204 25696
rect 23159 25656 23204 25684
rect 23198 25644 23204 25656
rect 23256 25644 23262 25696
rect 28166 25684 28172 25696
rect 28127 25656 28172 25684
rect 28166 25644 28172 25656
rect 28224 25644 28230 25696
rect 33318 25644 33324 25696
rect 33376 25684 33382 25696
rect 34517 25687 34575 25693
rect 34517 25684 34529 25687
rect 33376 25656 34529 25684
rect 33376 25644 33382 25656
rect 34517 25653 34529 25656
rect 34563 25653 34575 25687
rect 34517 25647 34575 25653
rect 38749 25687 38807 25693
rect 38749 25653 38761 25687
rect 38795 25684 38807 25687
rect 38838 25684 38844 25696
rect 38795 25656 38844 25684
rect 38795 25653 38807 25656
rect 38749 25647 38807 25653
rect 38838 25644 38844 25656
rect 38896 25684 38902 25696
rect 41046 25684 41052 25696
rect 38896 25656 41052 25684
rect 38896 25644 38902 25656
rect 41046 25644 41052 25656
rect 41104 25644 41110 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 5353 25483 5411 25489
rect 5353 25449 5365 25483
rect 5399 25480 5411 25483
rect 5626 25480 5632 25492
rect 5399 25452 5632 25480
rect 5399 25449 5411 25452
rect 5353 25443 5411 25449
rect 5626 25440 5632 25452
rect 5684 25440 5690 25492
rect 6546 25440 6552 25492
rect 6604 25480 6610 25492
rect 7193 25483 7251 25489
rect 7193 25480 7205 25483
rect 6604 25452 7205 25480
rect 6604 25440 6610 25452
rect 7193 25449 7205 25452
rect 7239 25449 7251 25483
rect 7193 25443 7251 25449
rect 21450 25440 21456 25492
rect 21508 25480 21514 25492
rect 23566 25480 23572 25492
rect 21508 25452 23572 25480
rect 21508 25440 21514 25452
rect 23566 25440 23572 25452
rect 23624 25480 23630 25492
rect 24118 25480 24124 25492
rect 23624 25452 24124 25480
rect 23624 25440 23630 25452
rect 24118 25440 24124 25452
rect 24176 25440 24182 25492
rect 24854 25440 24860 25492
rect 24912 25480 24918 25492
rect 25593 25483 25651 25489
rect 25593 25480 25605 25483
rect 24912 25452 25605 25480
rect 24912 25440 24918 25452
rect 25593 25449 25605 25452
rect 25639 25449 25651 25483
rect 25593 25443 25651 25449
rect 37642 25440 37648 25492
rect 37700 25480 37706 25492
rect 38105 25483 38163 25489
rect 38105 25480 38117 25483
rect 37700 25452 38117 25480
rect 37700 25440 37706 25452
rect 38105 25449 38117 25452
rect 38151 25480 38163 25483
rect 38286 25480 38292 25492
rect 38151 25452 38292 25480
rect 38151 25449 38163 25452
rect 38105 25443 38163 25449
rect 38286 25440 38292 25452
rect 38344 25440 38350 25492
rect 40034 25480 40040 25492
rect 39995 25452 40040 25480
rect 40034 25440 40040 25452
rect 40092 25440 40098 25492
rect 8386 25372 8392 25424
rect 8444 25412 8450 25424
rect 9125 25415 9183 25421
rect 9125 25412 9137 25415
rect 8444 25384 9137 25412
rect 8444 25372 8450 25384
rect 9125 25381 9137 25384
rect 9171 25381 9183 25415
rect 9125 25375 9183 25381
rect 11149 25415 11207 25421
rect 11149 25381 11161 25415
rect 11195 25412 11207 25415
rect 11698 25412 11704 25424
rect 11195 25384 11704 25412
rect 11195 25381 11207 25384
rect 11149 25375 11207 25381
rect 11698 25372 11704 25384
rect 11756 25372 11762 25424
rect 25222 25372 25228 25424
rect 25280 25412 25286 25424
rect 29178 25412 29184 25424
rect 25280 25384 29184 25412
rect 25280 25372 25286 25384
rect 29178 25372 29184 25384
rect 29236 25372 29242 25424
rect 3878 25304 3884 25356
rect 3936 25344 3942 25356
rect 4614 25344 4620 25356
rect 3936 25316 4200 25344
rect 3936 25304 3942 25316
rect 2866 25236 2872 25288
rect 2924 25276 2930 25288
rect 4062 25276 4068 25288
rect 2924 25248 4068 25276
rect 2924 25236 2930 25248
rect 4062 25236 4068 25248
rect 4120 25236 4126 25288
rect 4172 25285 4200 25316
rect 4356 25316 4620 25344
rect 4157 25279 4215 25285
rect 4157 25245 4169 25279
rect 4203 25245 4215 25279
rect 4157 25239 4215 25245
rect 4249 25279 4307 25285
rect 4249 25245 4261 25279
rect 4295 25276 4307 25279
rect 4356 25276 4384 25316
rect 4614 25304 4620 25316
rect 4672 25304 4678 25356
rect 6733 25347 6791 25353
rect 6733 25313 6745 25347
rect 6779 25344 6791 25347
rect 8202 25344 8208 25356
rect 6779 25316 8208 25344
rect 6779 25313 6791 25316
rect 6733 25307 6791 25313
rect 8202 25304 8208 25316
rect 8260 25304 8266 25356
rect 16666 25304 16672 25356
rect 16724 25344 16730 25356
rect 18141 25347 18199 25353
rect 18141 25344 18153 25347
rect 16724 25316 18153 25344
rect 16724 25304 16730 25316
rect 18141 25313 18153 25316
rect 18187 25313 18199 25347
rect 18141 25307 18199 25313
rect 18417 25347 18475 25353
rect 18417 25313 18429 25347
rect 18463 25344 18475 25347
rect 19242 25344 19248 25356
rect 18463 25316 19248 25344
rect 18463 25313 18475 25316
rect 18417 25307 18475 25313
rect 19242 25304 19248 25316
rect 19300 25304 19306 25356
rect 22922 25344 22928 25356
rect 22883 25316 22928 25344
rect 22922 25304 22928 25316
rect 22980 25304 22986 25356
rect 32309 25347 32367 25353
rect 32309 25313 32321 25347
rect 32355 25344 32367 25347
rect 33042 25344 33048 25356
rect 32355 25316 33048 25344
rect 32355 25313 32367 25316
rect 32309 25307 32367 25313
rect 4295 25248 4384 25276
rect 4433 25279 4491 25285
rect 4295 25245 4307 25248
rect 4249 25239 4307 25245
rect 4433 25245 4445 25279
rect 4479 25276 4491 25279
rect 4706 25276 4712 25288
rect 4479 25248 4712 25276
rect 4479 25245 4491 25248
rect 4433 25239 4491 25245
rect 4706 25236 4712 25248
rect 4764 25236 4770 25288
rect 6454 25236 6460 25288
rect 6512 25285 6518 25288
rect 6512 25276 6524 25285
rect 9309 25279 9367 25285
rect 6512 25248 6557 25276
rect 6512 25239 6524 25248
rect 9309 25245 9321 25279
rect 9355 25276 9367 25279
rect 9766 25276 9772 25288
rect 9355 25248 9772 25276
rect 9355 25245 9367 25248
rect 9309 25239 9367 25245
rect 6512 25236 6518 25239
rect 9766 25236 9772 25248
rect 9824 25236 9830 25288
rect 9861 25279 9919 25285
rect 9861 25245 9873 25279
rect 9907 25276 9919 25279
rect 13722 25276 13728 25288
rect 9907 25248 13728 25276
rect 9907 25245 9919 25248
rect 9861 25239 9919 25245
rect 13722 25236 13728 25248
rect 13780 25276 13786 25288
rect 15286 25276 15292 25288
rect 13780 25248 15292 25276
rect 13780 25236 13786 25248
rect 15286 25236 15292 25248
rect 15344 25236 15350 25288
rect 17770 25276 17776 25288
rect 16960 25248 17776 25276
rect 10042 25208 10048 25220
rect 10003 25180 10048 25208
rect 10042 25168 10048 25180
rect 10100 25168 10106 25220
rect 10965 25211 11023 25217
rect 10965 25208 10977 25211
rect 10152 25180 10977 25208
rect 3602 25100 3608 25152
rect 3660 25140 3666 25152
rect 3789 25143 3847 25149
rect 3789 25140 3801 25143
rect 3660 25112 3801 25140
rect 3660 25100 3666 25112
rect 3789 25109 3801 25112
rect 3835 25109 3847 25143
rect 3789 25103 3847 25109
rect 9950 25100 9956 25152
rect 10008 25140 10014 25152
rect 10152 25140 10180 25180
rect 10965 25177 10977 25180
rect 11011 25177 11023 25211
rect 15105 25211 15163 25217
rect 10965 25171 11023 25177
rect 14384 25180 15056 25208
rect 10008 25112 10180 25140
rect 10229 25143 10287 25149
rect 10008 25100 10014 25112
rect 10229 25109 10241 25143
rect 10275 25140 10287 25143
rect 10686 25140 10692 25152
rect 10275 25112 10692 25140
rect 10275 25109 10287 25112
rect 10229 25103 10287 25109
rect 10686 25100 10692 25112
rect 10744 25100 10750 25152
rect 12710 25100 12716 25152
rect 12768 25140 12774 25152
rect 13446 25140 13452 25152
rect 12768 25112 13452 25140
rect 12768 25100 12774 25112
rect 13446 25100 13452 25112
rect 13504 25100 13510 25152
rect 14182 25100 14188 25152
rect 14240 25140 14246 25152
rect 14384 25149 14412 25180
rect 14369 25143 14427 25149
rect 14369 25140 14381 25143
rect 14240 25112 14381 25140
rect 14240 25100 14246 25112
rect 14369 25109 14381 25112
rect 14415 25109 14427 25143
rect 14369 25103 14427 25109
rect 14734 25100 14740 25152
rect 14792 25140 14798 25152
rect 14921 25143 14979 25149
rect 14921 25140 14933 25143
rect 14792 25112 14933 25140
rect 14792 25100 14798 25112
rect 14921 25109 14933 25112
rect 14967 25109 14979 25143
rect 15028 25140 15056 25180
rect 15105 25177 15117 25211
rect 15151 25208 15163 25211
rect 15194 25208 15200 25220
rect 15151 25180 15200 25208
rect 15151 25177 15163 25180
rect 15105 25171 15163 25177
rect 15194 25168 15200 25180
rect 15252 25168 15258 25220
rect 16025 25211 16083 25217
rect 16025 25177 16037 25211
rect 16071 25177 16083 25211
rect 16025 25171 16083 25177
rect 16209 25211 16267 25217
rect 16209 25177 16221 25211
rect 16255 25208 16267 25211
rect 16666 25208 16672 25220
rect 16255 25180 16672 25208
rect 16255 25177 16267 25180
rect 16209 25171 16267 25177
rect 16040 25140 16068 25171
rect 16666 25168 16672 25180
rect 16724 25208 16730 25220
rect 16960 25217 16988 25248
rect 17770 25236 17776 25248
rect 17828 25236 17834 25288
rect 22669 25279 22727 25285
rect 22669 25245 22681 25279
rect 22715 25276 22727 25279
rect 23198 25276 23204 25288
rect 22715 25248 23204 25276
rect 22715 25245 22727 25248
rect 22669 25239 22727 25245
rect 23198 25236 23204 25248
rect 23256 25236 23262 25288
rect 25777 25279 25835 25285
rect 25777 25245 25789 25279
rect 25823 25276 25835 25279
rect 26970 25276 26976 25288
rect 25823 25248 26976 25276
rect 25823 25245 25835 25248
rect 25777 25239 25835 25245
rect 26970 25236 26976 25248
rect 27028 25236 27034 25288
rect 30926 25236 30932 25288
rect 30984 25276 30990 25288
rect 32324 25276 32352 25307
rect 33042 25304 33048 25316
rect 33100 25304 33106 25356
rect 30984 25248 32352 25276
rect 30984 25236 30990 25248
rect 36354 25236 36360 25288
rect 36412 25276 36418 25288
rect 37369 25279 37427 25285
rect 37369 25276 37381 25279
rect 36412 25248 37381 25276
rect 36412 25236 36418 25248
rect 37369 25245 37381 25248
rect 37415 25276 37427 25279
rect 38654 25276 38660 25288
rect 37415 25248 38660 25276
rect 37415 25245 37427 25248
rect 37369 25239 37427 25245
rect 38654 25236 38660 25248
rect 38712 25236 38718 25288
rect 40313 25279 40371 25285
rect 40313 25276 40325 25279
rect 39224 25248 40325 25276
rect 16945 25211 17003 25217
rect 16945 25208 16957 25211
rect 16724 25180 16957 25208
rect 16724 25168 16730 25180
rect 16945 25177 16957 25180
rect 16991 25177 17003 25211
rect 16945 25171 17003 25177
rect 17129 25211 17187 25217
rect 17129 25177 17141 25211
rect 17175 25208 17187 25211
rect 17310 25208 17316 25220
rect 17175 25180 17316 25208
rect 17175 25177 17187 25180
rect 17129 25171 17187 25177
rect 17310 25168 17316 25180
rect 17368 25208 17374 25220
rect 24486 25208 24492 25220
rect 17368 25180 24492 25208
rect 17368 25168 17374 25180
rect 24486 25168 24492 25180
rect 24544 25168 24550 25220
rect 25958 25208 25964 25220
rect 25919 25180 25964 25208
rect 25958 25168 25964 25180
rect 26016 25208 26022 25220
rect 27430 25208 27436 25220
rect 26016 25180 27436 25208
rect 26016 25168 26022 25180
rect 27430 25168 27436 25180
rect 27488 25168 27494 25220
rect 28258 25168 28264 25220
rect 28316 25208 28322 25220
rect 29641 25211 29699 25217
rect 29641 25208 29653 25211
rect 28316 25180 29653 25208
rect 28316 25168 28322 25180
rect 29641 25177 29653 25180
rect 29687 25177 29699 25211
rect 29641 25171 29699 25177
rect 29825 25211 29883 25217
rect 29825 25177 29837 25211
rect 29871 25208 29883 25211
rect 29871 25180 30972 25208
rect 29871 25177 29883 25180
rect 29825 25171 29883 25177
rect 15028 25112 16068 25140
rect 14921 25103 14979 25109
rect 17402 25100 17408 25152
rect 17460 25140 17466 25152
rect 17954 25140 17960 25152
rect 17460 25112 17960 25140
rect 17460 25100 17466 25112
rect 17954 25100 17960 25112
rect 18012 25100 18018 25152
rect 21545 25143 21603 25149
rect 21545 25109 21557 25143
rect 21591 25140 21603 25143
rect 22186 25140 22192 25152
rect 21591 25112 22192 25140
rect 21591 25109 21603 25112
rect 21545 25103 21603 25109
rect 22186 25100 22192 25112
rect 22244 25140 22250 25152
rect 23014 25140 23020 25152
rect 22244 25112 23020 25140
rect 22244 25100 22250 25112
rect 23014 25100 23020 25112
rect 23072 25100 23078 25152
rect 29086 25100 29092 25152
rect 29144 25140 29150 25152
rect 29840 25140 29868 25171
rect 29144 25112 29868 25140
rect 30009 25143 30067 25149
rect 29144 25100 29150 25112
rect 30009 25109 30021 25143
rect 30055 25140 30067 25143
rect 30282 25140 30288 25152
rect 30055 25112 30288 25140
rect 30055 25109 30067 25112
rect 30009 25103 30067 25109
rect 30282 25100 30288 25112
rect 30340 25100 30346 25152
rect 30944 25149 30972 25180
rect 31754 25168 31760 25220
rect 31812 25208 31818 25220
rect 32042 25211 32100 25217
rect 32042 25208 32054 25211
rect 31812 25180 32054 25208
rect 31812 25168 31818 25180
rect 32042 25177 32054 25180
rect 32088 25177 32100 25211
rect 32042 25171 32100 25177
rect 37124 25211 37182 25217
rect 37124 25177 37136 25211
rect 37170 25208 37182 25211
rect 37274 25208 37280 25220
rect 37170 25180 37280 25208
rect 37170 25177 37182 25180
rect 37124 25171 37182 25177
rect 37274 25168 37280 25180
rect 37332 25168 37338 25220
rect 39224 25152 39252 25248
rect 40313 25245 40325 25248
rect 40359 25245 40371 25279
rect 40313 25239 40371 25245
rect 40405 25279 40463 25285
rect 40405 25245 40417 25279
rect 40451 25245 40463 25279
rect 40405 25239 40463 25245
rect 40420 25208 40448 25239
rect 40494 25236 40500 25288
rect 40552 25276 40558 25288
rect 40681 25279 40739 25285
rect 40552 25248 40597 25276
rect 40552 25236 40558 25248
rect 40681 25245 40693 25279
rect 40727 25276 40739 25279
rect 40954 25276 40960 25288
rect 40727 25248 40960 25276
rect 40727 25245 40739 25248
rect 40681 25239 40739 25245
rect 40954 25236 40960 25248
rect 41012 25236 41018 25288
rect 58158 25276 58164 25288
rect 58119 25248 58164 25276
rect 58158 25236 58164 25248
rect 58216 25236 58222 25288
rect 40586 25208 40592 25220
rect 40420 25180 40592 25208
rect 40586 25168 40592 25180
rect 40644 25168 40650 25220
rect 30929 25143 30987 25149
rect 30929 25109 30941 25143
rect 30975 25109 30987 25143
rect 35986 25140 35992 25152
rect 35947 25112 35992 25140
rect 30929 25103 30987 25109
rect 35986 25100 35992 25112
rect 36044 25100 36050 25152
rect 39206 25140 39212 25152
rect 39167 25112 39212 25140
rect 39206 25100 39212 25112
rect 39264 25100 39270 25152
rect 40862 25100 40868 25152
rect 40920 25140 40926 25152
rect 41141 25143 41199 25149
rect 41141 25140 41153 25143
rect 40920 25112 41153 25140
rect 40920 25100 40926 25112
rect 41141 25109 41153 25112
rect 41187 25109 41199 25143
rect 41141 25103 41199 25109
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 4706 24936 4712 24948
rect 4667 24908 4712 24936
rect 4706 24896 4712 24908
rect 4764 24896 4770 24948
rect 7834 24896 7840 24948
rect 7892 24936 7898 24948
rect 10410 24936 10416 24948
rect 7892 24908 10416 24936
rect 7892 24896 7898 24908
rect 10410 24896 10416 24908
rect 10468 24896 10474 24948
rect 10778 24896 10784 24948
rect 10836 24936 10842 24948
rect 10965 24939 11023 24945
rect 10965 24936 10977 24939
rect 10836 24908 10977 24936
rect 10836 24896 10842 24908
rect 10965 24905 10977 24908
rect 11011 24936 11023 24939
rect 11330 24936 11336 24948
rect 11011 24908 11336 24936
rect 11011 24905 11023 24908
rect 10965 24899 11023 24905
rect 11330 24896 11336 24908
rect 11388 24896 11394 24948
rect 12618 24936 12624 24948
rect 12579 24908 12624 24936
rect 12618 24896 12624 24908
rect 12676 24896 12682 24948
rect 14550 24936 14556 24948
rect 12728 24908 14556 24936
rect 10870 24868 10876 24880
rect 3528 24840 3832 24868
rect 2406 24760 2412 24812
rect 2464 24800 2470 24812
rect 3528 24800 3556 24840
rect 2464 24772 3556 24800
rect 2464 24760 2470 24772
rect 3602 24760 3608 24812
rect 3660 24809 3666 24812
rect 3660 24800 3672 24809
rect 3804 24800 3832 24840
rect 10428 24840 10876 24868
rect 3660 24772 3705 24800
rect 3804 24772 3924 24800
rect 3660 24763 3672 24772
rect 3660 24760 3666 24763
rect 3896 24744 3924 24772
rect 4062 24760 4068 24812
rect 4120 24800 4126 24812
rect 5261 24803 5319 24809
rect 5261 24800 5273 24803
rect 4120 24772 5273 24800
rect 4120 24760 4126 24772
rect 5261 24769 5273 24772
rect 5307 24769 5319 24803
rect 10045 24803 10103 24809
rect 10045 24800 10057 24803
rect 5261 24763 5319 24769
rect 9232 24772 10057 24800
rect 3878 24732 3884 24744
rect 3839 24704 3884 24732
rect 3878 24692 3884 24704
rect 3936 24692 3942 24744
rect 5258 24624 5264 24676
rect 5316 24664 5322 24676
rect 9232 24673 9260 24772
rect 10045 24769 10057 24772
rect 10091 24769 10103 24803
rect 10045 24763 10103 24769
rect 10137 24803 10195 24809
rect 10137 24769 10149 24803
rect 10183 24769 10195 24803
rect 10137 24763 10195 24769
rect 10152 24732 10180 24763
rect 10226 24760 10232 24812
rect 10284 24800 10290 24812
rect 10428 24809 10456 24840
rect 10870 24828 10876 24840
rect 10928 24868 10934 24880
rect 12728 24868 12756 24908
rect 14550 24896 14556 24908
rect 14608 24896 14614 24948
rect 15102 24936 15108 24948
rect 14657 24908 15108 24936
rect 14657 24868 14685 24908
rect 15102 24896 15108 24908
rect 15160 24896 15166 24948
rect 15194 24896 15200 24948
rect 15252 24936 15258 24948
rect 15749 24939 15807 24945
rect 15749 24936 15761 24939
rect 15252 24908 15761 24936
rect 15252 24896 15258 24908
rect 15749 24905 15761 24908
rect 15795 24905 15807 24939
rect 24026 24936 24032 24948
rect 15749 24899 15807 24905
rect 15856 24908 24032 24936
rect 10928 24840 12756 24868
rect 13004 24840 14685 24868
rect 10928 24828 10934 24840
rect 10413 24803 10471 24809
rect 10284 24772 10329 24800
rect 10284 24760 10290 24772
rect 10413 24769 10425 24803
rect 10459 24769 10471 24803
rect 10413 24763 10471 24769
rect 11609 24803 11667 24809
rect 11609 24769 11621 24803
rect 11655 24800 11667 24803
rect 11698 24800 11704 24812
rect 11655 24772 11704 24800
rect 11655 24769 11667 24772
rect 11609 24763 11667 24769
rect 11698 24760 11704 24772
rect 11756 24800 11762 24812
rect 12710 24800 12716 24812
rect 11756 24772 12716 24800
rect 11756 24760 11762 24772
rect 12710 24760 12716 24772
rect 12768 24760 12774 24812
rect 12802 24760 12808 24812
rect 12860 24809 12866 24812
rect 13004 24809 13032 24840
rect 14918 24828 14924 24880
rect 14976 24868 14982 24880
rect 15856 24868 15884 24908
rect 24026 24896 24032 24908
rect 24084 24896 24090 24948
rect 27522 24896 27528 24948
rect 27580 24936 27586 24948
rect 30466 24936 30472 24948
rect 27580 24908 30472 24936
rect 27580 24896 27586 24908
rect 30466 24896 30472 24908
rect 30524 24896 30530 24948
rect 18322 24868 18328 24880
rect 14976 24840 15884 24868
rect 17867 24840 18328 24868
rect 14976 24828 14982 24840
rect 12860 24803 12909 24809
rect 12860 24769 12863 24803
rect 12897 24769 12909 24803
rect 12860 24763 12909 24769
rect 12989 24803 13047 24809
rect 12989 24769 13001 24803
rect 13035 24769 13047 24803
rect 12989 24763 13047 24769
rect 12860 24760 12866 24763
rect 11422 24732 11428 24744
rect 10152 24704 11428 24732
rect 11422 24692 11428 24704
rect 11480 24732 11486 24744
rect 13004 24732 13032 24763
rect 13078 24760 13084 24812
rect 13136 24800 13142 24812
rect 13265 24803 13323 24809
rect 13136 24772 13178 24800
rect 13136 24760 13142 24772
rect 13265 24769 13277 24803
rect 13311 24800 13323 24803
rect 13446 24800 13452 24812
rect 13311 24772 13452 24800
rect 13311 24769 13323 24772
rect 13265 24763 13323 24769
rect 13446 24760 13452 24772
rect 13504 24760 13510 24812
rect 14274 24760 14280 24812
rect 14332 24800 14338 24812
rect 14625 24803 14683 24809
rect 14625 24800 14637 24803
rect 14332 24772 14637 24800
rect 14332 24760 14338 24772
rect 14625 24769 14637 24772
rect 14671 24769 14683 24803
rect 14625 24763 14683 24769
rect 16758 24760 16764 24812
rect 16816 24800 16822 24812
rect 16945 24803 17003 24809
rect 16945 24800 16957 24803
rect 16816 24772 16957 24800
rect 16816 24760 16822 24772
rect 16945 24769 16957 24772
rect 16991 24769 17003 24803
rect 16945 24763 17003 24769
rect 17402 24760 17408 24812
rect 17460 24800 17466 24812
rect 17867 24809 17895 24840
rect 18322 24828 18328 24840
rect 18380 24828 18386 24880
rect 21269 24871 21327 24877
rect 21269 24837 21281 24871
rect 21315 24868 21327 24871
rect 21450 24868 21456 24880
rect 21315 24840 21456 24868
rect 21315 24837 21327 24840
rect 21269 24831 21327 24837
rect 21450 24828 21456 24840
rect 21508 24828 21514 24880
rect 23566 24868 23572 24880
rect 22480 24840 23572 24868
rect 17589 24803 17647 24809
rect 17589 24800 17601 24803
rect 17460 24772 17601 24800
rect 17460 24760 17466 24772
rect 17589 24769 17601 24772
rect 17635 24769 17647 24803
rect 17752 24803 17810 24809
rect 17752 24800 17764 24803
rect 17589 24763 17647 24769
rect 17696 24772 17764 24800
rect 11480 24704 13032 24732
rect 14369 24735 14427 24741
rect 11480 24692 11486 24704
rect 14369 24701 14381 24735
rect 14415 24701 14427 24735
rect 14369 24695 14427 24701
rect 9217 24667 9275 24673
rect 9217 24664 9229 24667
rect 5316 24636 9229 24664
rect 5316 24624 5322 24636
rect 9217 24633 9229 24636
rect 9263 24633 9275 24667
rect 12342 24664 12348 24676
rect 9217 24627 9275 24633
rect 12084 24636 12348 24664
rect 2501 24599 2559 24605
rect 2501 24565 2513 24599
rect 2547 24596 2559 24599
rect 2958 24596 2964 24608
rect 2547 24568 2964 24596
rect 2547 24565 2559 24568
rect 2501 24559 2559 24565
rect 2958 24556 2964 24568
rect 3016 24556 3022 24608
rect 7190 24556 7196 24608
rect 7248 24596 7254 24608
rect 7285 24599 7343 24605
rect 7285 24596 7297 24599
rect 7248 24568 7297 24596
rect 7248 24556 7254 24568
rect 7285 24565 7297 24568
rect 7331 24565 7343 24599
rect 9766 24596 9772 24608
rect 9727 24568 9772 24596
rect 7285 24559 7343 24565
rect 9766 24556 9772 24568
rect 9824 24556 9830 24608
rect 11974 24556 11980 24608
rect 12032 24596 12038 24608
rect 12084 24605 12112 24636
rect 12342 24624 12348 24636
rect 12400 24664 12406 24676
rect 12802 24664 12808 24676
rect 12400 24636 12808 24664
rect 12400 24624 12406 24636
rect 12802 24624 12808 24636
rect 12860 24624 12866 24676
rect 12069 24599 12127 24605
rect 12069 24596 12081 24599
rect 12032 24568 12081 24596
rect 12032 24556 12038 24568
rect 12069 24565 12081 24568
rect 12115 24565 12127 24599
rect 12069 24559 12127 24565
rect 12158 24556 12164 24608
rect 12216 24596 12222 24608
rect 13814 24596 13820 24608
rect 12216 24568 13820 24596
rect 12216 24556 12222 24568
rect 13814 24556 13820 24568
rect 13872 24556 13878 24608
rect 14384 24596 14412 24695
rect 17696 24676 17724 24772
rect 17752 24769 17764 24772
rect 17798 24769 17810 24803
rect 17752 24763 17810 24769
rect 17865 24803 17923 24809
rect 17865 24769 17877 24803
rect 17911 24769 17923 24803
rect 17865 24763 17923 24769
rect 18003 24803 18061 24809
rect 18003 24769 18015 24803
rect 18049 24800 18061 24803
rect 18506 24800 18512 24812
rect 18049 24772 18512 24800
rect 18049 24769 18061 24772
rect 18003 24763 18061 24769
rect 18506 24760 18512 24772
rect 18564 24760 18570 24812
rect 18690 24800 18696 24812
rect 18651 24772 18696 24800
rect 18690 24760 18696 24772
rect 18748 24760 18754 24812
rect 21818 24809 21824 24812
rect 18949 24803 19007 24809
rect 18949 24800 18961 24803
rect 18800 24772 18961 24800
rect 18233 24735 18291 24741
rect 18233 24701 18245 24735
rect 18279 24732 18291 24735
rect 18800 24732 18828 24772
rect 18949 24769 18961 24772
rect 18995 24769 19007 24803
rect 18949 24763 19007 24769
rect 21809 24803 21824 24809
rect 21809 24769 21821 24803
rect 21809 24763 21824 24769
rect 21818 24760 21824 24763
rect 21876 24760 21882 24812
rect 22002 24809 22008 24812
rect 22000 24800 22008 24809
rect 21963 24772 22008 24800
rect 22000 24763 22008 24772
rect 22002 24760 22008 24763
rect 22060 24760 22066 24812
rect 22097 24803 22155 24809
rect 22097 24769 22109 24803
rect 22143 24769 22155 24803
rect 22097 24763 22155 24769
rect 22209 24803 22267 24809
rect 22209 24769 22221 24803
rect 22255 24800 22267 24803
rect 22480 24800 22508 24840
rect 23566 24828 23572 24840
rect 23624 24828 23630 24880
rect 28166 24828 28172 24880
rect 28224 24868 28230 24880
rect 28629 24871 28687 24877
rect 28629 24868 28641 24871
rect 28224 24840 28641 24868
rect 28224 24828 28230 24840
rect 28629 24837 28641 24840
rect 28675 24837 28687 24871
rect 28629 24831 28687 24837
rect 31018 24828 31024 24880
rect 31076 24868 31082 24880
rect 32950 24868 32956 24880
rect 31076 24840 32956 24868
rect 31076 24828 31082 24840
rect 32950 24828 32956 24840
rect 33008 24828 33014 24880
rect 38286 24868 38292 24880
rect 38247 24840 38292 24868
rect 38286 24828 38292 24840
rect 38344 24828 38350 24880
rect 22255 24772 22508 24800
rect 22255 24769 22267 24772
rect 22209 24763 22267 24769
rect 18279 24704 18828 24732
rect 18279 24701 18291 24704
rect 18233 24695 18291 24701
rect 22112 24676 22140 24763
rect 22830 24760 22836 24812
rect 22888 24800 22894 24812
rect 22925 24803 22983 24809
rect 22925 24800 22937 24803
rect 22888 24772 22937 24800
rect 22888 24760 22894 24772
rect 22925 24769 22937 24772
rect 22971 24769 22983 24803
rect 22925 24763 22983 24769
rect 23014 24760 23020 24812
rect 23072 24800 23078 24812
rect 23198 24800 23204 24812
rect 23072 24772 23117 24800
rect 23159 24772 23204 24800
rect 23072 24760 23078 24772
rect 23198 24760 23204 24772
rect 23256 24760 23262 24812
rect 23293 24803 23351 24809
rect 23293 24769 23305 24803
rect 23339 24769 23351 24803
rect 23293 24763 23351 24769
rect 23308 24732 23336 24763
rect 23382 24760 23388 24812
rect 23440 24809 23446 24812
rect 23440 24800 23448 24809
rect 23440 24772 23485 24800
rect 23440 24763 23448 24772
rect 23440 24760 23446 24763
rect 28258 24760 28264 24812
rect 28316 24800 28322 24812
rect 28445 24803 28503 24809
rect 28445 24800 28457 24803
rect 28316 24772 28457 24800
rect 28316 24760 28322 24772
rect 28445 24769 28457 24772
rect 28491 24769 28503 24803
rect 28445 24763 28503 24769
rect 29454 24760 29460 24812
rect 29512 24800 29518 24812
rect 30386 24803 30444 24809
rect 30386 24800 30398 24803
rect 29512 24772 30398 24800
rect 29512 24760 29518 24772
rect 30386 24769 30398 24772
rect 30432 24769 30444 24803
rect 30386 24763 30444 24769
rect 30653 24803 30711 24809
rect 30653 24769 30665 24803
rect 30699 24800 30711 24803
rect 30926 24800 30932 24812
rect 30699 24772 30932 24800
rect 30699 24769 30711 24772
rect 30653 24763 30711 24769
rect 30926 24760 30932 24772
rect 30984 24760 30990 24812
rect 28902 24732 28908 24744
rect 23308 24704 28908 24732
rect 28902 24692 28908 24704
rect 28960 24732 28966 24744
rect 28960 24704 29316 24732
rect 28960 24692 28966 24704
rect 16761 24667 16819 24673
rect 16761 24633 16773 24667
rect 16807 24664 16819 24667
rect 17126 24664 17132 24676
rect 16807 24636 17132 24664
rect 16807 24633 16819 24636
rect 16761 24627 16819 24633
rect 17126 24624 17132 24636
rect 17184 24624 17190 24676
rect 17678 24624 17684 24676
rect 17736 24624 17742 24676
rect 22094 24624 22100 24676
rect 22152 24624 22158 24676
rect 25593 24667 25651 24673
rect 25593 24664 25605 24667
rect 22296 24636 25605 24664
rect 15470 24596 15476 24608
rect 14384 24568 15476 24596
rect 15470 24556 15476 24568
rect 15528 24556 15534 24608
rect 20073 24599 20131 24605
rect 20073 24565 20085 24599
rect 20119 24596 20131 24599
rect 20898 24596 20904 24608
rect 20119 24568 20904 24596
rect 20119 24565 20131 24568
rect 20073 24559 20131 24565
rect 20898 24556 20904 24568
rect 20956 24556 20962 24608
rect 20990 24556 20996 24608
rect 21048 24596 21054 24608
rect 22296 24596 22324 24636
rect 25593 24633 25605 24636
rect 25639 24664 25651 24667
rect 26050 24664 26056 24676
rect 25639 24636 26056 24664
rect 25639 24633 25651 24636
rect 25593 24627 25651 24633
rect 26050 24624 26056 24636
rect 26108 24624 26114 24676
rect 28350 24624 28356 24676
rect 28408 24664 28414 24676
rect 29086 24664 29092 24676
rect 28408 24636 29092 24664
rect 28408 24624 28414 24636
rect 29086 24624 29092 24636
rect 29144 24624 29150 24676
rect 29288 24673 29316 24704
rect 29273 24667 29331 24673
rect 29273 24633 29285 24667
rect 29319 24633 29331 24667
rect 29273 24627 29331 24633
rect 21048 24568 22324 24596
rect 22465 24599 22523 24605
rect 21048 24556 21054 24568
rect 22465 24565 22477 24599
rect 22511 24596 22523 24599
rect 23474 24596 23480 24608
rect 22511 24568 23480 24596
rect 22511 24565 22523 24568
rect 22465 24559 22523 24565
rect 23474 24556 23480 24568
rect 23532 24556 23538 24608
rect 23566 24556 23572 24608
rect 23624 24596 23630 24608
rect 26234 24596 26240 24608
rect 23624 24568 23669 24596
rect 26195 24568 26240 24596
rect 23624 24556 23630 24568
rect 26234 24556 26240 24568
rect 26292 24556 26298 24608
rect 28810 24596 28816 24608
rect 28771 24568 28816 24596
rect 28810 24556 28816 24568
rect 28868 24556 28874 24608
rect 37366 24596 37372 24608
rect 37327 24568 37372 24596
rect 37366 24556 37372 24568
rect 37424 24556 37430 24608
rect 38654 24556 38660 24608
rect 38712 24596 38718 24608
rect 39577 24599 39635 24605
rect 39577 24596 39589 24599
rect 38712 24568 39589 24596
rect 38712 24556 38718 24568
rect 39577 24565 39589 24568
rect 39623 24565 39635 24599
rect 39577 24559 39635 24565
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 3878 24352 3884 24404
rect 3936 24392 3942 24404
rect 5445 24395 5503 24401
rect 5445 24392 5457 24395
rect 3936 24364 5457 24392
rect 3936 24352 3942 24364
rect 5445 24361 5457 24364
rect 5491 24361 5503 24395
rect 5445 24355 5503 24361
rect 7834 24352 7840 24404
rect 7892 24392 7898 24404
rect 8021 24395 8079 24401
rect 8021 24392 8033 24395
rect 7892 24364 8033 24392
rect 7892 24352 7898 24364
rect 8021 24361 8033 24364
rect 8067 24392 8079 24395
rect 8067 24364 9904 24392
rect 8067 24361 8079 24364
rect 8021 24355 8079 24361
rect 9876 24324 9904 24364
rect 10134 24352 10140 24404
rect 10192 24392 10198 24404
rect 16574 24392 16580 24404
rect 10192 24364 16580 24392
rect 10192 24352 10198 24364
rect 16574 24352 16580 24364
rect 16632 24352 16638 24404
rect 17678 24352 17684 24404
rect 17736 24392 17742 24404
rect 19245 24395 19303 24401
rect 19245 24392 19257 24395
rect 17736 24364 19257 24392
rect 17736 24352 17742 24364
rect 19245 24361 19257 24364
rect 19291 24361 19303 24395
rect 28166 24392 28172 24404
rect 19245 24355 19303 24361
rect 21192 24364 28172 24392
rect 11330 24324 11336 24336
rect 9876 24296 11336 24324
rect 11330 24284 11336 24296
rect 11388 24284 11394 24336
rect 14274 24324 14280 24336
rect 14235 24296 14280 24324
rect 14274 24284 14280 24296
rect 14332 24284 14338 24336
rect 20162 24324 20168 24336
rect 14476 24296 20168 24324
rect 8202 24216 8208 24268
rect 8260 24256 8266 24268
rect 8941 24259 8999 24265
rect 8941 24256 8953 24259
rect 8260 24228 8953 24256
rect 8260 24216 8266 24228
rect 8941 24225 8953 24228
rect 8987 24225 8999 24259
rect 8941 24219 8999 24225
rect 6914 24188 6920 24200
rect 6875 24160 6920 24188
rect 6914 24148 6920 24160
rect 6972 24148 6978 24200
rect 7190 24188 7196 24200
rect 7103 24160 7196 24188
rect 7190 24148 7196 24160
rect 7248 24148 7254 24200
rect 9208 24191 9266 24197
rect 9208 24157 9220 24191
rect 9254 24188 9266 24191
rect 9766 24188 9772 24200
rect 9254 24160 9772 24188
rect 9254 24157 9266 24160
rect 9208 24151 9266 24157
rect 9766 24148 9772 24160
rect 9824 24148 9830 24200
rect 11287 24191 11345 24197
rect 11287 24188 11299 24191
rect 10796 24160 11299 24188
rect 4154 24120 4160 24132
rect 4115 24092 4160 24120
rect 4154 24080 4160 24092
rect 4212 24080 4218 24132
rect 7208 24120 7236 24148
rect 10796 24132 10824 24160
rect 11287 24157 11299 24160
rect 11333 24157 11345 24191
rect 11422 24188 11428 24200
rect 11383 24160 11428 24188
rect 11287 24151 11345 24157
rect 11422 24148 11428 24160
rect 11480 24148 11486 24200
rect 11517 24191 11575 24197
rect 11517 24157 11529 24191
rect 11563 24157 11575 24191
rect 11517 24151 11575 24157
rect 9858 24120 9864 24132
rect 7208 24092 9864 24120
rect 9858 24080 9864 24092
rect 9916 24080 9922 24132
rect 10778 24120 10784 24132
rect 9968 24092 10784 24120
rect 6546 24012 6552 24064
rect 6604 24052 6610 24064
rect 9968 24052 9996 24092
rect 10778 24080 10784 24092
rect 10836 24080 10842 24132
rect 11532 24120 11560 24151
rect 11698 24148 11704 24200
rect 11756 24188 11762 24200
rect 12161 24191 12219 24197
rect 11756 24160 11801 24188
rect 11756 24148 11762 24160
rect 12161 24157 12173 24191
rect 12207 24188 12219 24191
rect 12894 24188 12900 24200
rect 12207 24160 12900 24188
rect 12207 24157 12219 24160
rect 12161 24151 12219 24157
rect 12894 24148 12900 24160
rect 12952 24148 12958 24200
rect 13814 24148 13820 24200
rect 13872 24188 13878 24200
rect 14476 24188 14504 24296
rect 20162 24284 20168 24296
rect 20220 24284 20226 24336
rect 17773 24259 17831 24265
rect 17773 24225 17785 24259
rect 17819 24256 17831 24259
rect 18322 24256 18328 24268
rect 17819 24228 18328 24256
rect 17819 24225 17831 24228
rect 17773 24219 17831 24225
rect 18322 24216 18328 24228
rect 18380 24216 18386 24268
rect 19444 24228 20944 24256
rect 14533 24191 14591 24197
rect 14533 24188 14545 24191
rect 13872 24160 14545 24188
rect 13872 24148 13878 24160
rect 14533 24157 14545 24160
rect 14579 24157 14591 24191
rect 14533 24151 14591 24157
rect 14626 24191 14684 24197
rect 14626 24157 14638 24191
rect 14672 24157 14684 24191
rect 14626 24151 14684 24157
rect 11790 24120 11796 24132
rect 11532 24092 11796 24120
rect 11790 24080 11796 24092
rect 11848 24080 11854 24132
rect 12428 24123 12486 24129
rect 12428 24089 12440 24123
rect 12474 24120 12486 24123
rect 12618 24120 12624 24132
rect 12474 24092 12624 24120
rect 12474 24089 12486 24092
rect 12428 24083 12486 24089
rect 12618 24080 12624 24092
rect 12676 24080 12682 24132
rect 14640 24120 14668 24151
rect 14734 24148 14740 24200
rect 14792 24185 14798 24200
rect 14792 24157 14834 24185
rect 14792 24148 14798 24157
rect 14918 24148 14924 24200
rect 14976 24188 14982 24200
rect 16666 24188 16672 24200
rect 14976 24160 15021 24188
rect 16627 24160 16672 24188
rect 14976 24148 14982 24160
rect 16666 24148 16672 24160
rect 16724 24148 16730 24200
rect 17494 24188 17500 24200
rect 17455 24160 17500 24188
rect 17494 24148 17500 24160
rect 17552 24148 17558 24200
rect 19444 24197 19472 24228
rect 20916 24200 20944 24228
rect 19429 24191 19487 24197
rect 19429 24157 19441 24191
rect 19475 24157 19487 24191
rect 19429 24151 19487 24157
rect 20809 24191 20867 24197
rect 20809 24157 20821 24191
rect 20855 24157 20867 24191
rect 20809 24151 20867 24157
rect 15102 24120 15108 24132
rect 14640 24092 15108 24120
rect 15102 24080 15108 24092
rect 15160 24080 15166 24132
rect 16209 24123 16267 24129
rect 16209 24089 16221 24123
rect 16255 24120 16267 24123
rect 16758 24120 16764 24132
rect 16255 24092 16764 24120
rect 16255 24089 16267 24092
rect 16209 24083 16267 24089
rect 16758 24080 16764 24092
rect 16816 24080 16822 24132
rect 17218 24080 17224 24132
rect 17276 24120 17282 24132
rect 18230 24120 18236 24132
rect 17276 24092 18236 24120
rect 17276 24080 17282 24092
rect 18230 24080 18236 24092
rect 18288 24080 18294 24132
rect 19150 24080 19156 24132
rect 19208 24120 19214 24132
rect 19613 24123 19671 24129
rect 19613 24120 19625 24123
rect 19208 24092 19625 24120
rect 19208 24080 19214 24092
rect 19613 24089 19625 24092
rect 19659 24089 19671 24123
rect 19613 24083 19671 24089
rect 10318 24052 10324 24064
rect 6604 24024 9996 24052
rect 10279 24024 10324 24052
rect 6604 24012 6610 24024
rect 10318 24012 10324 24024
rect 10376 24012 10382 24064
rect 11054 24052 11060 24064
rect 11015 24024 11060 24052
rect 11054 24012 11060 24024
rect 11112 24012 11118 24064
rect 13538 24052 13544 24064
rect 13451 24024 13544 24052
rect 13538 24012 13544 24024
rect 13596 24052 13602 24064
rect 14550 24052 14556 24064
rect 13596 24024 14556 24052
rect 13596 24012 13602 24024
rect 14550 24012 14556 24024
rect 14608 24012 14614 24064
rect 15286 24012 15292 24064
rect 15344 24052 15350 24064
rect 15565 24055 15623 24061
rect 15565 24052 15577 24055
rect 15344 24024 15577 24052
rect 15344 24012 15350 24024
rect 15565 24021 15577 24024
rect 15611 24021 15623 24055
rect 20824 24052 20852 24151
rect 20898 24148 20904 24200
rect 20956 24188 20962 24200
rect 21192 24197 21220 24364
rect 28166 24352 28172 24364
rect 28224 24352 28230 24404
rect 28353 24395 28411 24401
rect 28353 24361 28365 24395
rect 28399 24392 28411 24395
rect 28994 24392 29000 24404
rect 28399 24364 29000 24392
rect 28399 24361 28411 24364
rect 28353 24355 28411 24361
rect 28994 24352 29000 24364
rect 29052 24352 29058 24404
rect 30745 24395 30803 24401
rect 30745 24361 30757 24395
rect 30791 24392 30803 24395
rect 31754 24392 31760 24404
rect 30791 24364 31760 24392
rect 30791 24361 30803 24364
rect 30745 24355 30803 24361
rect 31754 24352 31760 24364
rect 31812 24352 31818 24404
rect 37274 24392 37280 24404
rect 37235 24364 37280 24392
rect 37274 24352 37280 24364
rect 37332 24352 37338 24404
rect 40862 24392 40868 24404
rect 37844 24364 40868 24392
rect 22738 24284 22744 24336
rect 22796 24324 22802 24336
rect 26234 24324 26240 24336
rect 22796 24296 26240 24324
rect 22796 24284 22802 24296
rect 26234 24284 26240 24296
rect 26292 24324 26298 24336
rect 29270 24324 29276 24336
rect 26292 24296 26464 24324
rect 26292 24284 26298 24296
rect 22186 24216 22192 24268
rect 22244 24256 22250 24268
rect 25866 24256 25872 24268
rect 22244 24228 22452 24256
rect 22244 24216 22250 24228
rect 21177 24191 21235 24197
rect 20956 24160 21001 24188
rect 20956 24148 20962 24160
rect 21177 24157 21189 24191
rect 21223 24157 21235 24191
rect 21177 24151 21235 24157
rect 21315 24191 21373 24197
rect 21315 24157 21327 24191
rect 21361 24188 21373 24191
rect 21634 24188 21640 24200
rect 21361 24160 21640 24188
rect 21361 24157 21373 24160
rect 21315 24151 21373 24157
rect 21634 24148 21640 24160
rect 21692 24188 21698 24200
rect 22424 24197 22452 24228
rect 24964 24228 25872 24256
rect 24964 24200 24992 24228
rect 25866 24216 25872 24228
rect 25924 24256 25930 24268
rect 25924 24228 26188 24256
rect 25924 24216 25930 24228
rect 22053 24191 22111 24197
rect 22053 24188 22065 24191
rect 21692 24160 22065 24188
rect 21692 24148 21698 24160
rect 22053 24157 22065 24160
rect 22099 24157 22111 24191
rect 22053 24151 22111 24157
rect 22409 24191 22467 24197
rect 22409 24157 22421 24191
rect 22455 24157 22467 24191
rect 22409 24151 22467 24157
rect 22557 24191 22615 24197
rect 22557 24157 22569 24191
rect 22603 24188 22615 24191
rect 22646 24188 22652 24200
rect 22603 24160 22652 24188
rect 22603 24157 22615 24160
rect 22557 24151 22615 24157
rect 22646 24148 22652 24160
rect 22704 24148 22710 24200
rect 24486 24148 24492 24200
rect 24544 24188 24550 24200
rect 24673 24191 24731 24197
rect 24673 24188 24685 24191
rect 24544 24160 24685 24188
rect 24544 24148 24550 24160
rect 24673 24157 24685 24160
rect 24719 24157 24731 24191
rect 24836 24191 24894 24197
rect 24836 24188 24848 24191
rect 24673 24151 24731 24157
rect 24780 24160 24848 24188
rect 20990 24080 20996 24132
rect 21048 24120 21054 24132
rect 21085 24123 21143 24129
rect 21085 24120 21097 24123
rect 21048 24092 21097 24120
rect 21048 24080 21054 24092
rect 21085 24089 21097 24092
rect 21131 24089 21143 24123
rect 21542 24120 21548 24132
rect 21085 24083 21143 24089
rect 21376 24092 21548 24120
rect 21376 24052 21404 24092
rect 21542 24080 21548 24092
rect 21600 24080 21606 24132
rect 22189 24123 22247 24129
rect 22189 24089 22201 24123
rect 22235 24089 22247 24123
rect 22189 24083 22247 24089
rect 22281 24123 22339 24129
rect 22281 24089 22293 24123
rect 22327 24120 22339 24123
rect 23198 24120 23204 24132
rect 22327 24092 23204 24120
rect 22327 24089 22339 24092
rect 22281 24083 22339 24089
rect 20824 24024 21404 24052
rect 21453 24055 21511 24061
rect 15565 24015 15623 24021
rect 21453 24021 21465 24055
rect 21499 24052 21511 24055
rect 21818 24052 21824 24064
rect 21499 24024 21824 24052
rect 21499 24021 21511 24024
rect 21453 24015 21511 24021
rect 21818 24012 21824 24024
rect 21876 24012 21882 24064
rect 21910 24012 21916 24064
rect 21968 24052 21974 24064
rect 22204 24052 22232 24083
rect 23198 24080 23204 24092
rect 23256 24080 23262 24132
rect 24578 24080 24584 24132
rect 24636 24120 24642 24132
rect 24780 24120 24808 24160
rect 24836 24157 24848 24160
rect 24882 24157 24894 24191
rect 24836 24151 24894 24157
rect 24946 24148 24952 24200
rect 25004 24188 25010 24200
rect 25087 24191 25145 24197
rect 25004 24160 25049 24188
rect 25004 24148 25010 24160
rect 25087 24157 25099 24191
rect 25133 24188 25145 24191
rect 25406 24188 25412 24200
rect 25133 24160 25412 24188
rect 25133 24157 25145 24160
rect 25087 24151 25145 24157
rect 25406 24148 25412 24160
rect 25464 24148 25470 24200
rect 26050 24188 26056 24200
rect 26011 24160 26056 24188
rect 26050 24148 26056 24160
rect 26108 24148 26114 24200
rect 26160 24197 26188 24228
rect 26145 24191 26203 24197
rect 26145 24157 26157 24191
rect 26191 24157 26203 24191
rect 26145 24151 26203 24157
rect 26234 24148 26240 24200
rect 26292 24188 26298 24200
rect 26436 24197 26464 24296
rect 28644 24296 29276 24324
rect 28644 24197 28672 24296
rect 29270 24284 29276 24296
rect 29328 24324 29334 24336
rect 29328 24296 31754 24324
rect 29328 24284 29334 24296
rect 30006 24256 30012 24268
rect 28736 24228 30012 24256
rect 28736 24197 28764 24228
rect 30006 24216 30012 24228
rect 30064 24256 30070 24268
rect 30064 24228 30420 24256
rect 30064 24216 30070 24228
rect 26421 24191 26479 24197
rect 26292 24160 26337 24188
rect 26292 24148 26298 24160
rect 26421 24157 26433 24191
rect 26467 24157 26479 24191
rect 26421 24151 26479 24157
rect 27893 24191 27951 24197
rect 27893 24157 27905 24191
rect 27939 24188 27951 24191
rect 28629 24191 28687 24197
rect 28629 24188 28641 24191
rect 27939 24160 28641 24188
rect 27939 24157 27951 24160
rect 27893 24151 27951 24157
rect 28629 24157 28641 24160
rect 28675 24157 28687 24191
rect 28629 24151 28687 24157
rect 28721 24191 28779 24197
rect 28721 24157 28733 24191
rect 28767 24157 28779 24191
rect 28721 24151 28779 24157
rect 28350 24120 28356 24132
rect 24636 24092 24808 24120
rect 25148 24092 28356 24120
rect 24636 24080 24642 24092
rect 25148 24052 25176 24092
rect 28350 24080 28356 24092
rect 28408 24080 28414 24132
rect 28442 24080 28448 24132
rect 28500 24120 28506 24132
rect 28736 24120 28764 24151
rect 28810 24148 28816 24200
rect 28868 24188 28874 24200
rect 28997 24191 29055 24197
rect 28868 24160 28913 24188
rect 28868 24148 28874 24160
rect 28997 24157 29009 24191
rect 29043 24188 29055 24191
rect 30098 24188 30104 24200
rect 29043 24160 29132 24188
rect 29043 24157 29055 24160
rect 28997 24151 29055 24157
rect 28500 24092 28764 24120
rect 28500 24080 28506 24092
rect 25314 24052 25320 24064
rect 21968 24024 22013 24052
rect 22204 24024 25176 24052
rect 25275 24024 25320 24052
rect 21968 24012 21974 24024
rect 25314 24012 25320 24024
rect 25372 24012 25378 24064
rect 25777 24055 25835 24061
rect 25777 24021 25789 24055
rect 25823 24052 25835 24055
rect 25866 24052 25872 24064
rect 25823 24024 25872 24052
rect 25823 24021 25835 24024
rect 25777 24015 25835 24021
rect 25866 24012 25872 24024
rect 25924 24012 25930 24064
rect 27249 24055 27307 24061
rect 27249 24021 27261 24055
rect 27295 24052 27307 24055
rect 28810 24052 28816 24064
rect 27295 24024 28816 24052
rect 27295 24021 27307 24024
rect 27249 24015 27307 24021
rect 28810 24012 28816 24024
rect 28868 24052 28874 24064
rect 29104 24052 29132 24160
rect 29564 24160 30104 24188
rect 29564 24061 29592 24160
rect 30098 24148 30104 24160
rect 30156 24148 30162 24200
rect 30282 24188 30288 24200
rect 30243 24160 30288 24188
rect 30282 24148 30288 24160
rect 30340 24148 30346 24200
rect 30392 24197 30420 24228
rect 30377 24191 30435 24197
rect 30377 24157 30389 24191
rect 30423 24157 30435 24191
rect 30377 24151 30435 24157
rect 30469 24191 30527 24197
rect 30469 24157 30481 24191
rect 30515 24157 30527 24191
rect 30469 24151 30527 24157
rect 29549 24055 29607 24061
rect 29549 24052 29561 24055
rect 28868 24024 29561 24052
rect 28868 24012 28874 24024
rect 29549 24021 29561 24024
rect 29595 24021 29607 24055
rect 30484 24052 30512 24151
rect 31726 24120 31754 24296
rect 33594 24284 33600 24336
rect 33652 24324 33658 24336
rect 37844 24324 37872 24364
rect 40862 24352 40868 24364
rect 40920 24352 40926 24404
rect 40954 24324 40960 24336
rect 33652 24296 37872 24324
rect 37936 24296 40960 24324
rect 33652 24284 33658 24296
rect 36449 24259 36507 24265
rect 36449 24225 36461 24259
rect 36495 24256 36507 24259
rect 36495 24228 37780 24256
rect 36495 24225 36507 24228
rect 36449 24219 36507 24225
rect 35986 24148 35992 24200
rect 36044 24188 36050 24200
rect 36633 24191 36691 24197
rect 36633 24188 36645 24191
rect 36044 24160 36645 24188
rect 36044 24148 36050 24160
rect 36633 24157 36645 24160
rect 36679 24157 36691 24191
rect 37366 24188 37372 24200
rect 36633 24151 36691 24157
rect 36740 24160 37372 24188
rect 36740 24120 36768 24160
rect 37366 24148 37372 24160
rect 37424 24188 37430 24200
rect 37752 24197 37780 24228
rect 37936 24197 37964 24296
rect 40954 24284 40960 24296
rect 41012 24284 41018 24336
rect 38746 24216 38752 24268
rect 38804 24256 38810 24268
rect 38804 24228 41368 24256
rect 38804 24216 38810 24228
rect 37553 24191 37611 24197
rect 37553 24188 37565 24191
rect 37424 24160 37565 24188
rect 37424 24148 37430 24160
rect 37553 24157 37565 24160
rect 37599 24157 37611 24191
rect 37553 24151 37611 24157
rect 37645 24191 37703 24197
rect 37645 24157 37657 24191
rect 37691 24157 37703 24191
rect 37645 24151 37703 24157
rect 37737 24191 37795 24197
rect 37737 24157 37749 24191
rect 37783 24157 37795 24191
rect 37737 24151 37795 24157
rect 37921 24191 37979 24197
rect 37921 24157 37933 24191
rect 37967 24157 37979 24191
rect 37921 24151 37979 24157
rect 31726 24092 36768 24120
rect 36817 24123 36875 24129
rect 36817 24089 36829 24123
rect 36863 24089 36875 24123
rect 36817 24083 36875 24089
rect 31297 24055 31355 24061
rect 31297 24052 31309 24055
rect 30484 24024 31309 24052
rect 29549 24015 29607 24021
rect 31297 24021 31309 24024
rect 31343 24052 31355 24055
rect 31570 24052 31576 24064
rect 31343 24024 31576 24052
rect 31343 24021 31355 24024
rect 31297 24015 31355 24021
rect 31570 24012 31576 24024
rect 31628 24012 31634 24064
rect 36832 24052 36860 24083
rect 37550 24052 37556 24064
rect 36832 24024 37556 24052
rect 37550 24012 37556 24024
rect 37608 24012 37614 24064
rect 37660 24052 37688 24151
rect 38562 24148 38568 24200
rect 38620 24188 38626 24200
rect 41340 24197 41368 24228
rect 40497 24191 40555 24197
rect 40497 24188 40509 24191
rect 38620 24160 40509 24188
rect 38620 24148 38626 24160
rect 40497 24157 40509 24160
rect 40543 24157 40555 24191
rect 40497 24151 40555 24157
rect 41325 24191 41383 24197
rect 41325 24157 41337 24191
rect 41371 24157 41383 24191
rect 58158 24188 58164 24200
rect 58119 24160 58164 24188
rect 41325 24151 41383 24157
rect 58158 24148 58164 24160
rect 58216 24148 58222 24200
rect 39574 24080 39580 24132
rect 39632 24120 39638 24132
rect 39850 24120 39856 24132
rect 39632 24092 39856 24120
rect 39632 24080 39638 24092
rect 39850 24080 39856 24092
rect 39908 24120 39914 24132
rect 40313 24123 40371 24129
rect 40313 24120 40325 24123
rect 39908 24092 40325 24120
rect 39908 24080 39914 24092
rect 40313 24089 40325 24092
rect 40359 24120 40371 24123
rect 41141 24123 41199 24129
rect 41141 24120 41153 24123
rect 40359 24092 41153 24120
rect 40359 24089 40371 24092
rect 40313 24083 40371 24089
rect 41141 24089 41153 24092
rect 41187 24089 41199 24123
rect 41141 24083 41199 24089
rect 40586 24052 40592 24064
rect 37660 24024 40592 24052
rect 40586 24012 40592 24024
rect 40644 24012 40650 24064
rect 40681 24055 40739 24061
rect 40681 24021 40693 24055
rect 40727 24052 40739 24055
rect 41046 24052 41052 24064
rect 40727 24024 41052 24052
rect 40727 24021 40739 24024
rect 40681 24015 40739 24021
rect 41046 24012 41052 24024
rect 41104 24012 41110 24064
rect 41506 24052 41512 24064
rect 41467 24024 41512 24052
rect 41506 24012 41512 24024
rect 41564 24012 41570 24064
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 4154 23808 4160 23860
rect 4212 23848 4218 23860
rect 6457 23851 6515 23857
rect 6457 23848 6469 23851
rect 4212 23820 6469 23848
rect 4212 23808 4218 23820
rect 6457 23817 6469 23820
rect 6503 23848 6515 23851
rect 9306 23848 9312 23860
rect 6503 23820 9312 23848
rect 6503 23817 6515 23820
rect 6457 23811 6515 23817
rect 9306 23808 9312 23820
rect 9364 23808 9370 23860
rect 9766 23848 9772 23860
rect 9679 23820 9772 23848
rect 9766 23808 9772 23820
rect 9824 23848 9830 23860
rect 10042 23848 10048 23860
rect 9824 23820 10048 23848
rect 9824 23808 9830 23820
rect 10042 23808 10048 23820
rect 10100 23808 10106 23860
rect 13078 23808 13084 23860
rect 13136 23848 13142 23860
rect 13357 23851 13415 23857
rect 13357 23848 13369 23851
rect 13136 23820 13369 23848
rect 13136 23808 13142 23820
rect 13357 23817 13369 23820
rect 13403 23817 13415 23851
rect 13357 23811 13415 23817
rect 13446 23808 13452 23860
rect 13504 23848 13510 23860
rect 14461 23851 14519 23857
rect 14461 23848 14473 23851
rect 13504 23820 14473 23848
rect 13504 23808 13510 23820
rect 14461 23817 14473 23820
rect 14507 23848 14519 23851
rect 14918 23848 14924 23860
rect 14507 23820 14924 23848
rect 14507 23817 14519 23820
rect 14461 23811 14519 23817
rect 14918 23808 14924 23820
rect 14976 23808 14982 23860
rect 15028 23820 16068 23848
rect 8656 23783 8714 23789
rect 8656 23749 8668 23783
rect 8702 23780 8714 23783
rect 10229 23783 10287 23789
rect 10229 23780 10241 23783
rect 8702 23752 10241 23780
rect 8702 23749 8714 23752
rect 8656 23743 8714 23749
rect 10229 23749 10241 23752
rect 10275 23749 10287 23783
rect 10229 23743 10287 23749
rect 11054 23740 11060 23792
rect 11112 23780 11118 23792
rect 12630 23783 12688 23789
rect 12630 23780 12642 23783
rect 11112 23752 12642 23780
rect 11112 23740 11118 23752
rect 12630 23749 12642 23752
rect 12676 23749 12688 23783
rect 12630 23743 12688 23749
rect 13464 23752 14964 23780
rect 1946 23672 1952 23724
rect 2004 23712 2010 23724
rect 2133 23715 2191 23721
rect 2133 23712 2145 23715
rect 2004 23684 2145 23712
rect 2004 23672 2010 23684
rect 2133 23681 2145 23684
rect 2179 23681 2191 23715
rect 2133 23675 2191 23681
rect 2317 23715 2375 23721
rect 2317 23681 2329 23715
rect 2363 23712 2375 23715
rect 3234 23712 3240 23724
rect 2363 23684 3240 23712
rect 2363 23681 2375 23684
rect 2317 23675 2375 23681
rect 2148 23644 2176 23675
rect 3234 23672 3240 23684
rect 3292 23672 3298 23724
rect 7834 23712 7840 23724
rect 7795 23684 7840 23712
rect 7834 23672 7840 23684
rect 7892 23672 7898 23724
rect 8202 23672 8208 23724
rect 8260 23712 8266 23724
rect 8389 23715 8447 23721
rect 8389 23712 8401 23715
rect 8260 23684 8401 23712
rect 8260 23672 8266 23684
rect 8389 23681 8401 23684
rect 8435 23681 8447 23715
rect 10502 23712 10508 23724
rect 10463 23684 10508 23712
rect 8389 23675 8447 23681
rect 10502 23672 10508 23684
rect 10560 23672 10566 23724
rect 10594 23715 10652 23721
rect 10594 23681 10606 23715
rect 10640 23681 10652 23715
rect 10594 23675 10652 23681
rect 3786 23644 3792 23656
rect 2148 23616 3792 23644
rect 3786 23604 3792 23616
rect 3844 23604 3850 23656
rect 6730 23604 6736 23656
rect 6788 23644 6794 23656
rect 7561 23647 7619 23653
rect 7561 23644 7573 23647
rect 6788 23616 7573 23644
rect 6788 23604 6794 23616
rect 7561 23613 7573 23616
rect 7607 23613 7619 23647
rect 10609 23644 10637 23675
rect 10686 23672 10692 23724
rect 10744 23715 10750 23724
rect 10744 23687 10786 23715
rect 10744 23672 10750 23687
rect 10870 23672 10876 23724
rect 10928 23712 10934 23724
rect 10928 23684 10973 23712
rect 10928 23672 10934 23684
rect 11238 23672 11244 23724
rect 11296 23712 11302 23724
rect 13464 23712 13492 23752
rect 11296 23684 13492 23712
rect 11296 23672 11302 23684
rect 13538 23672 13544 23724
rect 13596 23712 13602 23724
rect 13596 23684 13641 23712
rect 13596 23672 13602 23684
rect 13722 23672 13728 23724
rect 13780 23712 13786 23724
rect 14936 23721 14964 23752
rect 14921 23715 14979 23721
rect 13780 23684 13825 23712
rect 13780 23672 13786 23684
rect 14921 23681 14933 23715
rect 14967 23681 14979 23715
rect 15028 23712 15056 23820
rect 15194 23780 15200 23792
rect 15155 23752 15200 23780
rect 15194 23740 15200 23752
rect 15252 23740 15258 23792
rect 16040 23789 16068 23820
rect 18506 23808 18512 23860
rect 18564 23848 18570 23860
rect 18693 23851 18751 23857
rect 18693 23848 18705 23851
rect 18564 23820 18705 23848
rect 18564 23808 18570 23820
rect 18693 23817 18705 23820
rect 18739 23817 18751 23851
rect 23106 23848 23112 23860
rect 18693 23811 18751 23817
rect 22664 23820 23112 23848
rect 16025 23783 16083 23789
rect 16025 23749 16037 23783
rect 16071 23780 16083 23783
rect 22664 23780 22692 23820
rect 23106 23808 23112 23820
rect 23164 23808 23170 23860
rect 24578 23808 24584 23860
rect 24636 23848 24642 23860
rect 26973 23851 27031 23857
rect 26973 23848 26985 23851
rect 24636 23820 26985 23848
rect 24636 23808 24642 23820
rect 26973 23817 26985 23820
rect 27019 23817 27031 23851
rect 29086 23848 29092 23860
rect 26973 23811 27031 23817
rect 27080 23820 29092 23848
rect 16071 23752 22692 23780
rect 22741 23783 22799 23789
rect 16071 23749 16083 23752
rect 16025 23743 16083 23749
rect 22741 23749 22753 23783
rect 22787 23780 22799 23783
rect 23198 23780 23204 23792
rect 22787 23752 23204 23780
rect 22787 23749 22799 23752
rect 22741 23743 22799 23749
rect 15102 23712 15108 23724
rect 15028 23684 15108 23712
rect 14921 23675 14979 23681
rect 15102 23672 15108 23684
rect 15160 23712 15166 23724
rect 15160 23684 15253 23712
rect 15160 23672 15166 23684
rect 15286 23672 15292 23724
rect 15344 23712 15350 23724
rect 18049 23715 18107 23721
rect 15344 23684 15389 23712
rect 15344 23672 15350 23684
rect 18049 23681 18061 23715
rect 18095 23712 18107 23715
rect 18598 23712 18604 23724
rect 18095 23684 18604 23712
rect 18095 23681 18107 23684
rect 18049 23675 18107 23681
rect 18598 23672 18604 23684
rect 18656 23672 18662 23724
rect 22462 23712 22468 23724
rect 22423 23684 22468 23712
rect 22462 23672 22468 23684
rect 22520 23672 22526 23724
rect 22554 23672 22560 23724
rect 22612 23712 22618 23724
rect 22612 23684 22657 23712
rect 22612 23672 22618 23684
rect 11422 23644 11428 23656
rect 10609 23616 11428 23644
rect 7561 23607 7619 23613
rect 11422 23604 11428 23616
rect 11480 23604 11486 23656
rect 12894 23604 12900 23656
rect 12952 23644 12958 23656
rect 15470 23644 15476 23656
rect 12952 23616 15476 23644
rect 12952 23604 12958 23616
rect 15470 23604 15476 23616
rect 15528 23604 15534 23656
rect 15654 23604 15660 23656
rect 15712 23644 15718 23656
rect 20990 23644 20996 23656
rect 15712 23616 20996 23644
rect 15712 23604 15718 23616
rect 20990 23604 20996 23616
rect 21048 23644 21054 23656
rect 22756 23644 22784 23743
rect 23198 23740 23204 23752
rect 23256 23740 23262 23792
rect 24486 23780 24492 23792
rect 24447 23752 24492 23780
rect 24486 23740 24492 23752
rect 24544 23740 24550 23792
rect 25590 23780 25596 23792
rect 25056 23752 25596 23780
rect 22833 23715 22891 23721
rect 22833 23681 22845 23715
rect 22879 23681 22891 23715
rect 22833 23675 22891 23681
rect 22971 23715 23029 23721
rect 22971 23681 22983 23715
rect 23017 23712 23029 23715
rect 23382 23712 23388 23724
rect 23017 23684 23388 23712
rect 23017 23681 23029 23684
rect 22971 23675 23029 23681
rect 21048 23616 22784 23644
rect 22848 23644 22876 23675
rect 23382 23672 23388 23684
rect 23440 23672 23446 23724
rect 25056 23721 25084 23752
rect 25590 23740 25596 23752
rect 25648 23740 25654 23792
rect 27080 23780 27108 23820
rect 29086 23808 29092 23820
rect 29144 23808 29150 23860
rect 29454 23848 29460 23860
rect 29415 23820 29460 23848
rect 29454 23808 29460 23820
rect 29512 23808 29518 23860
rect 38746 23848 38752 23860
rect 36004 23820 38752 23848
rect 26344 23752 27108 23780
rect 27157 23783 27215 23789
rect 25314 23721 25320 23724
rect 25041 23715 25099 23721
rect 25041 23681 25053 23715
rect 25087 23681 25099 23715
rect 25308 23712 25320 23721
rect 25275 23684 25320 23712
rect 25041 23675 25099 23681
rect 25308 23675 25320 23684
rect 25314 23672 25320 23675
rect 25372 23672 25378 23724
rect 22848 23616 25084 23644
rect 21048 23604 21054 23616
rect 17402 23576 17408 23588
rect 13648 23548 17408 23576
rect 13648 23520 13676 23548
rect 17402 23536 17408 23548
rect 17460 23536 17466 23588
rect 18233 23579 18291 23585
rect 18233 23545 18245 23579
rect 18279 23576 18291 23579
rect 19150 23576 19156 23588
rect 18279 23548 19156 23576
rect 18279 23545 18291 23548
rect 18233 23539 18291 23545
rect 19150 23536 19156 23548
rect 19208 23536 19214 23588
rect 21634 23536 21640 23588
rect 21692 23576 21698 23588
rect 23382 23576 23388 23588
rect 21692 23548 23388 23576
rect 21692 23536 21698 23548
rect 23382 23536 23388 23548
rect 23440 23536 23446 23588
rect 2501 23511 2559 23517
rect 2501 23477 2513 23511
rect 2547 23508 2559 23511
rect 2682 23508 2688 23520
rect 2547 23480 2688 23508
rect 2547 23477 2559 23480
rect 2501 23471 2559 23477
rect 2682 23468 2688 23480
rect 2740 23468 2746 23520
rect 11517 23511 11575 23517
rect 11517 23477 11529 23511
rect 11563 23508 11575 23511
rect 11606 23508 11612 23520
rect 11563 23480 11612 23508
rect 11563 23477 11575 23480
rect 11517 23471 11575 23477
rect 11606 23468 11612 23480
rect 11664 23468 11670 23520
rect 13630 23468 13636 23520
rect 13688 23468 13694 23520
rect 15378 23468 15384 23520
rect 15436 23508 15442 23520
rect 15473 23511 15531 23517
rect 15473 23508 15485 23511
rect 15436 23480 15485 23508
rect 15436 23468 15442 23480
rect 15473 23477 15485 23480
rect 15519 23477 15531 23511
rect 15473 23471 15531 23477
rect 22830 23468 22836 23520
rect 22888 23508 22894 23520
rect 23109 23511 23167 23517
rect 23109 23508 23121 23511
rect 22888 23480 23121 23508
rect 22888 23468 22894 23480
rect 23109 23477 23121 23480
rect 23155 23477 23167 23511
rect 25056 23508 25084 23616
rect 26344 23576 26372 23752
rect 27157 23749 27169 23783
rect 27203 23780 27215 23783
rect 27614 23780 27620 23792
rect 27203 23752 27620 23780
rect 27203 23749 27215 23752
rect 27157 23743 27215 23749
rect 25976 23548 26372 23576
rect 26421 23579 26479 23585
rect 25976 23508 26004 23548
rect 26421 23545 26433 23579
rect 26467 23576 26479 23579
rect 27172 23576 27200 23743
rect 27614 23740 27620 23752
rect 27672 23740 27678 23792
rect 28813 23783 28871 23789
rect 28813 23749 28825 23783
rect 28859 23780 28871 23783
rect 28902 23780 28908 23792
rect 28859 23752 28908 23780
rect 28859 23749 28871 23752
rect 28813 23743 28871 23749
rect 28902 23740 28908 23752
rect 28960 23740 28966 23792
rect 36004 23789 36032 23820
rect 38746 23808 38752 23820
rect 38804 23808 38810 23860
rect 40862 23808 40868 23860
rect 40920 23848 40926 23860
rect 41693 23851 41751 23857
rect 41693 23848 41705 23851
rect 40920 23820 41705 23848
rect 40920 23808 40926 23820
rect 41693 23817 41705 23820
rect 41739 23817 41751 23851
rect 41693 23811 41751 23817
rect 28997 23783 29055 23789
rect 28997 23749 29009 23783
rect 29043 23780 29055 23783
rect 35989 23783 36047 23789
rect 29043 23752 29960 23780
rect 29043 23749 29055 23752
rect 28997 23743 29055 23749
rect 27341 23715 27399 23721
rect 27341 23712 27353 23715
rect 26467 23548 27200 23576
rect 27264 23684 27353 23712
rect 26467 23545 26479 23548
rect 26421 23539 26479 23545
rect 25056 23480 26004 23508
rect 23109 23471 23167 23477
rect 26050 23468 26056 23520
rect 26108 23508 26114 23520
rect 27264 23508 27292 23684
rect 27341 23681 27353 23684
rect 27387 23681 27399 23715
rect 27341 23675 27399 23681
rect 28258 23672 28264 23724
rect 28316 23712 28322 23724
rect 29932 23721 29960 23752
rect 35989 23749 36001 23783
rect 36035 23749 36047 23783
rect 35989 23743 36047 23749
rect 38654 23740 38660 23792
rect 38712 23780 38718 23792
rect 39758 23780 39764 23792
rect 38712 23752 39764 23780
rect 38712 23740 38718 23752
rect 39758 23740 39764 23752
rect 39816 23780 39822 23792
rect 39816 23752 40172 23780
rect 39816 23740 39822 23752
rect 28629 23715 28687 23721
rect 28629 23712 28641 23715
rect 28316 23684 28641 23712
rect 28316 23672 28322 23684
rect 28629 23681 28641 23684
rect 28675 23681 28687 23715
rect 29713 23715 29771 23721
rect 29713 23712 29725 23715
rect 28629 23675 28687 23681
rect 29656 23684 29725 23712
rect 29656 23576 29684 23684
rect 29713 23681 29725 23684
rect 29759 23681 29771 23715
rect 29713 23675 29771 23681
rect 29806 23715 29864 23721
rect 29806 23681 29818 23715
rect 29852 23681 29864 23715
rect 29806 23675 29864 23681
rect 29917 23715 29975 23721
rect 29917 23681 29929 23715
rect 29963 23681 29975 23715
rect 29917 23675 29975 23681
rect 29809 23644 29837 23675
rect 30098 23672 30104 23724
rect 30156 23712 30162 23724
rect 35894 23712 35900 23724
rect 30156 23684 30201 23712
rect 35855 23684 35900 23712
rect 30156 23672 30162 23684
rect 35894 23672 35900 23684
rect 35952 23672 35958 23724
rect 36081 23715 36139 23721
rect 36081 23681 36093 23715
rect 36127 23712 36139 23715
rect 36170 23712 36176 23724
rect 36127 23684 36176 23712
rect 36127 23681 36139 23684
rect 36081 23675 36139 23681
rect 36170 23672 36176 23684
rect 36228 23672 36234 23724
rect 36265 23715 36323 23721
rect 36265 23681 36277 23715
rect 36311 23681 36323 23715
rect 36265 23675 36323 23681
rect 30006 23644 30012 23656
rect 29809 23616 30012 23644
rect 30006 23604 30012 23616
rect 30064 23604 30070 23656
rect 36280 23644 36308 23675
rect 36354 23672 36360 23724
rect 36412 23712 36418 23724
rect 37461 23715 37519 23721
rect 37461 23712 37473 23715
rect 36412 23684 37473 23712
rect 36412 23672 36418 23684
rect 37461 23681 37473 23684
rect 37507 23681 37519 23715
rect 37461 23675 37519 23681
rect 37645 23715 37703 23721
rect 37645 23681 37657 23715
rect 37691 23712 37703 23715
rect 39574 23712 39580 23724
rect 37691 23684 39580 23712
rect 37691 23681 37703 23684
rect 37645 23675 37703 23681
rect 39574 23672 39580 23684
rect 39632 23672 39638 23724
rect 40144 23721 40172 23752
rect 39873 23715 39931 23721
rect 39873 23681 39885 23715
rect 39919 23712 39931 23715
rect 40129 23715 40187 23721
rect 39919 23684 40080 23712
rect 39919 23681 39931 23684
rect 39873 23675 39931 23681
rect 38838 23644 38844 23656
rect 36280 23616 38844 23644
rect 38838 23604 38844 23616
rect 38896 23604 38902 23656
rect 40052 23644 40080 23684
rect 40129 23681 40141 23715
rect 40175 23681 40187 23715
rect 40862 23712 40868 23724
rect 40823 23684 40868 23712
rect 40129 23675 40187 23681
rect 40862 23672 40868 23684
rect 40920 23672 40926 23724
rect 40957 23715 41015 23721
rect 40957 23681 40969 23715
rect 41003 23681 41015 23715
rect 40957 23675 41015 23681
rect 40589 23647 40647 23653
rect 40589 23644 40601 23647
rect 40052 23616 40601 23644
rect 40589 23613 40601 23616
rect 40635 23613 40647 23647
rect 40589 23607 40647 23613
rect 40770 23604 40776 23656
rect 40828 23644 40834 23656
rect 40972 23644 41000 23675
rect 41046 23672 41052 23724
rect 41104 23712 41110 23724
rect 41104 23684 41149 23712
rect 41104 23672 41110 23684
rect 41230 23672 41236 23724
rect 41288 23712 41294 23724
rect 41288 23684 41333 23712
rect 41288 23672 41294 23684
rect 40828 23616 41000 23644
rect 40828 23604 40834 23616
rect 30561 23579 30619 23585
rect 29656 23548 30052 23576
rect 30024 23520 30052 23548
rect 30561 23545 30573 23579
rect 30607 23545 30619 23579
rect 30561 23539 30619 23545
rect 26108 23480 27292 23508
rect 26108 23468 26114 23480
rect 30006 23468 30012 23520
rect 30064 23508 30070 23520
rect 30576 23508 30604 23539
rect 31570 23536 31576 23588
rect 31628 23576 31634 23588
rect 37182 23576 37188 23588
rect 31628 23548 37188 23576
rect 31628 23536 31634 23548
rect 37182 23536 37188 23548
rect 37240 23536 37246 23588
rect 37458 23536 37464 23588
rect 37516 23576 37522 23588
rect 38562 23576 38568 23588
rect 37516 23548 38568 23576
rect 37516 23536 37522 23548
rect 38562 23536 38568 23548
rect 38620 23576 38626 23588
rect 38749 23579 38807 23585
rect 38749 23576 38761 23579
rect 38620 23548 38761 23576
rect 38620 23536 38626 23548
rect 38749 23545 38761 23548
rect 38795 23545 38807 23579
rect 38749 23539 38807 23545
rect 30064 23480 30604 23508
rect 30064 23468 30070 23480
rect 33778 23468 33784 23520
rect 33836 23508 33842 23520
rect 35713 23511 35771 23517
rect 35713 23508 35725 23511
rect 33836 23480 35725 23508
rect 33836 23468 33842 23480
rect 35713 23477 35725 23480
rect 35759 23477 35771 23511
rect 35713 23471 35771 23477
rect 37277 23511 37335 23517
rect 37277 23477 37289 23511
rect 37323 23508 37335 23511
rect 37734 23508 37740 23520
rect 37323 23480 37740 23508
rect 37323 23477 37335 23480
rect 37277 23471 37335 23477
rect 37734 23468 37740 23480
rect 37792 23468 37798 23520
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 3881 23307 3939 23313
rect 3881 23304 3893 23307
rect 2746 23276 3893 23304
rect 2746 23236 2774 23276
rect 3881 23273 3893 23276
rect 3927 23304 3939 23307
rect 4062 23304 4068 23316
rect 3927 23276 4068 23304
rect 3927 23273 3939 23276
rect 3881 23267 3939 23273
rect 4062 23264 4068 23276
rect 4120 23264 4126 23316
rect 4522 23264 4528 23316
rect 4580 23304 4586 23316
rect 4798 23304 4804 23316
rect 4580 23276 4804 23304
rect 4580 23264 4586 23276
rect 4798 23264 4804 23276
rect 4856 23304 4862 23316
rect 5074 23304 5080 23316
rect 4856 23276 5080 23304
rect 4856 23264 4862 23276
rect 5074 23264 5080 23276
rect 5132 23264 5138 23316
rect 10226 23304 10232 23316
rect 10187 23276 10232 23304
rect 10226 23264 10232 23276
rect 10284 23264 10290 23316
rect 11790 23264 11796 23316
rect 11848 23304 11854 23316
rect 11885 23307 11943 23313
rect 11885 23304 11897 23307
rect 11848 23276 11897 23304
rect 11848 23264 11854 23276
rect 11885 23273 11897 23276
rect 11931 23273 11943 23307
rect 11885 23267 11943 23273
rect 20438 23264 20444 23316
rect 20496 23304 20502 23316
rect 20990 23304 20996 23316
rect 20496 23276 20996 23304
rect 20496 23264 20502 23276
rect 20990 23264 20996 23276
rect 21048 23264 21054 23316
rect 21358 23264 21364 23316
rect 21416 23304 21422 23316
rect 22649 23307 22707 23313
rect 22649 23304 22661 23307
rect 21416 23276 22661 23304
rect 21416 23264 21422 23276
rect 22649 23273 22661 23276
rect 22695 23273 22707 23307
rect 32214 23304 32220 23316
rect 22649 23267 22707 23273
rect 32048 23276 32220 23304
rect 2608 23208 2774 23236
rect 2608 23109 2636 23208
rect 5534 23196 5540 23248
rect 5592 23196 5598 23248
rect 5718 23196 5724 23248
rect 5776 23236 5782 23248
rect 7834 23236 7840 23248
rect 5776 23208 5856 23236
rect 7747 23208 7840 23236
rect 5776 23196 5782 23208
rect 5552 23168 5580 23196
rect 5552 23140 5672 23168
rect 2593 23103 2651 23109
rect 2593 23069 2605 23103
rect 2639 23069 2651 23103
rect 2593 23063 2651 23069
rect 2685 23103 2743 23109
rect 2685 23069 2697 23103
rect 2731 23069 2743 23103
rect 2685 23063 2743 23069
rect 2700 23032 2728 23063
rect 2774 23060 2780 23112
rect 2832 23100 2838 23112
rect 2832 23072 2877 23100
rect 2832 23060 2838 23072
rect 2958 23060 2964 23112
rect 3016 23100 3022 23112
rect 5644 23109 5672 23140
rect 5353 23103 5411 23109
rect 3016 23072 4936 23100
rect 3016 23060 3022 23072
rect 2608 23004 2728 23032
rect 2608 22976 2636 23004
rect 4908 22976 4936 23072
rect 5353 23069 5365 23103
rect 5399 23069 5411 23103
rect 5353 23063 5411 23069
rect 5537 23103 5595 23109
rect 5537 23069 5549 23103
rect 5583 23069 5595 23103
rect 5537 23063 5595 23069
rect 5629 23103 5687 23109
rect 5629 23069 5641 23103
rect 5675 23069 5687 23103
rect 5629 23063 5687 23069
rect 5721 23103 5779 23109
rect 5721 23069 5733 23103
rect 5767 23100 5779 23103
rect 5828 23100 5856 23208
rect 7834 23196 7840 23208
rect 7892 23236 7898 23248
rect 11238 23236 11244 23248
rect 7892 23208 11244 23236
rect 7892 23196 7898 23208
rect 11238 23196 11244 23208
rect 11296 23196 11302 23248
rect 11330 23196 11336 23248
rect 11388 23236 11394 23248
rect 12250 23236 12256 23248
rect 11388 23208 12256 23236
rect 11388 23196 11394 23208
rect 12250 23196 12256 23208
rect 12308 23196 12314 23248
rect 16666 23196 16672 23248
rect 16724 23236 16730 23248
rect 16724 23208 19334 23236
rect 16724 23196 16730 23208
rect 9306 23128 9312 23180
rect 9364 23168 9370 23180
rect 14461 23171 14519 23177
rect 14461 23168 14473 23171
rect 9364 23140 14473 23168
rect 9364 23128 9370 23140
rect 14461 23137 14473 23140
rect 14507 23168 14519 23171
rect 19306 23168 19334 23208
rect 23753 23171 23811 23177
rect 23753 23168 23765 23171
rect 14507 23140 16804 23168
rect 19306 23140 23765 23168
rect 14507 23137 14519 23140
rect 14461 23131 14519 23137
rect 5767 23072 5856 23100
rect 5767 23069 5779 23072
rect 5721 23063 5779 23069
rect 2314 22964 2320 22976
rect 2275 22936 2320 22964
rect 2314 22924 2320 22936
rect 2372 22924 2378 22976
rect 2590 22924 2596 22976
rect 2648 22924 2654 22976
rect 4890 22924 4896 22976
rect 4948 22964 4954 22976
rect 5368 22964 5396 23063
rect 5552 23032 5580 23063
rect 6086 23060 6092 23112
rect 6144 23100 6150 23112
rect 6457 23103 6515 23109
rect 6457 23100 6469 23103
rect 6144 23072 6469 23100
rect 6144 23060 6150 23072
rect 6457 23069 6469 23072
rect 6503 23069 6515 23103
rect 6457 23063 6515 23069
rect 9214 23060 9220 23112
rect 9272 23100 9278 23112
rect 10045 23103 10103 23109
rect 9272 23072 9996 23100
rect 9272 23060 9278 23072
rect 5902 23032 5908 23044
rect 5552 23004 5908 23032
rect 5902 22992 5908 23004
rect 5960 22992 5966 23044
rect 5997 23035 6055 23041
rect 5997 23001 6009 23035
rect 6043 23032 6055 23035
rect 6702 23035 6760 23041
rect 6702 23032 6714 23035
rect 6043 23004 6714 23032
rect 6043 23001 6055 23004
rect 5997 22995 6055 23001
rect 6702 23001 6714 23004
rect 6748 23001 6760 23035
rect 6702 22995 6760 23001
rect 9861 23035 9919 23041
rect 9861 23001 9873 23035
rect 9907 23001 9919 23035
rect 9968 23032 9996 23072
rect 10045 23069 10057 23103
rect 10091 23100 10103 23103
rect 10318 23100 10324 23112
rect 10091 23072 10324 23100
rect 10091 23069 10103 23072
rect 10045 23063 10103 23069
rect 10318 23060 10324 23072
rect 10376 23060 10382 23112
rect 11238 23100 11244 23112
rect 10428 23072 11244 23100
rect 10428 23032 10456 23072
rect 11238 23060 11244 23072
rect 11296 23060 11302 23112
rect 11422 23100 11428 23112
rect 11383 23072 11428 23100
rect 11422 23060 11428 23072
rect 11480 23060 11486 23112
rect 13722 23100 13728 23112
rect 12406 23072 13728 23100
rect 9968 23004 10456 23032
rect 9861 22995 9919 23001
rect 6914 22964 6920 22976
rect 4948 22936 6920 22964
rect 4948 22924 4954 22936
rect 6914 22924 6920 22936
rect 6972 22924 6978 22976
rect 9876 22964 9904 22995
rect 11606 22992 11612 23044
rect 11664 23032 11670 23044
rect 12069 23035 12127 23041
rect 12069 23032 12081 23035
rect 11664 23004 12081 23032
rect 11664 22992 11670 23004
rect 12069 23001 12081 23004
rect 12115 23001 12127 23035
rect 12069 22995 12127 23001
rect 12253 23035 12311 23041
rect 12253 23001 12265 23035
rect 12299 23032 12311 23035
rect 12406 23032 12434 23072
rect 13722 23060 13728 23072
rect 13780 23060 13786 23112
rect 16776 23109 16804 23140
rect 23753 23137 23765 23140
rect 23799 23168 23811 23171
rect 23799 23140 24900 23168
rect 23799 23137 23811 23140
rect 23753 23131 23811 23137
rect 16761 23103 16819 23109
rect 16761 23069 16773 23103
rect 16807 23069 16819 23103
rect 16761 23063 16819 23069
rect 18509 23103 18567 23109
rect 18509 23069 18521 23103
rect 18555 23100 18567 23103
rect 19334 23100 19340 23112
rect 18555 23072 19340 23100
rect 18555 23069 18567 23072
rect 18509 23063 18567 23069
rect 19334 23060 19340 23072
rect 19392 23060 19398 23112
rect 22741 23103 22799 23109
rect 22741 23069 22753 23103
rect 22787 23069 22799 23103
rect 22741 23063 22799 23069
rect 12299 23004 12434 23032
rect 12299 23001 12311 23004
rect 12253 22995 12311 23001
rect 12268 22964 12296 22995
rect 18598 22992 18604 23044
rect 18656 23032 18662 23044
rect 18693 23035 18751 23041
rect 18693 23032 18705 23035
rect 18656 23004 18705 23032
rect 18656 22992 18662 23004
rect 18693 23001 18705 23004
rect 18739 23001 18751 23035
rect 22756 23032 22784 23063
rect 22830 23060 22836 23112
rect 22888 23100 22894 23112
rect 24872 23109 24900 23140
rect 24857 23103 24915 23109
rect 22888 23072 22933 23100
rect 22888 23060 22894 23072
rect 24857 23069 24869 23103
rect 24903 23069 24915 23103
rect 25590 23100 25596 23112
rect 25551 23072 25596 23100
rect 24857 23063 24915 23069
rect 25590 23060 25596 23072
rect 25648 23060 25654 23112
rect 25866 23109 25872 23112
rect 25860 23100 25872 23109
rect 25827 23072 25872 23100
rect 25860 23063 25872 23072
rect 25866 23060 25872 23063
rect 25924 23060 25930 23112
rect 26970 23060 26976 23112
rect 27028 23100 27034 23112
rect 31757 23103 31815 23109
rect 31757 23100 31769 23103
rect 27028 23072 31769 23100
rect 27028 23060 27034 23072
rect 31757 23069 31769 23072
rect 31803 23069 31815 23103
rect 31757 23063 31815 23069
rect 31941 23103 31999 23109
rect 31941 23069 31953 23103
rect 31987 23100 31999 23103
rect 32048 23100 32076 23276
rect 32214 23264 32220 23276
rect 32272 23304 32278 23316
rect 34238 23304 34244 23316
rect 32272 23276 34244 23304
rect 32272 23264 32278 23276
rect 34238 23264 34244 23276
rect 34296 23264 34302 23316
rect 36173 23307 36231 23313
rect 35452 23276 36124 23304
rect 35452 23236 35480 23276
rect 34164 23208 35480 23236
rect 33042 23168 33048 23180
rect 32140 23140 33048 23168
rect 32140 23109 32168 23140
rect 33042 23128 33048 23140
rect 33100 23128 33106 23180
rect 34164 23177 34192 23208
rect 34149 23171 34207 23177
rect 34149 23137 34161 23171
rect 34195 23137 34207 23171
rect 35894 23168 35900 23180
rect 34149 23131 34207 23137
rect 35360 23140 35900 23168
rect 35360 23112 35388 23140
rect 35894 23128 35900 23140
rect 35952 23128 35958 23180
rect 31987 23072 32076 23100
rect 32125 23103 32183 23109
rect 31987 23069 31999 23072
rect 31941 23063 31999 23069
rect 32125 23069 32137 23103
rect 32171 23069 32183 23103
rect 33410 23100 33416 23112
rect 32125 23063 32183 23069
rect 32232 23072 33416 23100
rect 24486 23032 24492 23044
rect 22756 23004 24492 23032
rect 18693 22995 18751 23001
rect 24486 22992 24492 23004
rect 24544 22992 24550 23044
rect 25041 23035 25099 23041
rect 25041 23001 25053 23035
rect 25087 23032 25099 23035
rect 25314 23032 25320 23044
rect 25087 23004 25320 23032
rect 25087 23001 25099 23004
rect 25041 22995 25099 23001
rect 25314 22992 25320 23004
rect 25372 23032 25378 23044
rect 31846 23032 31852 23044
rect 25372 23004 31852 23032
rect 25372 22992 25378 23004
rect 31846 22992 31852 23004
rect 31904 22992 31910 23044
rect 32033 23035 32091 23041
rect 32033 23001 32045 23035
rect 32079 23032 32091 23035
rect 32232 23032 32260 23072
rect 33410 23060 33416 23072
rect 33468 23060 33474 23112
rect 35342 23100 35348 23112
rect 35255 23072 35348 23100
rect 35342 23060 35348 23072
rect 35400 23060 35406 23112
rect 35618 23060 35624 23112
rect 35676 23060 35682 23112
rect 35713 23103 35771 23109
rect 35713 23069 35725 23103
rect 35759 23100 35771 23103
rect 35986 23100 35992 23112
rect 35759 23072 35992 23100
rect 35759 23069 35771 23072
rect 35713 23063 35771 23069
rect 35986 23060 35992 23072
rect 36044 23060 36050 23112
rect 36096 23100 36124 23276
rect 36173 23273 36185 23307
rect 36219 23304 36231 23307
rect 36354 23304 36360 23316
rect 36219 23276 36360 23304
rect 36219 23273 36231 23276
rect 36173 23267 36231 23273
rect 36354 23264 36360 23276
rect 36412 23264 36418 23316
rect 37182 23264 37188 23316
rect 37240 23304 37246 23316
rect 39206 23304 39212 23316
rect 37240 23276 39212 23304
rect 37240 23264 37246 23276
rect 39206 23264 39212 23276
rect 39264 23264 39270 23316
rect 37553 23103 37611 23109
rect 37553 23100 37565 23103
rect 36096 23072 37565 23100
rect 37553 23069 37565 23072
rect 37599 23100 37611 23103
rect 38654 23100 38660 23112
rect 37599 23072 38660 23100
rect 37599 23069 37611 23072
rect 37553 23063 37611 23069
rect 38654 23060 38660 23072
rect 38712 23060 38718 23112
rect 39224 23100 39252 23264
rect 41506 23168 41512 23180
rect 40788 23140 41512 23168
rect 40788 23109 40816 23140
rect 41506 23128 41512 23140
rect 41564 23128 41570 23180
rect 40589 23103 40647 23109
rect 40589 23100 40601 23103
rect 39224 23072 40601 23100
rect 40589 23069 40601 23072
rect 40635 23069 40647 23103
rect 40589 23063 40647 23069
rect 40681 23103 40739 23109
rect 40681 23069 40693 23103
rect 40727 23069 40739 23103
rect 40681 23063 40739 23069
rect 40773 23103 40831 23109
rect 40773 23069 40785 23103
rect 40819 23069 40831 23103
rect 40773 23063 40831 23069
rect 40957 23103 41015 23109
rect 40957 23069 40969 23103
rect 41003 23100 41015 23103
rect 41230 23100 41236 23112
rect 41003 23072 41236 23100
rect 41003 23069 41015 23072
rect 40957 23063 41015 23069
rect 33226 23032 33232 23044
rect 32079 23004 32260 23032
rect 32324 23004 33232 23032
rect 32079 23001 32091 23004
rect 32033 22995 32091 23001
rect 15470 22964 15476 22976
rect 9876 22936 12296 22964
rect 15383 22936 15476 22964
rect 15470 22924 15476 22936
rect 15528 22964 15534 22976
rect 16666 22964 16672 22976
rect 15528 22936 16672 22964
rect 15528 22924 15534 22936
rect 16666 22924 16672 22936
rect 16724 22924 16730 22976
rect 18046 22924 18052 22976
rect 18104 22964 18110 22976
rect 18325 22967 18383 22973
rect 18325 22964 18337 22967
rect 18104 22936 18337 22964
rect 18104 22924 18110 22936
rect 18325 22933 18337 22936
rect 18371 22933 18383 22967
rect 18325 22927 18383 22933
rect 22465 22967 22523 22973
rect 22465 22933 22477 22967
rect 22511 22964 22523 22967
rect 22922 22964 22928 22976
rect 22511 22936 22928 22964
rect 22511 22933 22523 22936
rect 22465 22927 22523 22933
rect 22922 22924 22928 22936
rect 22980 22924 22986 22976
rect 26970 22964 26976 22976
rect 26931 22936 26976 22964
rect 26970 22924 26976 22936
rect 27028 22924 27034 22976
rect 28166 22924 28172 22976
rect 28224 22964 28230 22976
rect 28810 22964 28816 22976
rect 28224 22936 28816 22964
rect 28224 22924 28230 22936
rect 28810 22924 28816 22936
rect 28868 22964 28874 22976
rect 32324 22973 32352 23004
rect 33226 22992 33232 23004
rect 33284 22992 33290 23044
rect 33318 22992 33324 23044
rect 33376 23032 33382 23044
rect 33882 23035 33940 23041
rect 33882 23032 33894 23035
rect 33376 23004 33894 23032
rect 33376 22992 33382 23004
rect 33882 23001 33894 23004
rect 33928 23001 33940 23035
rect 33882 22995 33940 23001
rect 35437 23035 35495 23041
rect 35437 23001 35449 23035
rect 35483 23001 35495 23035
rect 35437 22995 35495 23001
rect 35529 23035 35587 23041
rect 35529 23001 35541 23035
rect 35575 23032 35587 23035
rect 35636 23032 35664 23060
rect 37274 23032 37280 23044
rect 37332 23041 37338 23044
rect 35575 23004 35664 23032
rect 37244 23004 37280 23032
rect 35575 23001 35587 23004
rect 35529 22995 35587 23001
rect 29549 22967 29607 22973
rect 29549 22964 29561 22967
rect 28868 22936 29561 22964
rect 28868 22924 28874 22936
rect 29549 22933 29561 22936
rect 29595 22933 29607 22967
rect 29549 22927 29607 22933
rect 32309 22967 32367 22973
rect 32309 22933 32321 22967
rect 32355 22933 32367 22967
rect 32766 22964 32772 22976
rect 32727 22936 32772 22964
rect 32309 22927 32367 22933
rect 32766 22924 32772 22936
rect 32824 22924 32830 22976
rect 34514 22924 34520 22976
rect 34572 22964 34578 22976
rect 35161 22967 35219 22973
rect 35161 22964 35173 22967
rect 34572 22936 35173 22964
rect 34572 22924 34578 22936
rect 35161 22933 35173 22936
rect 35207 22933 35219 22967
rect 35452 22964 35480 22995
rect 37274 22992 37280 23004
rect 37332 22995 37344 23041
rect 40696 23032 40724 23063
rect 41230 23060 41236 23072
rect 41288 23060 41294 23112
rect 40696 23004 40816 23032
rect 37332 22992 37338 22995
rect 40788 22976 40816 23004
rect 36354 22964 36360 22976
rect 35452 22936 36360 22964
rect 35161 22927 35219 22933
rect 36354 22924 36360 22936
rect 36412 22924 36418 22976
rect 40034 22924 40040 22976
rect 40092 22964 40098 22976
rect 40313 22967 40371 22973
rect 40313 22964 40325 22967
rect 40092 22936 40325 22964
rect 40092 22924 40098 22936
rect 40313 22933 40325 22936
rect 40359 22933 40371 22967
rect 40313 22927 40371 22933
rect 40770 22924 40776 22976
rect 40828 22924 40834 22976
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 1581 22763 1639 22769
rect 1581 22729 1593 22763
rect 1627 22760 1639 22763
rect 2774 22760 2780 22772
rect 1627 22732 2780 22760
rect 1627 22729 1639 22732
rect 1581 22723 1639 22729
rect 2774 22720 2780 22732
rect 2832 22720 2838 22772
rect 5718 22760 5724 22772
rect 5679 22732 5724 22760
rect 5718 22720 5724 22732
rect 5776 22720 5782 22772
rect 5902 22720 5908 22772
rect 5960 22760 5966 22772
rect 6365 22763 6423 22769
rect 6365 22760 6377 22763
rect 5960 22732 6377 22760
rect 5960 22720 5966 22732
rect 6365 22729 6377 22732
rect 6411 22729 6423 22763
rect 7193 22763 7251 22769
rect 7193 22760 7205 22763
rect 6365 22723 6423 22729
rect 6472 22732 7205 22760
rect 1946 22692 1952 22704
rect 1907 22664 1952 22692
rect 1946 22652 1952 22664
rect 2004 22652 2010 22704
rect 2314 22652 2320 22704
rect 2372 22692 2378 22704
rect 2654 22695 2712 22701
rect 2654 22692 2666 22695
rect 2372 22664 2666 22692
rect 2372 22652 2378 22664
rect 2654 22661 2666 22664
rect 2700 22661 2712 22695
rect 2654 22655 2712 22661
rect 3786 22652 3792 22704
rect 3844 22692 3850 22704
rect 3844 22664 5120 22692
rect 3844 22652 3850 22664
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22624 1823 22627
rect 2406 22624 2412 22636
rect 1811 22596 1900 22624
rect 2367 22596 2412 22624
rect 1811 22593 1823 22596
rect 1765 22587 1823 22593
rect 1872 22420 1900 22596
rect 2406 22584 2412 22596
rect 2464 22584 2470 22636
rect 4522 22624 4528 22636
rect 4483 22596 4528 22624
rect 4522 22584 4528 22596
rect 4580 22584 4586 22636
rect 4617 22627 4675 22633
rect 4617 22593 4629 22627
rect 4663 22593 4675 22627
rect 4617 22587 4675 22593
rect 4632 22556 4660 22587
rect 4706 22584 4712 22636
rect 4764 22624 4770 22636
rect 4764 22596 4809 22624
rect 4764 22584 4770 22596
rect 4890 22584 4896 22636
rect 4948 22624 4954 22636
rect 5092 22624 5120 22664
rect 6472 22624 6500 22732
rect 7193 22729 7205 22732
rect 7239 22729 7251 22763
rect 7193 22723 7251 22729
rect 9858 22720 9864 22772
rect 9916 22760 9922 22772
rect 10137 22763 10195 22769
rect 10137 22760 10149 22763
rect 9916 22732 10149 22760
rect 9916 22720 9922 22732
rect 10137 22729 10149 22732
rect 10183 22760 10195 22763
rect 10502 22760 10508 22772
rect 10183 22732 10508 22760
rect 10183 22729 10195 22732
rect 10137 22723 10195 22729
rect 10502 22720 10508 22732
rect 10560 22720 10566 22772
rect 11238 22720 11244 22772
rect 11296 22760 11302 22772
rect 11609 22763 11667 22769
rect 11609 22760 11621 22763
rect 11296 22732 11621 22760
rect 11296 22720 11302 22732
rect 11609 22729 11621 22732
rect 11655 22760 11667 22763
rect 13814 22760 13820 22772
rect 11655 22732 13820 22760
rect 11655 22729 11667 22732
rect 11609 22723 11667 22729
rect 13814 22720 13820 22732
rect 13872 22720 13878 22772
rect 15102 22720 15108 22772
rect 15160 22760 15166 22772
rect 15289 22763 15347 22769
rect 15289 22760 15301 22763
rect 15160 22732 15301 22760
rect 15160 22720 15166 22732
rect 15289 22729 15301 22732
rect 15335 22729 15347 22763
rect 15289 22723 15347 22729
rect 19334 22720 19340 22772
rect 19392 22760 19398 22772
rect 19613 22763 19671 22769
rect 19613 22760 19625 22763
rect 19392 22732 19625 22760
rect 19392 22720 19398 22732
rect 19613 22729 19625 22732
rect 19659 22760 19671 22763
rect 20438 22760 20444 22772
rect 19659 22732 20444 22760
rect 19659 22729 19671 22732
rect 19613 22723 19671 22729
rect 20438 22720 20444 22732
rect 20496 22720 20502 22772
rect 22278 22760 22284 22772
rect 20548 22732 22284 22760
rect 6549 22695 6607 22701
rect 6549 22661 6561 22695
rect 6595 22692 6607 22695
rect 7834 22692 7840 22704
rect 6595 22664 7840 22692
rect 6595 22661 6607 22664
rect 6549 22655 6607 22661
rect 7834 22652 7840 22664
rect 7892 22652 7898 22704
rect 14550 22692 14556 22704
rect 14511 22664 14556 22692
rect 14550 22652 14556 22664
rect 14608 22652 14614 22704
rect 14645 22695 14703 22701
rect 14645 22661 14657 22695
rect 14691 22692 14703 22695
rect 15120 22692 15148 22720
rect 14691 22664 15148 22692
rect 16761 22695 16819 22701
rect 14691 22661 14703 22664
rect 14645 22655 14703 22661
rect 16761 22661 16773 22695
rect 16807 22692 16819 22695
rect 20548 22692 20576 22732
rect 22278 22720 22284 22732
rect 22336 22720 22342 22772
rect 26234 22720 26240 22772
rect 26292 22760 26298 22772
rect 26329 22763 26387 22769
rect 26329 22760 26341 22763
rect 26292 22732 26341 22760
rect 26292 22720 26298 22732
rect 26329 22729 26341 22732
rect 26375 22729 26387 22763
rect 26329 22723 26387 22729
rect 27614 22720 27620 22772
rect 27672 22760 27678 22772
rect 33318 22760 33324 22772
rect 27672 22732 33180 22760
rect 33279 22732 33324 22760
rect 27672 22720 27678 22732
rect 26145 22695 26203 22701
rect 16807 22664 20576 22692
rect 21192 22664 25544 22692
rect 16807 22661 16819 22664
rect 16761 22655 16819 22661
rect 6733 22627 6791 22633
rect 6733 22624 6745 22627
rect 4948 22596 4993 22624
rect 5092 22596 6745 22624
rect 4948 22584 4954 22596
rect 6733 22593 6745 22596
rect 6779 22593 6791 22627
rect 6733 22587 6791 22593
rect 7377 22627 7435 22633
rect 7377 22593 7389 22627
rect 7423 22624 7435 22627
rect 14461 22627 14519 22633
rect 7423 22596 7972 22624
rect 7423 22593 7435 22596
rect 7377 22587 7435 22593
rect 5534 22556 5540 22568
rect 4632 22528 5540 22556
rect 5534 22516 5540 22528
rect 5592 22556 5598 22568
rect 6638 22556 6644 22568
rect 5592 22528 6644 22556
rect 5592 22516 5598 22528
rect 6638 22516 6644 22528
rect 6696 22516 6702 22568
rect 7944 22497 7972 22596
rect 14461 22593 14473 22627
rect 14507 22593 14519 22627
rect 14826 22624 14832 22636
rect 14787 22596 14832 22624
rect 14461 22587 14519 22593
rect 14476 22556 14504 22587
rect 14826 22584 14832 22596
rect 14884 22584 14890 22636
rect 15286 22624 15292 22636
rect 14936 22596 15292 22624
rect 14936 22556 14964 22596
rect 15286 22584 15292 22596
rect 15344 22624 15350 22636
rect 16776 22624 16804 22655
rect 18506 22633 18512 22636
rect 15344 22596 16804 22624
rect 15344 22584 15350 22596
rect 18500 22587 18512 22633
rect 18564 22624 18570 22636
rect 21192 22633 21220 22664
rect 21177 22627 21235 22633
rect 18564 22596 18600 22624
rect 18506 22584 18512 22587
rect 18564 22584 18570 22596
rect 21177 22593 21189 22627
rect 21223 22593 21235 22627
rect 21177 22587 21235 22593
rect 21269 22627 21327 22633
rect 21269 22593 21281 22627
rect 21315 22593 21327 22627
rect 21818 22624 21824 22636
rect 21779 22596 21824 22624
rect 21269 22587 21327 22593
rect 14476 22528 14964 22556
rect 16666 22516 16672 22568
rect 16724 22556 16730 22568
rect 18233 22559 18291 22565
rect 18233 22556 18245 22559
rect 16724 22528 18245 22556
rect 16724 22516 16730 22528
rect 18233 22525 18245 22528
rect 18279 22525 18291 22559
rect 21284 22556 21312 22587
rect 21818 22584 21824 22596
rect 21876 22584 21882 22636
rect 22002 22624 22008 22636
rect 21963 22596 22008 22624
rect 22002 22584 22008 22596
rect 22060 22584 22066 22636
rect 23566 22624 23572 22636
rect 22848 22596 23572 22624
rect 22848 22556 22876 22596
rect 23566 22584 23572 22596
rect 23624 22584 23630 22636
rect 24121 22627 24179 22633
rect 24121 22593 24133 22627
rect 24167 22624 24179 22627
rect 24946 22624 24952 22636
rect 24167 22596 24952 22624
rect 24167 22593 24179 22596
rect 24121 22587 24179 22593
rect 24946 22584 24952 22596
rect 25004 22584 25010 22636
rect 21284 22528 22876 22556
rect 18233 22519 18291 22525
rect 23106 22516 23112 22568
rect 23164 22556 23170 22568
rect 23845 22559 23903 22565
rect 23845 22556 23857 22559
rect 23164 22528 23857 22556
rect 23164 22516 23170 22528
rect 23845 22525 23857 22528
rect 23891 22525 23903 22559
rect 23845 22519 23903 22525
rect 3789 22491 3847 22497
rect 3789 22457 3801 22491
rect 3835 22488 3847 22491
rect 7929 22491 7987 22497
rect 3835 22460 7328 22488
rect 3835 22457 3847 22460
rect 3789 22451 3847 22457
rect 3804 22420 3832 22451
rect 1872 22392 3832 22420
rect 4249 22423 4307 22429
rect 4249 22389 4261 22423
rect 4295 22420 4307 22423
rect 4614 22420 4620 22432
rect 4295 22392 4620 22420
rect 4295 22389 4307 22392
rect 4249 22383 4307 22389
rect 4614 22380 4620 22392
rect 4672 22380 4678 22432
rect 7300 22420 7328 22460
rect 7929 22457 7941 22491
rect 7975 22488 7987 22491
rect 16114 22488 16120 22500
rect 7975 22460 16120 22488
rect 7975 22457 7987 22460
rect 7929 22451 7987 22457
rect 16114 22448 16120 22460
rect 16172 22448 16178 22500
rect 8386 22420 8392 22432
rect 7300 22392 8392 22420
rect 8386 22380 8392 22392
rect 8444 22380 8450 22432
rect 14274 22420 14280 22432
rect 14235 22392 14280 22420
rect 14274 22380 14280 22392
rect 14332 22380 14338 22432
rect 15746 22380 15752 22432
rect 15804 22420 15810 22432
rect 15841 22423 15899 22429
rect 15841 22420 15853 22423
rect 15804 22392 15853 22420
rect 15804 22380 15810 22392
rect 15841 22389 15853 22392
rect 15887 22389 15899 22423
rect 15841 22383 15899 22389
rect 17402 22380 17408 22432
rect 17460 22420 17466 22432
rect 17681 22423 17739 22429
rect 17681 22420 17693 22423
rect 17460 22392 17693 22420
rect 17460 22380 17466 22392
rect 17681 22389 17693 22392
rect 17727 22389 17739 22423
rect 17681 22383 17739 22389
rect 17770 22380 17776 22432
rect 17828 22420 17834 22432
rect 20901 22423 20959 22429
rect 20901 22420 20913 22423
rect 17828 22392 20913 22420
rect 17828 22380 17834 22392
rect 20901 22389 20913 22392
rect 20947 22389 20959 22423
rect 21082 22420 21088 22432
rect 21043 22392 21088 22420
rect 20901 22383 20959 22389
rect 21082 22380 21088 22392
rect 21140 22380 21146 22432
rect 21726 22380 21732 22432
rect 21784 22420 21790 22432
rect 21821 22423 21879 22429
rect 21821 22420 21833 22423
rect 21784 22392 21833 22420
rect 21784 22380 21790 22392
rect 21821 22389 21833 22392
rect 21867 22389 21879 22423
rect 21821 22383 21879 22389
rect 22189 22423 22247 22429
rect 22189 22389 22201 22423
rect 22235 22420 22247 22423
rect 22462 22420 22468 22432
rect 22235 22392 22468 22420
rect 22235 22389 22247 22392
rect 22189 22383 22247 22389
rect 22462 22380 22468 22392
rect 22520 22380 22526 22432
rect 22554 22380 22560 22432
rect 22612 22420 22618 22432
rect 22649 22423 22707 22429
rect 22649 22420 22661 22423
rect 22612 22392 22661 22420
rect 22612 22380 22618 22392
rect 22649 22389 22661 22392
rect 22695 22389 22707 22423
rect 22649 22383 22707 22389
rect 23293 22423 23351 22429
rect 23293 22389 23305 22423
rect 23339 22420 23351 22423
rect 23382 22420 23388 22432
rect 23339 22392 23388 22420
rect 23339 22389 23351 22392
rect 23293 22383 23351 22389
rect 23382 22380 23388 22392
rect 23440 22380 23446 22432
rect 25516 22420 25544 22664
rect 26145 22661 26157 22695
rect 26191 22692 26203 22695
rect 26970 22692 26976 22704
rect 26191 22664 26976 22692
rect 26191 22661 26203 22664
rect 26145 22655 26203 22661
rect 26970 22652 26976 22664
rect 27028 22652 27034 22704
rect 32582 22652 32588 22704
rect 32640 22692 32646 22704
rect 33152 22692 33180 22732
rect 33318 22720 33324 22732
rect 33376 22720 33382 22772
rect 33502 22720 33508 22772
rect 33560 22760 33566 22772
rect 35713 22763 35771 22769
rect 33560 22732 34836 22760
rect 33560 22720 33566 22732
rect 34808 22701 34836 22732
rect 35713 22729 35725 22763
rect 35759 22729 35771 22763
rect 37274 22760 37280 22772
rect 37235 22732 37280 22760
rect 35713 22723 35771 22729
rect 34793 22695 34851 22701
rect 32640 22664 32996 22692
rect 33152 22664 34376 22692
rect 32640 22652 32646 22664
rect 25958 22624 25964 22636
rect 25919 22596 25964 22624
rect 25958 22584 25964 22596
rect 26016 22584 26022 22636
rect 27982 22633 27988 22636
rect 27976 22587 27988 22633
rect 28040 22624 28046 22636
rect 28040 22596 28076 22624
rect 27982 22584 27988 22587
rect 28040 22584 28046 22596
rect 31846 22584 31852 22636
rect 31904 22624 31910 22636
rect 32490 22624 32496 22636
rect 31904 22596 32496 22624
rect 31904 22584 31910 22596
rect 32490 22584 32496 22596
rect 32548 22624 32554 22636
rect 32677 22627 32735 22633
rect 32677 22624 32689 22627
rect 32548 22596 32689 22624
rect 32548 22584 32554 22596
rect 32677 22593 32689 22596
rect 32723 22593 32735 22627
rect 32858 22624 32864 22636
rect 32819 22596 32864 22624
rect 32677 22587 32735 22593
rect 32858 22584 32864 22596
rect 32916 22584 32922 22636
rect 32968 22633 32996 22664
rect 32953 22627 33011 22633
rect 32953 22593 32965 22627
rect 32999 22593 33011 22627
rect 32953 22587 33011 22593
rect 33045 22627 33103 22633
rect 33045 22593 33057 22627
rect 33091 22593 33103 22627
rect 33045 22587 33103 22593
rect 25590 22516 25596 22568
rect 25648 22556 25654 22568
rect 27709 22559 27767 22565
rect 27709 22556 27721 22559
rect 25648 22528 27721 22556
rect 25648 22516 25654 22528
rect 27709 22525 27721 22528
rect 27755 22525 27767 22559
rect 27709 22519 27767 22525
rect 32122 22516 32128 22568
rect 32180 22556 32186 22568
rect 33060 22556 33088 22587
rect 33134 22584 33140 22636
rect 33192 22624 33198 22636
rect 33965 22627 34023 22633
rect 33965 22624 33977 22627
rect 33192 22596 33977 22624
rect 33192 22584 33198 22596
rect 33965 22593 33977 22596
rect 34011 22593 34023 22627
rect 33965 22587 34023 22593
rect 34054 22584 34060 22636
rect 34112 22624 34118 22636
rect 34238 22633 34244 22636
rect 34195 22627 34244 22633
rect 34112 22596 34157 22624
rect 34112 22584 34118 22596
rect 34195 22593 34207 22627
rect 34241 22593 34244 22627
rect 34195 22587 34244 22593
rect 34238 22584 34244 22587
rect 34296 22584 34302 22636
rect 34348 22633 34376 22664
rect 34793 22661 34805 22695
rect 34839 22661 34851 22695
rect 34793 22655 34851 22661
rect 34333 22627 34391 22633
rect 34333 22593 34345 22627
rect 34379 22593 34391 22627
rect 34333 22587 34391 22593
rect 35069 22627 35127 22633
rect 35069 22593 35081 22627
rect 35115 22624 35127 22627
rect 35728 22624 35756 22723
rect 37274 22720 37280 22732
rect 37332 22720 37338 22772
rect 40770 22760 40776 22772
rect 37660 22732 40776 22760
rect 35989 22695 36047 22701
rect 35989 22661 36001 22695
rect 36035 22692 36047 22695
rect 37458 22692 37464 22704
rect 36035 22664 37464 22692
rect 36035 22661 36047 22664
rect 35989 22655 36047 22661
rect 37458 22652 37464 22664
rect 37516 22652 37522 22704
rect 35894 22624 35900 22636
rect 35115 22596 35756 22624
rect 35855 22596 35900 22624
rect 35115 22593 35127 22596
rect 35069 22587 35127 22593
rect 35894 22584 35900 22596
rect 35952 22584 35958 22636
rect 36081 22627 36139 22633
rect 36081 22593 36093 22627
rect 36127 22624 36139 22627
rect 36170 22624 36176 22636
rect 36127 22596 36176 22624
rect 36127 22593 36139 22596
rect 36081 22587 36139 22593
rect 33594 22556 33600 22568
rect 32180 22528 33600 22556
rect 32180 22516 32186 22528
rect 33594 22516 33600 22528
rect 33652 22516 33658 22568
rect 34606 22516 34612 22568
rect 34664 22556 34670 22568
rect 34885 22559 34943 22565
rect 34885 22556 34897 22559
rect 34664 22528 34897 22556
rect 34664 22516 34670 22528
rect 34885 22525 34897 22528
rect 34931 22525 34943 22559
rect 34885 22519 34943 22525
rect 35618 22516 35624 22568
rect 35676 22556 35682 22568
rect 36096 22556 36124 22587
rect 36170 22584 36176 22596
rect 36228 22584 36234 22636
rect 36262 22584 36268 22636
rect 36320 22624 36326 22636
rect 36320 22596 36365 22624
rect 36320 22584 36326 22596
rect 37366 22584 37372 22636
rect 37424 22624 37430 22636
rect 37660 22633 37688 22732
rect 40770 22720 40776 22732
rect 40828 22720 40834 22772
rect 39758 22652 39764 22704
rect 39816 22692 39822 22704
rect 39816 22664 40172 22692
rect 39816 22652 39822 22664
rect 37553 22627 37611 22633
rect 37553 22624 37565 22627
rect 37424 22596 37565 22624
rect 37424 22584 37430 22596
rect 37553 22593 37565 22596
rect 37599 22593 37611 22627
rect 37553 22587 37611 22593
rect 37645 22627 37703 22633
rect 37645 22593 37657 22627
rect 37691 22593 37703 22627
rect 37645 22587 37703 22593
rect 37734 22584 37740 22636
rect 37792 22624 37798 22636
rect 37921 22627 37979 22633
rect 37792 22596 37837 22624
rect 37792 22584 37798 22596
rect 37921 22593 37933 22627
rect 37967 22593 37979 22627
rect 37921 22587 37979 22593
rect 39873 22627 39931 22633
rect 39873 22593 39885 22627
rect 39919 22624 39931 22627
rect 40034 22624 40040 22636
rect 39919 22596 40040 22624
rect 39919 22593 39931 22596
rect 39873 22587 39931 22593
rect 35676 22528 36124 22556
rect 35676 22516 35682 22528
rect 36630 22516 36636 22568
rect 36688 22556 36694 22568
rect 37936 22556 37964 22587
rect 40034 22584 40040 22596
rect 40092 22584 40098 22636
rect 40144 22633 40172 22664
rect 40129 22627 40187 22633
rect 40129 22593 40141 22627
rect 40175 22593 40187 22627
rect 40129 22587 40187 22593
rect 36688 22528 37964 22556
rect 36688 22516 36694 22528
rect 28644 22460 32260 22488
rect 28644 22420 28672 22460
rect 29086 22420 29092 22432
rect 25516 22392 28672 22420
rect 29047 22392 29092 22420
rect 29086 22380 29092 22392
rect 29144 22380 29150 22432
rect 30006 22380 30012 22432
rect 30064 22420 30070 22432
rect 32122 22420 32128 22432
rect 30064 22392 32128 22420
rect 30064 22380 30070 22392
rect 32122 22380 32128 22392
rect 32180 22380 32186 22432
rect 32232 22420 32260 22460
rect 32674 22448 32680 22500
rect 32732 22488 32738 22500
rect 32858 22488 32864 22500
rect 32732 22460 32864 22488
rect 32732 22448 32738 22460
rect 32858 22448 32864 22460
rect 32916 22448 32922 22500
rect 35253 22491 35311 22497
rect 35253 22488 35265 22491
rect 33428 22460 35265 22488
rect 33428 22420 33456 22460
rect 35253 22457 35265 22460
rect 35299 22457 35311 22491
rect 38746 22488 38752 22500
rect 38707 22460 38752 22488
rect 35253 22451 35311 22457
rect 38746 22448 38752 22460
rect 38804 22448 38810 22500
rect 58158 22488 58164 22500
rect 58119 22460 58164 22488
rect 58158 22448 58164 22460
rect 58216 22448 58222 22500
rect 32232 22392 33456 22420
rect 33502 22380 33508 22432
rect 33560 22420 33566 22432
rect 33781 22423 33839 22429
rect 33781 22420 33793 22423
rect 33560 22392 33793 22420
rect 33560 22380 33566 22392
rect 33781 22389 33793 22392
rect 33827 22389 33839 22423
rect 33781 22383 33839 22389
rect 34422 22380 34428 22432
rect 34480 22420 34486 22432
rect 34793 22423 34851 22429
rect 34793 22420 34805 22423
rect 34480 22392 34805 22420
rect 34480 22380 34486 22392
rect 34793 22389 34805 22392
rect 34839 22389 34851 22423
rect 34793 22383 34851 22389
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 2590 22176 2596 22228
rect 2648 22216 2654 22228
rect 5534 22216 5540 22228
rect 2648 22188 5540 22216
rect 2648 22176 2654 22188
rect 5534 22176 5540 22188
rect 5592 22176 5598 22228
rect 9309 22219 9367 22225
rect 9309 22185 9321 22219
rect 9355 22216 9367 22219
rect 9674 22216 9680 22228
rect 9355 22188 9680 22216
rect 9355 22185 9367 22188
rect 9309 22179 9367 22185
rect 9674 22176 9680 22188
rect 9732 22216 9738 22228
rect 9732 22188 16528 22216
rect 9732 22176 9738 22188
rect 7377 22151 7435 22157
rect 7377 22117 7389 22151
rect 7423 22148 7435 22151
rect 14826 22148 14832 22160
rect 7423 22120 7457 22148
rect 11072 22120 14832 22148
rect 7423 22117 7435 22120
rect 7377 22111 7435 22117
rect 5994 22080 6000 22092
rect 5955 22052 6000 22080
rect 5994 22040 6000 22052
rect 6052 22040 6058 22092
rect 7392 22080 7420 22111
rect 11072 22080 11100 22120
rect 14826 22108 14832 22120
rect 14884 22108 14890 22160
rect 16500 22148 16528 22188
rect 16574 22176 16580 22228
rect 16632 22216 16638 22228
rect 19981 22219 20039 22225
rect 16632 22188 18644 22216
rect 16632 22176 16638 22188
rect 17402 22148 17408 22160
rect 16500 22120 17408 22148
rect 17402 22108 17408 22120
rect 17460 22148 17466 22160
rect 17862 22148 17868 22160
rect 17460 22120 17868 22148
rect 17460 22108 17466 22120
rect 17862 22108 17868 22120
rect 17920 22108 17926 22160
rect 18506 22148 18512 22160
rect 18467 22120 18512 22148
rect 18506 22108 18512 22120
rect 18564 22108 18570 22160
rect 18616 22148 18644 22188
rect 19981 22185 19993 22219
rect 20027 22216 20039 22219
rect 20346 22216 20352 22228
rect 20027 22188 20352 22216
rect 20027 22185 20039 22188
rect 19981 22179 20039 22185
rect 20346 22176 20352 22188
rect 20404 22176 20410 22228
rect 22646 22176 22652 22228
rect 22704 22216 22710 22228
rect 23382 22216 23388 22228
rect 22704 22188 23388 22216
rect 22704 22176 22710 22188
rect 23382 22176 23388 22188
rect 23440 22176 23446 22228
rect 33502 22216 33508 22228
rect 33463 22188 33508 22216
rect 33502 22176 33508 22188
rect 33560 22176 33566 22228
rect 37366 22176 37372 22228
rect 37424 22216 37430 22228
rect 37461 22219 37519 22225
rect 37461 22216 37473 22219
rect 37424 22188 37473 22216
rect 37424 22176 37430 22188
rect 37461 22185 37473 22188
rect 37507 22185 37519 22219
rect 37461 22179 37519 22185
rect 21821 22151 21879 22157
rect 21821 22148 21833 22151
rect 18616 22120 21833 22148
rect 21821 22117 21833 22120
rect 21867 22148 21879 22151
rect 28074 22148 28080 22160
rect 21867 22120 28080 22148
rect 21867 22117 21879 22120
rect 21821 22111 21879 22117
rect 28074 22108 28080 22120
rect 28132 22108 28138 22160
rect 7392 22052 11100 22080
rect 11164 22052 11652 22080
rect 1857 22015 1915 22021
rect 1857 21981 1869 22015
rect 1903 22012 1915 22015
rect 3789 22015 3847 22021
rect 3789 22012 3801 22015
rect 1903 21984 3801 22012
rect 1903 21981 1915 21984
rect 1857 21975 1915 21981
rect 3789 21981 3801 21984
rect 3835 22012 3847 22015
rect 3878 22012 3884 22024
rect 3835 21984 3884 22012
rect 3835 21981 3847 21984
rect 3789 21975 3847 21981
rect 3878 21972 3884 21984
rect 3936 22012 3942 22024
rect 6012 22012 6040 22040
rect 7392 22012 7420 22052
rect 3936 21984 6040 22012
rect 6104 21984 7420 22012
rect 3936 21972 3942 21984
rect 2124 21947 2182 21953
rect 2124 21913 2136 21947
rect 2170 21944 2182 21947
rect 2222 21944 2228 21956
rect 2170 21916 2228 21944
rect 2170 21913 2182 21916
rect 2124 21907 2182 21913
rect 2222 21904 2228 21916
rect 2280 21904 2286 21956
rect 4056 21947 4114 21953
rect 4056 21913 4068 21947
rect 4102 21944 4114 21947
rect 4614 21944 4620 21956
rect 4102 21916 4620 21944
rect 4102 21913 4114 21916
rect 4056 21907 4114 21913
rect 4614 21904 4620 21916
rect 4672 21904 4678 21956
rect 5626 21904 5632 21956
rect 5684 21944 5690 21956
rect 6104 21944 6132 21984
rect 8386 21972 8392 22024
rect 8444 22012 8450 22024
rect 9861 22015 9919 22021
rect 9861 22012 9873 22015
rect 8444 21984 9873 22012
rect 8444 21972 8450 21984
rect 9861 21981 9873 21984
rect 9907 21981 9919 22015
rect 9861 21975 9919 21981
rect 10229 22015 10287 22021
rect 10229 21981 10241 22015
rect 10275 22012 10287 22015
rect 10410 22012 10416 22024
rect 10275 21984 10416 22012
rect 10275 21981 10287 21984
rect 10229 21975 10287 21981
rect 10410 21972 10416 21984
rect 10468 22012 10474 22024
rect 11164 22012 11192 22052
rect 10468 21984 11192 22012
rect 10468 21972 10474 21984
rect 11238 21972 11244 22024
rect 11296 22012 11302 22024
rect 11514 22012 11520 22024
rect 11296 21984 11341 22012
rect 11475 21984 11520 22012
rect 11296 21972 11302 21984
rect 11514 21972 11520 21984
rect 11572 21972 11578 22024
rect 11624 22021 11652 22052
rect 11698 22040 11704 22092
rect 11756 22080 11762 22092
rect 16761 22083 16819 22089
rect 16761 22080 16773 22083
rect 11756 22052 16773 22080
rect 11756 22040 11762 22052
rect 11609 22015 11667 22021
rect 11609 21981 11621 22015
rect 11655 22012 11667 22015
rect 14090 22012 14096 22024
rect 11655 21984 14096 22012
rect 11655 21981 11667 21984
rect 11609 21975 11667 21981
rect 14090 21972 14096 21984
rect 14148 21972 14154 22024
rect 15580 22021 15608 22052
rect 16761 22049 16773 22052
rect 16807 22049 16819 22083
rect 16761 22043 16819 22049
rect 17770 22040 17776 22092
rect 17828 22080 17834 22092
rect 19889 22083 19947 22089
rect 17828 22052 18276 22080
rect 17828 22040 17834 22052
rect 15565 22015 15623 22021
rect 15565 21981 15577 22015
rect 15611 21981 15623 22015
rect 15746 22012 15752 22024
rect 15707 21984 15752 22012
rect 15565 21975 15623 21981
rect 15746 21972 15752 21984
rect 15804 21972 15810 22024
rect 17037 22015 17095 22021
rect 17037 21981 17049 22015
rect 17083 22012 17095 22015
rect 17218 22012 17224 22024
rect 17083 21984 17224 22012
rect 17083 21981 17095 21984
rect 17037 21975 17095 21981
rect 17218 21972 17224 21984
rect 17276 21972 17282 22024
rect 17862 22012 17868 22024
rect 17823 21984 17868 22012
rect 17862 21972 17868 21984
rect 17920 21972 17926 22024
rect 18046 22012 18052 22024
rect 18007 21984 18052 22012
rect 18046 21972 18052 21984
rect 18104 21972 18110 22024
rect 18248 22021 18276 22052
rect 19889 22049 19901 22083
rect 19935 22080 19947 22083
rect 32950 22080 32956 22092
rect 19935 22052 32956 22080
rect 19935 22049 19947 22052
rect 19889 22043 19947 22049
rect 32950 22040 32956 22052
rect 33008 22040 33014 22092
rect 34514 22080 34520 22092
rect 33244 22052 34520 22080
rect 18141 22015 18199 22021
rect 18141 21981 18153 22015
rect 18187 21981 18199 22015
rect 18141 21975 18199 21981
rect 18233 22015 18291 22021
rect 18233 21981 18245 22015
rect 18279 22012 18291 22015
rect 18874 22012 18880 22024
rect 18279 21984 18880 22012
rect 18279 21981 18291 21984
rect 18233 21975 18291 21981
rect 5684 21916 6132 21944
rect 6264 21947 6322 21953
rect 5684 21904 5690 21916
rect 6264 21913 6276 21947
rect 6310 21944 6322 21947
rect 6362 21944 6368 21956
rect 6310 21916 6368 21944
rect 6310 21913 6322 21916
rect 6264 21907 6322 21913
rect 6362 21904 6368 21916
rect 6420 21904 6426 21956
rect 8938 21904 8944 21956
rect 8996 21944 9002 21956
rect 9217 21947 9275 21953
rect 9217 21944 9229 21947
rect 8996 21916 9229 21944
rect 8996 21904 9002 21916
rect 9217 21913 9229 21916
rect 9263 21913 9275 21947
rect 10042 21944 10048 21956
rect 10003 21916 10048 21944
rect 9217 21907 9275 21913
rect 10042 21904 10048 21916
rect 10100 21904 10106 21956
rect 10137 21947 10195 21953
rect 10137 21913 10149 21947
rect 10183 21944 10195 21947
rect 10318 21944 10324 21956
rect 10183 21916 10324 21944
rect 10183 21913 10195 21916
rect 10137 21907 10195 21913
rect 10318 21904 10324 21916
rect 10376 21904 10382 21956
rect 11422 21944 11428 21956
rect 11383 21916 11428 21944
rect 11422 21904 11428 21916
rect 11480 21944 11486 21956
rect 11698 21944 11704 21956
rect 11480 21916 11704 21944
rect 11480 21904 11486 21916
rect 11698 21904 11704 21916
rect 11756 21904 11762 21956
rect 15381 21947 15439 21953
rect 15381 21913 15393 21947
rect 15427 21944 15439 21947
rect 16114 21944 16120 21956
rect 15427 21916 16120 21944
rect 15427 21913 15439 21916
rect 15381 21907 15439 21913
rect 16114 21904 16120 21916
rect 16172 21904 16178 21956
rect 17494 21904 17500 21956
rect 17552 21944 17558 21956
rect 18156 21944 18184 21975
rect 18874 21972 18880 21984
rect 18932 21972 18938 22024
rect 19981 22015 20039 22021
rect 18984 21984 19748 22012
rect 17552 21916 18184 21944
rect 17552 21904 17558 21916
rect 3234 21876 3240 21888
rect 3195 21848 3240 21876
rect 3234 21836 3240 21848
rect 3292 21836 3298 21888
rect 3970 21836 3976 21888
rect 4028 21876 4034 21888
rect 5169 21879 5227 21885
rect 5169 21876 5181 21879
rect 4028 21848 5181 21876
rect 4028 21836 4034 21848
rect 5169 21845 5181 21848
rect 5215 21876 5227 21879
rect 9950 21876 9956 21888
rect 5215 21848 9956 21876
rect 5215 21845 5227 21848
rect 5169 21839 5227 21845
rect 9950 21836 9956 21848
rect 10008 21836 10014 21888
rect 10413 21879 10471 21885
rect 10413 21845 10425 21879
rect 10459 21876 10471 21879
rect 10962 21876 10968 21888
rect 10459 21848 10968 21876
rect 10459 21845 10471 21848
rect 10413 21839 10471 21845
rect 10962 21836 10968 21848
rect 11020 21836 11026 21888
rect 11793 21879 11851 21885
rect 11793 21845 11805 21879
rect 11839 21876 11851 21879
rect 12618 21876 12624 21888
rect 11839 21848 12624 21876
rect 11839 21845 11851 21848
rect 11793 21839 11851 21845
rect 12618 21836 12624 21848
rect 12676 21836 12682 21888
rect 14918 21876 14924 21888
rect 14879 21848 14924 21876
rect 14918 21836 14924 21848
rect 14976 21836 14982 21888
rect 16942 21836 16948 21888
rect 17000 21876 17006 21888
rect 18984 21876 19012 21984
rect 17000 21848 19012 21876
rect 17000 21836 17006 21848
rect 19334 21836 19340 21888
rect 19392 21876 19398 21888
rect 19613 21879 19671 21885
rect 19613 21876 19625 21879
rect 19392 21848 19625 21876
rect 19392 21836 19398 21848
rect 19613 21845 19625 21848
rect 19659 21845 19671 21879
rect 19720 21876 19748 21984
rect 19981 21981 19993 22015
rect 20027 22012 20039 22015
rect 21910 22012 21916 22024
rect 20027 21984 21916 22012
rect 20027 21981 20039 21984
rect 19981 21975 20039 21981
rect 21910 21972 21916 21984
rect 21968 21972 21974 22024
rect 22554 22012 22560 22024
rect 22066 21984 22560 22012
rect 20254 21904 20260 21956
rect 20312 21944 20318 21956
rect 20533 21947 20591 21953
rect 20533 21944 20545 21947
rect 20312 21916 20545 21944
rect 20312 21904 20318 21916
rect 20533 21913 20545 21916
rect 20579 21913 20591 21947
rect 20533 21907 20591 21913
rect 22066 21876 22094 21984
rect 22554 21972 22560 21984
rect 22612 22012 22618 22024
rect 23017 22015 23075 22021
rect 23017 22012 23029 22015
rect 22612 21984 23029 22012
rect 22612 21972 22618 21984
rect 23017 21981 23029 21984
rect 23063 21981 23075 22015
rect 23017 21975 23075 21981
rect 23106 22009 23164 22015
rect 23106 22002 23118 22009
rect 23152 22002 23164 22009
rect 23106 21950 23112 22002
rect 23164 21950 23170 22002
rect 23198 21972 23204 22024
rect 23256 22012 23262 22024
rect 23382 22012 23388 22024
rect 23256 21984 23301 22012
rect 23343 21984 23388 22012
rect 23256 21972 23262 21984
rect 23382 21972 23388 21984
rect 23440 21972 23446 22024
rect 24394 21972 24400 22024
rect 24452 22012 24458 22024
rect 24489 22015 24547 22021
rect 24489 22012 24501 22015
rect 24452 21984 24501 22012
rect 24452 21972 24458 21984
rect 24489 21981 24501 21984
rect 24535 21981 24547 22015
rect 24489 21975 24547 21981
rect 28445 22015 28503 22021
rect 28445 21981 28457 22015
rect 28491 22012 28503 22015
rect 29086 22012 29092 22024
rect 28491 21984 29092 22012
rect 28491 21981 28503 21984
rect 28445 21975 28503 21981
rect 29086 21972 29092 21984
rect 29144 21972 29150 22024
rect 30466 21972 30472 22024
rect 30524 22012 30530 22024
rect 32033 22015 32091 22021
rect 32033 22012 32045 22015
rect 30524 21984 32045 22012
rect 30524 21972 30530 21984
rect 32033 21981 32045 21984
rect 32079 21981 32091 22015
rect 32214 22012 32220 22024
rect 32175 21984 32220 22012
rect 32033 21975 32091 21981
rect 32214 21972 32220 21984
rect 32272 21972 32278 22024
rect 32398 21972 32404 22024
rect 32456 22012 32462 22024
rect 33042 22012 33048 22024
rect 32456 21984 33048 22012
rect 32456 21972 32462 21984
rect 33042 21972 33048 21984
rect 33100 21972 33106 22024
rect 33244 22021 33272 22052
rect 34514 22040 34520 22052
rect 34572 22040 34578 22092
rect 33229 22015 33287 22021
rect 33229 21981 33241 22015
rect 33275 21981 33287 22015
rect 33229 21975 33287 21981
rect 33318 21972 33324 22024
rect 33376 22012 33382 22024
rect 33505 22015 33563 22021
rect 33376 21984 33421 22012
rect 33376 21972 33382 21984
rect 33505 21981 33517 22015
rect 33551 22012 33563 22015
rect 34238 22012 34244 22024
rect 33551 21984 34244 22012
rect 33551 21981 33563 21984
rect 33505 21975 33563 21981
rect 34238 21972 34244 21984
rect 34296 21972 34302 22024
rect 28258 21944 28264 21956
rect 28219 21916 28264 21944
rect 28258 21904 28264 21916
rect 28316 21904 28322 21956
rect 32309 21947 32367 21953
rect 32309 21913 32321 21947
rect 32355 21944 32367 21947
rect 32766 21944 32772 21956
rect 32355 21916 32772 21944
rect 32355 21913 32367 21916
rect 32309 21907 32367 21913
rect 32766 21904 32772 21916
rect 32824 21904 32830 21956
rect 34422 21944 34428 21956
rect 32876 21916 34428 21944
rect 22738 21876 22744 21888
rect 19720 21848 22094 21876
rect 22699 21848 22744 21876
rect 19613 21839 19671 21845
rect 22738 21836 22744 21848
rect 22796 21836 22802 21888
rect 24673 21879 24731 21885
rect 24673 21845 24685 21879
rect 24719 21876 24731 21879
rect 25958 21876 25964 21888
rect 24719 21848 25964 21876
rect 24719 21845 24731 21848
rect 24673 21839 24731 21845
rect 25958 21836 25964 21848
rect 26016 21836 26022 21888
rect 28629 21879 28687 21885
rect 28629 21845 28641 21879
rect 28675 21876 28687 21879
rect 28718 21876 28724 21888
rect 28675 21848 28724 21876
rect 28675 21845 28687 21848
rect 28629 21839 28687 21845
rect 28718 21836 28724 21848
rect 28776 21836 28782 21888
rect 32585 21879 32643 21885
rect 32585 21845 32597 21879
rect 32631 21876 32643 21879
rect 32876 21876 32904 21916
rect 34422 21904 34428 21916
rect 34480 21904 34486 21956
rect 33042 21876 33048 21888
rect 32631 21848 32904 21876
rect 33003 21848 33048 21876
rect 32631 21845 32643 21848
rect 32585 21839 32643 21845
rect 33042 21836 33048 21848
rect 33100 21836 33106 21888
rect 36630 21836 36636 21888
rect 36688 21876 36694 21888
rect 36909 21879 36967 21885
rect 36909 21876 36921 21879
rect 36688 21848 36921 21876
rect 36688 21836 36694 21848
rect 36909 21845 36921 21848
rect 36955 21845 36967 21879
rect 36909 21839 36967 21845
rect 40313 21879 40371 21885
rect 40313 21845 40325 21879
rect 40359 21876 40371 21879
rect 40678 21876 40684 21888
rect 40359 21848 40684 21876
rect 40359 21845 40371 21848
rect 40313 21839 40371 21845
rect 40678 21836 40684 21848
rect 40736 21836 40742 21888
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 2222 21672 2228 21684
rect 2183 21644 2228 21672
rect 2222 21632 2228 21644
rect 2280 21632 2286 21684
rect 2590 21632 2596 21684
rect 2648 21632 2654 21684
rect 4157 21675 4215 21681
rect 4157 21641 4169 21675
rect 4203 21672 4215 21675
rect 4706 21672 4712 21684
rect 4203 21644 4712 21672
rect 4203 21641 4215 21644
rect 4157 21635 4215 21641
rect 4706 21632 4712 21644
rect 4764 21632 4770 21684
rect 6362 21672 6368 21684
rect 6323 21644 6368 21672
rect 6362 21632 6368 21644
rect 6420 21632 6426 21684
rect 6454 21632 6460 21684
rect 6512 21672 6518 21684
rect 6822 21672 6828 21684
rect 6512 21644 6828 21672
rect 6512 21632 6518 21644
rect 6822 21632 6828 21644
rect 6880 21672 6886 21684
rect 7469 21675 7527 21681
rect 7469 21672 7481 21675
rect 6880 21644 7481 21672
rect 6880 21632 6886 21644
rect 7469 21641 7481 21644
rect 7515 21641 7527 21675
rect 7469 21635 7527 21641
rect 10042 21632 10048 21684
rect 10100 21672 10106 21684
rect 11422 21672 11428 21684
rect 10100 21644 11428 21672
rect 10100 21632 10106 21644
rect 11422 21632 11428 21644
rect 11480 21632 11486 21684
rect 12158 21672 12164 21684
rect 12119 21644 12164 21672
rect 12158 21632 12164 21644
rect 12216 21632 12222 21684
rect 17862 21632 17868 21684
rect 17920 21672 17926 21684
rect 21085 21675 21143 21681
rect 21085 21672 21097 21675
rect 17920 21644 21097 21672
rect 17920 21632 17926 21644
rect 21085 21641 21097 21644
rect 21131 21672 21143 21675
rect 22094 21672 22100 21684
rect 21131 21644 22100 21672
rect 21131 21641 21143 21644
rect 21085 21635 21143 21641
rect 22094 21632 22100 21644
rect 22152 21632 22158 21684
rect 23198 21632 23204 21684
rect 23256 21672 23262 21684
rect 23753 21675 23811 21681
rect 23753 21672 23765 21675
rect 23256 21644 23765 21672
rect 23256 21632 23262 21644
rect 23753 21641 23765 21644
rect 23799 21641 23811 21675
rect 23753 21635 23811 21641
rect 27982 21632 27988 21684
rect 28040 21672 28046 21684
rect 28077 21675 28135 21681
rect 28077 21672 28089 21675
rect 28040 21644 28089 21672
rect 28040 21632 28046 21644
rect 28077 21641 28089 21644
rect 28123 21641 28135 21675
rect 28718 21672 28724 21684
rect 28077 21635 28135 21641
rect 28644 21644 28724 21672
rect 2498 21536 2504 21548
rect 2459 21508 2504 21536
rect 2498 21496 2504 21508
rect 2556 21496 2562 21548
rect 2608 21545 2636 21632
rect 3970 21604 3976 21616
rect 3931 21576 3976 21604
rect 3970 21564 3976 21576
rect 4028 21564 4034 21616
rect 5626 21604 5632 21616
rect 5587 21576 5632 21604
rect 5626 21564 5632 21576
rect 5684 21564 5690 21616
rect 5813 21607 5871 21613
rect 5813 21573 5825 21607
rect 5859 21604 5871 21607
rect 5859 21576 6868 21604
rect 5859 21573 5871 21576
rect 5813 21567 5871 21573
rect 2593 21539 2651 21545
rect 2593 21505 2605 21539
rect 2639 21505 2651 21539
rect 2593 21499 2651 21505
rect 2682 21496 2688 21548
rect 2740 21536 2746 21548
rect 2869 21539 2927 21545
rect 2740 21508 2785 21536
rect 2740 21496 2746 21508
rect 2869 21505 2881 21539
rect 2915 21536 2927 21539
rect 2958 21536 2964 21548
rect 2915 21508 2964 21536
rect 2915 21505 2927 21508
rect 2869 21499 2927 21505
rect 2958 21496 2964 21508
rect 3016 21496 3022 21548
rect 3786 21536 3792 21548
rect 3699 21508 3792 21536
rect 3786 21496 3792 21508
rect 3844 21536 3850 21548
rect 5445 21539 5503 21545
rect 5445 21536 5457 21539
rect 3844 21508 5457 21536
rect 3844 21496 3850 21508
rect 5445 21505 5457 21508
rect 5491 21505 5503 21539
rect 5445 21499 5503 21505
rect 6454 21496 6460 21548
rect 6512 21536 6518 21548
rect 6595 21539 6653 21545
rect 6595 21536 6607 21539
rect 6512 21508 6607 21536
rect 6512 21496 6518 21508
rect 6595 21505 6607 21508
rect 6641 21505 6653 21539
rect 6730 21536 6736 21548
rect 6691 21508 6736 21536
rect 6595 21499 6653 21505
rect 6730 21496 6736 21508
rect 6788 21496 6794 21548
rect 6840 21545 6868 21576
rect 9766 21564 9772 21616
rect 9824 21604 9830 21616
rect 10229 21607 10287 21613
rect 10229 21604 10241 21607
rect 9824 21576 10241 21604
rect 9824 21564 9830 21576
rect 10229 21573 10241 21576
rect 10275 21573 10287 21607
rect 10229 21567 10287 21573
rect 15289 21607 15347 21613
rect 15289 21573 15301 21607
rect 15335 21604 15347 21607
rect 18509 21607 18567 21613
rect 18509 21604 18521 21607
rect 15335 21576 18521 21604
rect 15335 21573 15347 21576
rect 15289 21567 15347 21573
rect 18509 21573 18521 21576
rect 18555 21604 18567 21607
rect 18598 21604 18604 21616
rect 18555 21576 18604 21604
rect 18555 21573 18567 21576
rect 18509 21567 18567 21573
rect 6825 21539 6883 21545
rect 6825 21505 6837 21539
rect 6871 21505 6883 21539
rect 7006 21536 7012 21548
rect 6967 21508 7012 21536
rect 6825 21499 6883 21505
rect 7006 21496 7012 21508
rect 7064 21496 7070 21548
rect 9950 21536 9956 21548
rect 9911 21508 9956 21536
rect 9950 21496 9956 21508
rect 10008 21496 10014 21548
rect 10042 21496 10048 21548
rect 10100 21536 10106 21548
rect 10137 21539 10195 21545
rect 10137 21536 10149 21539
rect 10100 21508 10149 21536
rect 10100 21496 10106 21508
rect 10137 21505 10149 21508
rect 10183 21505 10195 21539
rect 10137 21499 10195 21505
rect 10321 21539 10379 21545
rect 10321 21505 10333 21539
rect 10367 21536 10379 21539
rect 10410 21536 10416 21548
rect 10367 21508 10416 21536
rect 10367 21505 10379 21508
rect 10321 21499 10379 21505
rect 10410 21496 10416 21508
rect 10468 21496 10474 21548
rect 12158 21496 12164 21548
rect 12216 21536 12222 21548
rect 12253 21539 12311 21545
rect 12253 21536 12265 21539
rect 12216 21508 12265 21536
rect 12216 21496 12222 21508
rect 12253 21505 12265 21508
rect 12299 21505 12311 21539
rect 12253 21499 12311 21505
rect 14829 21539 14887 21545
rect 14829 21505 14841 21539
rect 14875 21536 14887 21539
rect 15304 21536 15332 21567
rect 18598 21564 18604 21576
rect 18656 21564 18662 21616
rect 23106 21604 23112 21616
rect 22940 21576 23112 21604
rect 15470 21536 15476 21548
rect 14875 21508 15332 21536
rect 15431 21508 15476 21536
rect 14875 21505 14887 21508
rect 14829 21499 14887 21505
rect 15470 21496 15476 21508
rect 15528 21496 15534 21548
rect 16942 21545 16948 21548
rect 16936 21499 16948 21545
rect 17000 21536 17006 21548
rect 18693 21539 18751 21545
rect 17000 21508 17036 21536
rect 16942 21496 16948 21499
rect 17000 21496 17006 21508
rect 18693 21505 18705 21539
rect 18739 21536 18751 21539
rect 20346 21536 20352 21548
rect 18739 21508 20352 21536
rect 18739 21505 18751 21508
rect 18693 21499 18751 21505
rect 3234 21428 3240 21480
rect 3292 21468 3298 21480
rect 11238 21468 11244 21480
rect 3292 21440 11244 21468
rect 3292 21428 3298 21440
rect 11238 21428 11244 21440
rect 11296 21428 11302 21480
rect 14918 21428 14924 21480
rect 14976 21468 14982 21480
rect 15657 21471 15715 21477
rect 15657 21468 15669 21471
rect 14976 21440 15669 21468
rect 14976 21428 14982 21440
rect 15657 21437 15669 21440
rect 15703 21437 15715 21471
rect 16666 21468 16672 21480
rect 16627 21440 16672 21468
rect 15657 21431 15715 21437
rect 16666 21428 16672 21440
rect 16724 21428 16730 21480
rect 18708 21468 18736 21499
rect 20346 21496 20352 21508
rect 20404 21496 20410 21548
rect 21082 21496 21088 21548
rect 21140 21536 21146 21548
rect 21177 21539 21235 21545
rect 21177 21536 21189 21539
rect 21140 21508 21189 21536
rect 21140 21496 21146 21508
rect 21177 21505 21189 21508
rect 21223 21505 21235 21539
rect 22646 21536 22652 21548
rect 22607 21508 22652 21536
rect 21177 21499 21235 21505
rect 22646 21496 22652 21508
rect 22704 21496 22710 21548
rect 22830 21536 22836 21548
rect 22791 21508 22836 21536
rect 22830 21496 22836 21508
rect 22888 21496 22894 21548
rect 22940 21545 22968 21576
rect 23106 21564 23112 21576
rect 23164 21564 23170 21616
rect 23658 21564 23664 21616
rect 23716 21604 23722 21616
rect 24121 21607 24179 21613
rect 24121 21604 24133 21607
rect 23716 21576 24133 21604
rect 23716 21564 23722 21576
rect 24121 21573 24133 21576
rect 24167 21604 24179 21607
rect 24394 21604 24400 21616
rect 24167 21576 24400 21604
rect 24167 21573 24179 21576
rect 24121 21567 24179 21573
rect 24394 21564 24400 21576
rect 24452 21564 24458 21616
rect 24486 21564 24492 21616
rect 24544 21604 24550 21616
rect 24544 21576 27292 21604
rect 24544 21564 24550 21576
rect 22925 21539 22983 21545
rect 22925 21505 22937 21539
rect 22971 21505 22983 21539
rect 22925 21499 22983 21505
rect 23017 21539 23075 21545
rect 23017 21505 23029 21539
rect 23063 21505 23075 21539
rect 23934 21536 23940 21548
rect 23895 21508 23940 21536
rect 23017 21499 23075 21505
rect 18064 21440 18736 21468
rect 10505 21403 10563 21409
rect 10505 21369 10517 21403
rect 10551 21400 10563 21403
rect 11514 21400 11520 21412
rect 10551 21372 11520 21400
rect 10551 21369 10563 21372
rect 10505 21363 10563 21369
rect 11514 21360 11520 21372
rect 11572 21360 11578 21412
rect 18064 21409 18092 21440
rect 18874 21428 18880 21480
rect 18932 21468 18938 21480
rect 22189 21471 22247 21477
rect 22189 21468 22201 21471
rect 18932 21440 22201 21468
rect 18932 21428 18938 21440
rect 22189 21437 22201 21440
rect 22235 21468 22247 21471
rect 23032 21468 23060 21499
rect 23934 21496 23940 21508
rect 23992 21496 23998 21548
rect 26421 21539 26479 21545
rect 26421 21505 26433 21539
rect 26467 21505 26479 21539
rect 26421 21499 26479 21505
rect 23842 21468 23848 21480
rect 22235 21440 23060 21468
rect 23124 21440 23848 21468
rect 22235 21437 22247 21440
rect 22189 21431 22247 21437
rect 18049 21403 18107 21409
rect 14476 21372 15884 21400
rect 14476 21344 14504 21372
rect 8938 21332 8944 21344
rect 8899 21304 8944 21332
rect 8938 21292 8944 21304
rect 8996 21292 9002 21344
rect 10778 21292 10784 21344
rect 10836 21332 10842 21344
rect 14185 21335 14243 21341
rect 14185 21332 14197 21335
rect 10836 21304 14197 21332
rect 10836 21292 10842 21304
rect 14185 21301 14197 21304
rect 14231 21332 14243 21335
rect 14458 21332 14464 21344
rect 14231 21304 14464 21332
rect 14231 21301 14243 21304
rect 14185 21295 14243 21301
rect 14458 21292 14464 21304
rect 14516 21292 14522 21344
rect 14642 21332 14648 21344
rect 14603 21304 14648 21332
rect 14642 21292 14648 21304
rect 14700 21292 14706 21344
rect 15856 21332 15884 21372
rect 18049 21369 18061 21403
rect 18095 21369 18107 21403
rect 18049 21363 18107 21369
rect 18708 21372 19012 21400
rect 18708 21332 18736 21372
rect 18874 21332 18880 21344
rect 15856 21304 18736 21332
rect 18835 21304 18880 21332
rect 18874 21292 18880 21304
rect 18932 21292 18938 21344
rect 18984 21332 19012 21372
rect 19242 21360 19248 21412
rect 19300 21400 19306 21412
rect 20254 21400 20260 21412
rect 19300 21372 20260 21400
rect 19300 21360 19306 21372
rect 20254 21360 20260 21372
rect 20312 21400 20318 21412
rect 20349 21403 20407 21409
rect 20349 21400 20361 21403
rect 20312 21372 20361 21400
rect 20312 21360 20318 21372
rect 20349 21369 20361 21372
rect 20395 21369 20407 21403
rect 20349 21363 20407 21369
rect 19797 21335 19855 21341
rect 19797 21332 19809 21335
rect 18984 21304 19809 21332
rect 19797 21301 19809 21304
rect 19843 21332 19855 21335
rect 21082 21332 21088 21344
rect 19843 21304 21088 21332
rect 19843 21301 19855 21304
rect 19797 21295 19855 21301
rect 21082 21292 21088 21304
rect 21140 21292 21146 21344
rect 21174 21292 21180 21344
rect 21232 21332 21238 21344
rect 23124 21332 23152 21440
rect 23842 21428 23848 21440
rect 23900 21428 23906 21480
rect 23198 21360 23204 21412
rect 23256 21400 23262 21412
rect 23256 21372 25176 21400
rect 23256 21360 23262 21372
rect 23290 21332 23296 21344
rect 21232 21304 23152 21332
rect 23251 21304 23296 21332
rect 21232 21292 21238 21304
rect 23290 21292 23296 21304
rect 23348 21292 23354 21344
rect 25148 21341 25176 21372
rect 25133 21335 25191 21341
rect 25133 21301 25145 21335
rect 25179 21332 25191 21335
rect 25682 21332 25688 21344
rect 25179 21304 25688 21332
rect 25179 21301 25191 21304
rect 25133 21295 25191 21301
rect 25682 21292 25688 21304
rect 25740 21292 25746 21344
rect 25958 21292 25964 21344
rect 26016 21332 26022 21344
rect 26436 21332 26464 21499
rect 27264 21400 27292 21576
rect 27614 21496 27620 21548
rect 27672 21536 27678 21548
rect 28307 21539 28365 21545
rect 28307 21536 28319 21539
rect 27672 21508 28319 21536
rect 27672 21496 27678 21508
rect 28307 21505 28319 21508
rect 28353 21505 28365 21539
rect 28439 21536 28445 21548
rect 28400 21508 28445 21536
rect 28307 21499 28365 21505
rect 28439 21496 28445 21508
rect 28497 21496 28503 21548
rect 28558 21545 28616 21551
rect 28558 21511 28570 21545
rect 28604 21542 28616 21545
rect 28644 21542 28672 21644
rect 28718 21632 28724 21644
rect 28776 21632 28782 21684
rect 32585 21675 32643 21681
rect 32585 21641 32597 21675
rect 32631 21672 32643 21675
rect 32674 21672 32680 21684
rect 32631 21644 32680 21672
rect 32631 21641 32643 21644
rect 32585 21635 32643 21641
rect 32674 21632 32680 21644
rect 32732 21632 32738 21684
rect 32950 21632 32956 21684
rect 33008 21672 33014 21684
rect 33045 21675 33103 21681
rect 33045 21672 33057 21675
rect 33008 21644 33057 21672
rect 33008 21632 33014 21644
rect 33045 21641 33057 21644
rect 33091 21641 33103 21675
rect 34698 21672 34704 21684
rect 33045 21635 33103 21641
rect 33244 21644 34704 21672
rect 30377 21607 30435 21613
rect 30377 21573 30389 21607
rect 30423 21604 30435 21607
rect 32401 21607 32459 21613
rect 30423 21576 32352 21604
rect 30423 21573 30435 21576
rect 30377 21567 30435 21573
rect 28604 21514 28672 21542
rect 28721 21539 28779 21545
rect 28604 21511 28616 21514
rect 28558 21505 28616 21511
rect 28721 21505 28733 21539
rect 28767 21505 28779 21539
rect 28721 21499 28779 21505
rect 30101 21539 30159 21545
rect 30101 21505 30113 21539
rect 30147 21536 30159 21539
rect 30926 21536 30932 21548
rect 30147 21508 30932 21536
rect 30147 21505 30159 21508
rect 30101 21499 30159 21505
rect 27706 21428 27712 21480
rect 27764 21468 27770 21480
rect 28736 21468 28764 21499
rect 30926 21496 30932 21508
rect 30984 21496 30990 21548
rect 32217 21539 32275 21545
rect 32217 21505 32229 21539
rect 32263 21505 32275 21539
rect 32324 21536 32352 21576
rect 32401 21573 32413 21607
rect 32447 21604 32459 21607
rect 32766 21604 32772 21616
rect 32447 21576 32772 21604
rect 32447 21573 32459 21576
rect 32401 21567 32459 21573
rect 32766 21564 32772 21576
rect 32824 21564 32830 21616
rect 33244 21604 33272 21644
rect 34698 21632 34704 21644
rect 34756 21632 34762 21684
rect 32876 21576 33272 21604
rect 33505 21607 33563 21613
rect 32876 21536 32904 21576
rect 33505 21573 33517 21607
rect 33551 21604 33563 21607
rect 34330 21604 34336 21616
rect 33551 21576 34336 21604
rect 33551 21573 33563 21576
rect 33505 21567 33563 21573
rect 34330 21564 34336 21576
rect 34388 21564 34394 21616
rect 39700 21607 39758 21613
rect 39700 21573 39712 21607
rect 39746 21604 39758 21607
rect 40405 21607 40463 21613
rect 40405 21604 40417 21607
rect 39746 21576 40417 21604
rect 39746 21573 39758 21576
rect 39700 21567 39758 21573
rect 40405 21573 40417 21576
rect 40451 21573 40463 21607
rect 40405 21567 40463 21573
rect 32324 21508 32904 21536
rect 33229 21539 33287 21545
rect 32217 21499 32275 21505
rect 33229 21505 33241 21539
rect 33275 21536 33287 21539
rect 33778 21536 33784 21548
rect 33275 21508 33784 21536
rect 33275 21505 33287 21508
rect 33229 21499 33287 21505
rect 29181 21471 29239 21477
rect 29181 21468 29193 21471
rect 27764 21440 29193 21468
rect 27764 21428 27770 21440
rect 29181 21437 29193 21440
rect 29227 21437 29239 21471
rect 30282 21468 30288 21480
rect 30243 21440 30288 21468
rect 29181 21431 29239 21437
rect 30282 21428 30288 21440
rect 30340 21428 30346 21480
rect 32232 21468 32260 21499
rect 33778 21496 33784 21508
rect 33836 21496 33842 21548
rect 39390 21496 39396 21548
rect 39448 21536 39454 21548
rect 40678 21536 40684 21548
rect 39448 21508 39988 21536
rect 40639 21508 40684 21536
rect 39448 21496 39454 21508
rect 32766 21468 32772 21480
rect 32232 21440 32772 21468
rect 32766 21428 32772 21440
rect 32824 21428 32830 21480
rect 33413 21471 33471 21477
rect 33413 21437 33425 21471
rect 33459 21468 33471 21471
rect 33686 21468 33692 21480
rect 33459 21440 33692 21468
rect 33459 21437 33471 21440
rect 33413 21431 33471 21437
rect 33686 21428 33692 21440
rect 33744 21428 33750 21480
rect 39960 21477 39988 21508
rect 40678 21496 40684 21508
rect 40736 21496 40742 21548
rect 40773 21539 40831 21545
rect 40773 21505 40785 21539
rect 40819 21505 40831 21539
rect 40773 21499 40831 21505
rect 39945 21471 40003 21477
rect 39945 21437 39957 21471
rect 39991 21437 40003 21471
rect 39945 21431 40003 21437
rect 40586 21428 40592 21480
rect 40644 21468 40650 21480
rect 40788 21468 40816 21499
rect 40862 21496 40868 21548
rect 40920 21536 40926 21548
rect 41049 21539 41107 21545
rect 40920 21508 40965 21536
rect 40920 21496 40926 21508
rect 41049 21505 41061 21539
rect 41095 21505 41107 21539
rect 41049 21499 41107 21505
rect 40644 21440 40816 21468
rect 40644 21428 40650 21440
rect 29917 21403 29975 21409
rect 29917 21400 29929 21403
rect 27264 21372 29929 21400
rect 29917 21369 29929 21372
rect 29963 21369 29975 21403
rect 29917 21363 29975 21369
rect 40494 21360 40500 21412
rect 40552 21400 40558 21412
rect 40954 21400 40960 21412
rect 40552 21372 40960 21400
rect 40552 21360 40558 21372
rect 40954 21360 40960 21372
rect 41012 21400 41018 21412
rect 41064 21400 41092 21499
rect 41012 21372 41092 21400
rect 41012 21360 41018 21372
rect 26973 21335 27031 21341
rect 26973 21332 26985 21335
rect 26016 21304 26985 21332
rect 26016 21292 26022 21304
rect 26973 21301 26985 21304
rect 27019 21301 27031 21335
rect 27614 21332 27620 21344
rect 27575 21304 27620 21332
rect 26973 21295 27031 21301
rect 27614 21292 27620 21304
rect 27672 21292 27678 21344
rect 30098 21332 30104 21344
rect 30059 21304 30104 21332
rect 30098 21292 30104 21304
rect 30156 21292 30162 21344
rect 33226 21332 33232 21344
rect 33187 21304 33232 21332
rect 33226 21292 33232 21304
rect 33284 21292 33290 21344
rect 38562 21332 38568 21344
rect 38523 21304 38568 21332
rect 38562 21292 38568 21304
rect 38620 21292 38626 21344
rect 58158 21332 58164 21344
rect 58119 21304 58164 21332
rect 58158 21292 58164 21304
rect 58216 21292 58222 21344
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 10870 21128 10876 21140
rect 10831 21100 10876 21128
rect 10870 21088 10876 21100
rect 10928 21088 10934 21140
rect 13170 21088 13176 21140
rect 13228 21128 13234 21140
rect 13630 21128 13636 21140
rect 13228 21100 13636 21128
rect 13228 21088 13234 21100
rect 13630 21088 13636 21100
rect 13688 21128 13694 21140
rect 14645 21131 14703 21137
rect 14645 21128 14657 21131
rect 13688 21100 14657 21128
rect 13688 21088 13694 21100
rect 14645 21097 14657 21100
rect 14691 21097 14703 21131
rect 14645 21091 14703 21097
rect 16577 21131 16635 21137
rect 16577 21097 16589 21131
rect 16623 21128 16635 21131
rect 16850 21128 16856 21140
rect 16623 21100 16856 21128
rect 16623 21097 16635 21100
rect 16577 21091 16635 21097
rect 16850 21088 16856 21100
rect 16908 21088 16914 21140
rect 16942 21088 16948 21140
rect 17000 21128 17006 21140
rect 17037 21131 17095 21137
rect 17037 21128 17049 21131
rect 17000 21100 17049 21128
rect 17000 21088 17006 21100
rect 17037 21097 17049 21100
rect 17083 21097 17095 21131
rect 17037 21091 17095 21097
rect 22002 21088 22008 21140
rect 22060 21128 22066 21140
rect 30098 21128 30104 21140
rect 22060 21100 26924 21128
rect 30059 21100 30104 21128
rect 22060 21088 22066 21100
rect 11609 21063 11667 21069
rect 11609 21029 11621 21063
rect 11655 21060 11667 21063
rect 13262 21060 13268 21072
rect 11655 21032 13268 21060
rect 11655 21029 11667 21032
rect 11609 21023 11667 21029
rect 13262 21020 13268 21032
rect 13320 21020 13326 21072
rect 13722 21020 13728 21072
rect 13780 21060 13786 21072
rect 16025 21063 16083 21069
rect 16025 21060 16037 21063
rect 13780 21032 16037 21060
rect 13780 21020 13786 21032
rect 16025 21029 16037 21032
rect 16071 21029 16083 21063
rect 21361 21063 21419 21069
rect 21361 21060 21373 21063
rect 16025 21023 16083 21029
rect 17236 21032 21373 21060
rect 13630 20952 13636 21004
rect 13688 20992 13694 21004
rect 13688 20964 15516 20992
rect 13688 20952 13694 20964
rect 10229 20927 10287 20933
rect 10229 20893 10241 20927
rect 10275 20924 10287 20927
rect 10778 20924 10784 20936
rect 10275 20896 10784 20924
rect 10275 20893 10287 20896
rect 10229 20887 10287 20893
rect 10778 20884 10784 20896
rect 10836 20884 10842 20936
rect 11422 20924 11428 20936
rect 11383 20896 11428 20924
rect 11422 20884 11428 20896
rect 11480 20884 11486 20936
rect 12805 20927 12863 20933
rect 12805 20893 12817 20927
rect 12851 20924 12863 20927
rect 14642 20924 14648 20936
rect 12851 20896 14648 20924
rect 12851 20893 12863 20896
rect 12805 20887 12863 20893
rect 12342 20816 12348 20868
rect 12400 20856 12406 20868
rect 12820 20856 12848 20887
rect 14642 20884 14648 20896
rect 14700 20884 14706 20936
rect 15378 20924 15384 20936
rect 15339 20896 15384 20924
rect 15378 20884 15384 20896
rect 15436 20884 15442 20936
rect 15488 20933 15516 20964
rect 15474 20927 15532 20933
rect 15474 20893 15486 20927
rect 15520 20893 15532 20927
rect 15474 20887 15532 20893
rect 15654 20884 15660 20936
rect 15712 20924 15718 20936
rect 15887 20927 15945 20933
rect 15712 20896 15757 20924
rect 15712 20884 15718 20896
rect 15887 20893 15899 20927
rect 15933 20924 15945 20927
rect 17236 20924 17264 21032
rect 21361 21029 21373 21032
rect 21407 21060 21419 21063
rect 21634 21060 21640 21072
rect 21407 21032 21640 21060
rect 21407 21029 21419 21032
rect 21361 21023 21419 21029
rect 21634 21020 21640 21032
rect 21692 21020 21698 21072
rect 26896 21060 26924 21100
rect 30098 21088 30104 21100
rect 30156 21088 30162 21140
rect 30926 21088 30932 21140
rect 30984 21128 30990 21140
rect 36541 21131 36599 21137
rect 36541 21128 36553 21131
rect 30984 21100 36553 21128
rect 30984 21088 30990 21100
rect 36541 21097 36553 21100
rect 36587 21097 36599 21131
rect 38562 21128 38568 21140
rect 36541 21091 36599 21097
rect 37108 21100 38568 21128
rect 33042 21060 33048 21072
rect 26896 21032 33048 21060
rect 33042 21020 33048 21032
rect 33100 21020 33106 21072
rect 18874 20992 18880 21004
rect 17512 20964 18880 20992
rect 17512 20933 17540 20964
rect 18874 20952 18880 20964
rect 18932 20952 18938 21004
rect 20364 20964 21220 20992
rect 15933 20896 17264 20924
rect 17293 20927 17351 20933
rect 17497 20927 17555 20933
rect 15933 20893 15945 20896
rect 15887 20887 15945 20893
rect 17293 20893 17305 20927
rect 17339 20924 17351 20927
rect 17339 20893 17356 20924
rect 17293 20887 17356 20893
rect 12400 20828 12848 20856
rect 12989 20859 13047 20865
rect 12400 20816 12406 20828
rect 12989 20825 13001 20859
rect 13035 20856 13047 20859
rect 13630 20856 13636 20868
rect 13035 20828 13636 20856
rect 13035 20825 13047 20828
rect 12989 20819 13047 20825
rect 13630 20816 13636 20828
rect 13688 20816 13694 20868
rect 14458 20816 14464 20868
rect 14516 20856 14522 20868
rect 14553 20859 14611 20865
rect 14553 20856 14565 20859
rect 14516 20828 14565 20856
rect 14516 20816 14522 20828
rect 14553 20825 14565 20828
rect 14599 20825 14611 20859
rect 15746 20856 15752 20868
rect 15707 20828 15752 20856
rect 14553 20819 14611 20825
rect 15746 20816 15752 20828
rect 15804 20816 15810 20868
rect 16850 20816 16856 20868
rect 16908 20856 16914 20868
rect 17328 20856 17356 20887
rect 17386 20921 17444 20927
rect 17386 20887 17398 20921
rect 17432 20918 17444 20921
rect 17432 20887 17448 20918
rect 17497 20893 17509 20927
rect 17543 20893 17555 20927
rect 17497 20887 17555 20893
rect 17681 20927 17739 20933
rect 17681 20893 17693 20927
rect 17727 20924 17739 20927
rect 17862 20924 17868 20936
rect 17727 20896 17868 20924
rect 17727 20893 17739 20896
rect 17681 20887 17739 20893
rect 17386 20881 17448 20887
rect 17862 20884 17868 20896
rect 17920 20884 17926 20936
rect 19978 20884 19984 20936
rect 20036 20924 20042 20936
rect 20119 20927 20177 20933
rect 20119 20924 20131 20927
rect 20036 20896 20131 20924
rect 20036 20884 20042 20896
rect 20119 20893 20131 20896
rect 20165 20924 20177 20927
rect 20364 20924 20392 20964
rect 20165 20896 20392 20924
rect 20165 20893 20177 20896
rect 20119 20887 20177 20893
rect 20438 20884 20444 20936
rect 20496 20933 20502 20936
rect 20496 20927 20535 20933
rect 20523 20893 20535 20927
rect 20496 20887 20535 20893
rect 20496 20884 20502 20887
rect 20622 20884 20628 20936
rect 20680 20924 20686 20936
rect 21192 20933 21220 20964
rect 24578 20952 24584 21004
rect 24636 20992 24642 21004
rect 26694 20992 26700 21004
rect 24636 20964 26700 20992
rect 24636 20952 24642 20964
rect 26694 20952 26700 20964
rect 26752 20952 26758 21004
rect 27062 20952 27068 21004
rect 27120 20992 27126 21004
rect 30834 20992 30840 21004
rect 27120 20964 30840 20992
rect 27120 20952 27126 20964
rect 30834 20952 30840 20964
rect 30892 20952 30898 21004
rect 21177 20927 21235 20933
rect 20680 20896 20725 20924
rect 20680 20884 20686 20896
rect 21177 20893 21189 20927
rect 21223 20893 21235 20927
rect 21177 20887 21235 20893
rect 22465 20927 22523 20933
rect 22465 20893 22477 20927
rect 22511 20924 22523 20927
rect 23198 20924 23204 20936
rect 22511 20896 23204 20924
rect 22511 20893 22523 20896
rect 22465 20887 22523 20893
rect 23198 20884 23204 20896
rect 23256 20884 23262 20936
rect 25774 20884 25780 20936
rect 25832 20924 25838 20936
rect 26145 20927 26203 20933
rect 26145 20924 26157 20927
rect 25832 20896 26157 20924
rect 25832 20884 25838 20896
rect 26145 20893 26157 20896
rect 26191 20893 26203 20927
rect 26145 20887 26203 20893
rect 29549 20927 29607 20933
rect 29549 20893 29561 20927
rect 29595 20924 29607 20927
rect 29638 20924 29644 20936
rect 29595 20896 29644 20924
rect 29595 20893 29607 20896
rect 29549 20887 29607 20893
rect 29638 20884 29644 20896
rect 29696 20884 29702 20936
rect 29914 20924 29920 20936
rect 29875 20896 29920 20924
rect 29914 20884 29920 20896
rect 29972 20884 29978 20936
rect 36725 20927 36783 20933
rect 36725 20893 36737 20927
rect 36771 20924 36783 20927
rect 36998 20924 37004 20936
rect 36771 20896 37004 20924
rect 36771 20893 36783 20896
rect 36725 20887 36783 20893
rect 36998 20884 37004 20896
rect 37056 20884 37062 20936
rect 37108 20933 37136 21100
rect 38562 21088 38568 21100
rect 38620 21128 38626 21140
rect 40589 21131 40647 21137
rect 38620 21100 40448 21128
rect 38620 21088 38626 21100
rect 39224 20964 40264 20992
rect 37093 20927 37151 20933
rect 37093 20893 37105 20927
rect 37139 20893 37151 20927
rect 37093 20887 37151 20893
rect 37550 20884 37556 20936
rect 37608 20924 37614 20936
rect 38194 20924 38200 20936
rect 37608 20896 38200 20924
rect 37608 20884 37614 20896
rect 38194 20884 38200 20896
rect 38252 20924 38258 20936
rect 39224 20924 39252 20964
rect 38252 20896 39252 20924
rect 39301 20927 39359 20933
rect 38252 20884 38258 20896
rect 39301 20893 39313 20927
rect 39347 20924 39359 20927
rect 39390 20924 39396 20936
rect 39347 20896 39396 20924
rect 39347 20893 39359 20896
rect 39301 20887 39359 20893
rect 39390 20884 39396 20896
rect 39448 20884 39454 20936
rect 40236 20933 40264 20964
rect 40420 20933 40448 21100
rect 40589 21097 40601 21131
rect 40635 21128 40647 21131
rect 40862 21128 40868 21140
rect 40635 21100 40868 21128
rect 40635 21097 40647 21100
rect 40589 21091 40647 21097
rect 40862 21088 40868 21100
rect 40920 21088 40926 21140
rect 40221 20927 40279 20933
rect 40221 20893 40233 20927
rect 40267 20893 40279 20927
rect 40221 20887 40279 20893
rect 40405 20927 40463 20933
rect 40405 20893 40417 20927
rect 40451 20893 40463 20927
rect 40405 20887 40463 20893
rect 16908 20828 17356 20856
rect 16908 20816 16914 20828
rect 2498 20748 2504 20800
rect 2556 20788 2562 20800
rect 3053 20791 3111 20797
rect 3053 20788 3065 20791
rect 2556 20760 3065 20788
rect 2556 20748 2562 20760
rect 3053 20757 3065 20760
rect 3099 20788 3111 20791
rect 4982 20788 4988 20800
rect 3099 20760 4988 20788
rect 3099 20757 3111 20760
rect 3053 20751 3111 20757
rect 4982 20748 4988 20760
rect 5040 20748 5046 20800
rect 12158 20788 12164 20800
rect 12119 20760 12164 20788
rect 12158 20748 12164 20760
rect 12216 20748 12222 20800
rect 13078 20748 13084 20800
rect 13136 20788 13142 20800
rect 13173 20791 13231 20797
rect 13173 20788 13185 20791
rect 13136 20760 13185 20788
rect 13136 20748 13142 20760
rect 13173 20757 13185 20760
rect 13219 20757 13231 20791
rect 13173 20751 13231 20757
rect 13262 20748 13268 20800
rect 13320 20788 13326 20800
rect 16868 20788 16896 20816
rect 13320 20760 16896 20788
rect 17420 20788 17448 20881
rect 20254 20856 20260 20868
rect 20215 20828 20260 20856
rect 20254 20816 20260 20828
rect 20312 20816 20318 20868
rect 22738 20865 22744 20868
rect 20349 20859 20407 20865
rect 20349 20825 20361 20859
rect 20395 20825 20407 20859
rect 22732 20856 22744 20865
rect 22699 20828 22744 20856
rect 20349 20819 20407 20825
rect 22732 20819 22744 20828
rect 17494 20788 17500 20800
rect 17420 20760 17500 20788
rect 13320 20748 13326 20760
rect 17494 20748 17500 20760
rect 17552 20748 17558 20800
rect 17954 20748 17960 20800
rect 18012 20788 18018 20800
rect 19981 20791 20039 20797
rect 19981 20788 19993 20791
rect 18012 20760 19993 20788
rect 18012 20748 18018 20760
rect 19981 20757 19993 20760
rect 20027 20757 20039 20791
rect 19981 20751 20039 20757
rect 20162 20748 20168 20800
rect 20220 20788 20226 20800
rect 20364 20788 20392 20819
rect 22738 20816 22744 20819
rect 22796 20816 22802 20868
rect 23382 20816 23388 20868
rect 23440 20856 23446 20868
rect 25961 20859 26019 20865
rect 25961 20856 25973 20859
rect 23440 20828 25973 20856
rect 23440 20816 23446 20828
rect 25961 20825 25973 20828
rect 26007 20856 26019 20859
rect 28258 20856 28264 20868
rect 26007 20828 28264 20856
rect 26007 20825 26019 20828
rect 25961 20819 26019 20825
rect 28258 20816 28264 20828
rect 28316 20816 28322 20868
rect 29733 20859 29791 20865
rect 29733 20856 29745 20859
rect 29656 20828 29745 20856
rect 29656 20800 29684 20828
rect 29733 20825 29745 20828
rect 29779 20825 29791 20859
rect 29733 20819 29791 20825
rect 29825 20859 29883 20865
rect 29825 20825 29837 20859
rect 29871 20856 29883 20859
rect 31110 20856 31116 20868
rect 29871 20828 31116 20856
rect 29871 20825 29883 20828
rect 29825 20819 29883 20825
rect 31110 20816 31116 20828
rect 31168 20816 31174 20868
rect 36817 20859 36875 20865
rect 36817 20825 36829 20859
rect 36863 20825 36875 20859
rect 36817 20819 36875 20825
rect 36909 20859 36967 20865
rect 36909 20825 36921 20859
rect 36955 20856 36967 20859
rect 37182 20856 37188 20868
rect 36955 20828 37188 20856
rect 36955 20825 36967 20828
rect 36909 20819 36967 20825
rect 20220 20760 20392 20788
rect 22005 20791 22063 20797
rect 20220 20748 20226 20760
rect 22005 20757 22017 20791
rect 22051 20788 22063 20791
rect 22646 20788 22652 20800
rect 22051 20760 22652 20788
rect 22051 20757 22063 20760
rect 22005 20751 22063 20757
rect 22646 20748 22652 20760
rect 22704 20748 22710 20800
rect 23845 20791 23903 20797
rect 23845 20757 23857 20791
rect 23891 20788 23903 20791
rect 23934 20788 23940 20800
rect 23891 20760 23940 20788
rect 23891 20757 23903 20760
rect 23845 20751 23903 20757
rect 23934 20748 23940 20760
rect 23992 20788 23998 20800
rect 24486 20788 24492 20800
rect 23992 20760 24492 20788
rect 23992 20748 23998 20760
rect 24486 20748 24492 20760
rect 24544 20748 24550 20800
rect 26234 20748 26240 20800
rect 26292 20788 26298 20800
rect 26329 20791 26387 20797
rect 26329 20788 26341 20791
rect 26292 20760 26341 20788
rect 26292 20748 26298 20760
rect 26329 20757 26341 20760
rect 26375 20757 26387 20791
rect 27246 20788 27252 20800
rect 27207 20760 27252 20788
rect 26329 20751 26387 20757
rect 27246 20748 27252 20760
rect 27304 20748 27310 20800
rect 29638 20748 29644 20800
rect 29696 20748 29702 20800
rect 30098 20748 30104 20800
rect 30156 20788 30162 20800
rect 31386 20788 31392 20800
rect 30156 20760 31392 20788
rect 30156 20748 30162 20760
rect 31386 20748 31392 20760
rect 31444 20748 31450 20800
rect 32401 20791 32459 20797
rect 32401 20757 32413 20791
rect 32447 20788 32459 20791
rect 32858 20788 32864 20800
rect 32447 20760 32864 20788
rect 32447 20757 32459 20760
rect 32401 20751 32459 20757
rect 32858 20748 32864 20760
rect 32916 20748 32922 20800
rect 33318 20748 33324 20800
rect 33376 20788 33382 20800
rect 33870 20788 33876 20800
rect 33376 20760 33876 20788
rect 33376 20748 33382 20760
rect 33870 20748 33876 20760
rect 33928 20748 33934 20800
rect 36832 20788 36860 20819
rect 37182 20816 37188 20828
rect 37240 20816 37246 20868
rect 39056 20859 39114 20865
rect 39056 20825 39068 20859
rect 39102 20856 39114 20859
rect 40126 20856 40132 20868
rect 39102 20828 40132 20856
rect 39102 20825 39114 20828
rect 39056 20819 39114 20825
rect 40126 20816 40132 20828
rect 40184 20816 40190 20868
rect 37921 20791 37979 20797
rect 37921 20788 37933 20791
rect 36832 20760 37933 20788
rect 37921 20757 37933 20760
rect 37967 20788 37979 20791
rect 40402 20788 40408 20800
rect 37967 20760 40408 20788
rect 37967 20757 37979 20760
rect 37921 20751 37979 20757
rect 40402 20748 40408 20760
rect 40460 20748 40466 20800
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 7745 20587 7803 20593
rect 7745 20553 7757 20587
rect 7791 20584 7803 20587
rect 11974 20584 11980 20596
rect 7791 20556 11980 20584
rect 7791 20553 7803 20556
rect 7745 20547 7803 20553
rect 11974 20544 11980 20556
rect 12032 20544 12038 20596
rect 13630 20584 13636 20596
rect 13591 20556 13636 20584
rect 13630 20544 13636 20556
rect 13688 20544 13694 20596
rect 15654 20584 15660 20596
rect 15615 20556 15660 20584
rect 15654 20544 15660 20556
rect 15712 20544 15718 20596
rect 20162 20544 20168 20596
rect 20220 20544 20226 20596
rect 29086 20544 29092 20596
rect 29144 20584 29150 20596
rect 29362 20584 29368 20596
rect 29144 20556 29368 20584
rect 29144 20544 29150 20556
rect 29362 20544 29368 20556
rect 29420 20544 29426 20596
rect 31110 20544 31116 20596
rect 31168 20584 31174 20596
rect 31662 20584 31668 20596
rect 31168 20556 31668 20584
rect 31168 20544 31174 20556
rect 31662 20544 31668 20556
rect 31720 20584 31726 20596
rect 33597 20587 33655 20593
rect 33597 20584 33609 20587
rect 31720 20556 33609 20584
rect 31720 20544 31726 20556
rect 33597 20553 33609 20556
rect 33643 20553 33655 20587
rect 33597 20547 33655 20553
rect 40126 20544 40132 20596
rect 40184 20584 40190 20596
rect 40497 20587 40555 20593
rect 40497 20584 40509 20587
rect 40184 20556 40509 20584
rect 40184 20544 40190 20556
rect 40497 20553 40509 20556
rect 40543 20553 40555 20587
rect 40497 20547 40555 20553
rect 40770 20544 40776 20596
rect 40828 20584 40834 20596
rect 40828 20556 40908 20584
rect 40828 20544 40834 20556
rect 5350 20476 5356 20528
rect 5408 20516 5414 20528
rect 12158 20516 12164 20528
rect 5408 20488 12164 20516
rect 5408 20476 5414 20488
rect 12158 20476 12164 20488
rect 12216 20476 12222 20528
rect 13722 20516 13728 20528
rect 12406 20488 13728 20516
rect 7742 20408 7748 20460
rect 7800 20448 7806 20460
rect 7837 20451 7895 20457
rect 7837 20448 7849 20451
rect 7800 20420 7849 20448
rect 7800 20408 7806 20420
rect 7837 20417 7849 20420
rect 7883 20448 7895 20451
rect 8389 20451 8447 20457
rect 8389 20448 8401 20451
rect 7883 20420 8401 20448
rect 7883 20417 7895 20420
rect 7837 20411 7895 20417
rect 8389 20417 8401 20420
rect 8435 20417 8447 20451
rect 8389 20411 8447 20417
rect 9585 20451 9643 20457
rect 9585 20417 9597 20451
rect 9631 20448 9643 20451
rect 12406 20448 12434 20488
rect 13722 20476 13728 20488
rect 13780 20476 13786 20528
rect 19794 20516 19800 20528
rect 15580 20488 19800 20516
rect 12526 20457 12532 20460
rect 9631 20420 12434 20448
rect 9631 20417 9643 20420
rect 9585 20411 9643 20417
rect 12520 20411 12532 20457
rect 12584 20448 12590 20460
rect 12584 20420 12620 20448
rect 12526 20408 12532 20411
rect 12584 20408 12590 20420
rect 13262 20408 13268 20460
rect 13320 20448 13326 20460
rect 14369 20451 14427 20457
rect 14369 20448 14381 20451
rect 13320 20420 14381 20448
rect 13320 20408 13326 20420
rect 14369 20417 14381 20420
rect 14415 20417 14427 20451
rect 14369 20411 14427 20417
rect 15194 20408 15200 20460
rect 15252 20448 15258 20460
rect 15470 20448 15476 20460
rect 15252 20420 15476 20448
rect 15252 20408 15258 20420
rect 15470 20408 15476 20420
rect 15528 20448 15534 20460
rect 15580 20457 15608 20488
rect 19794 20476 19800 20488
rect 19852 20516 19858 20528
rect 20180 20516 20208 20544
rect 23290 20525 23296 20528
rect 20257 20519 20315 20525
rect 20257 20516 20269 20519
rect 19852 20488 20269 20516
rect 19852 20476 19858 20488
rect 20257 20485 20269 20488
rect 20303 20485 20315 20519
rect 23284 20516 23296 20525
rect 23251 20488 23296 20516
rect 20257 20479 20315 20485
rect 23284 20479 23296 20488
rect 23290 20476 23296 20479
rect 23348 20476 23354 20528
rect 27430 20516 27436 20528
rect 26068 20488 27436 20516
rect 15565 20451 15623 20457
rect 15565 20448 15577 20451
rect 15528 20420 15577 20448
rect 15528 20408 15534 20420
rect 15565 20417 15577 20420
rect 15611 20417 15623 20451
rect 17678 20448 17684 20460
rect 17639 20420 17684 20448
rect 15565 20411 15623 20417
rect 17678 20408 17684 20420
rect 17736 20408 17742 20460
rect 17773 20451 17831 20457
rect 17773 20417 17785 20451
rect 17819 20448 17831 20451
rect 19518 20448 19524 20460
rect 17819 20420 19524 20448
rect 17819 20417 17831 20420
rect 17773 20411 17831 20417
rect 19518 20408 19524 20420
rect 19576 20408 19582 20460
rect 19886 20408 19892 20460
rect 19944 20448 19950 20460
rect 20027 20451 20085 20457
rect 20027 20448 20039 20451
rect 19944 20420 20039 20448
rect 19944 20408 19950 20420
rect 20027 20417 20039 20420
rect 20073 20417 20085 20451
rect 20162 20448 20168 20460
rect 20123 20420 20168 20448
rect 20027 20411 20085 20417
rect 20162 20408 20168 20420
rect 20220 20408 20226 20460
rect 20346 20408 20352 20460
rect 20404 20457 20410 20460
rect 20404 20451 20443 20457
rect 20431 20417 20443 20451
rect 20404 20411 20443 20417
rect 20404 20408 20410 20411
rect 20530 20408 20536 20460
rect 20588 20448 20594 20460
rect 23017 20451 23075 20457
rect 20588 20420 20633 20448
rect 20588 20408 20594 20420
rect 23017 20417 23029 20451
rect 23063 20448 23075 20451
rect 23106 20448 23112 20460
rect 23063 20420 23112 20448
rect 23063 20417 23075 20420
rect 23017 20411 23075 20417
rect 23106 20408 23112 20420
rect 23164 20408 23170 20460
rect 26068 20457 26096 20488
rect 27430 20476 27436 20488
rect 27488 20476 27494 20528
rect 32398 20516 32404 20528
rect 30116 20488 32404 20516
rect 25317 20451 25375 20457
rect 25317 20417 25329 20451
rect 25363 20448 25375 20451
rect 26053 20451 26111 20457
rect 26053 20448 26065 20451
rect 25363 20420 26065 20448
rect 25363 20417 25375 20420
rect 25317 20411 25375 20417
rect 26053 20417 26065 20420
rect 26099 20417 26111 20451
rect 26053 20411 26111 20417
rect 26145 20451 26203 20457
rect 26145 20417 26157 20451
rect 26191 20417 26203 20451
rect 26145 20411 26203 20417
rect 9493 20383 9551 20389
rect 9493 20349 9505 20383
rect 9539 20380 9551 20383
rect 12250 20380 12256 20392
rect 9539 20352 10180 20380
rect 12211 20352 12256 20380
rect 9539 20349 9551 20352
rect 9493 20343 9551 20349
rect 9122 20272 9128 20324
rect 9180 20312 9186 20324
rect 9180 20284 9444 20312
rect 9180 20272 9186 20284
rect 9214 20244 9220 20256
rect 9175 20216 9220 20244
rect 9214 20204 9220 20216
rect 9272 20204 9278 20256
rect 9416 20253 9444 20284
rect 10152 20253 10180 20352
rect 12250 20340 12256 20352
rect 12308 20340 12314 20392
rect 14090 20380 14096 20392
rect 14003 20352 14096 20380
rect 14090 20340 14096 20352
rect 14148 20380 14154 20392
rect 17494 20380 17500 20392
rect 14148 20352 17500 20380
rect 14148 20340 14154 20352
rect 17494 20340 17500 20352
rect 17552 20340 17558 20392
rect 24854 20340 24860 20392
rect 24912 20380 24918 20392
rect 26160 20380 26188 20411
rect 26234 20408 26240 20460
rect 26292 20448 26298 20460
rect 26292 20420 26337 20448
rect 26292 20408 26298 20420
rect 26418 20408 26424 20460
rect 26476 20448 26482 20460
rect 26476 20420 26521 20448
rect 26476 20408 26482 20420
rect 26878 20408 26884 20460
rect 26936 20448 26942 20460
rect 27246 20448 27252 20460
rect 26936 20420 27252 20448
rect 26936 20408 26942 20420
rect 27246 20408 27252 20420
rect 27304 20448 27310 20460
rect 27525 20451 27583 20457
rect 27525 20448 27537 20451
rect 27304 20420 27537 20448
rect 27304 20408 27310 20420
rect 27525 20417 27537 20420
rect 27571 20417 27583 20451
rect 28626 20448 28632 20460
rect 28539 20420 28632 20448
rect 27525 20411 27583 20417
rect 28626 20408 28632 20420
rect 28684 20448 28690 20460
rect 29089 20451 29147 20457
rect 29089 20448 29101 20451
rect 28684 20420 29101 20448
rect 28684 20408 28690 20420
rect 29089 20417 29101 20420
rect 29135 20448 29147 20451
rect 29454 20448 29460 20460
rect 29135 20420 29460 20448
rect 29135 20417 29147 20420
rect 29089 20411 29147 20417
rect 29454 20408 29460 20420
rect 29512 20408 29518 20460
rect 30116 20457 30144 20488
rect 30101 20451 30159 20457
rect 30101 20417 30113 20451
rect 30147 20417 30159 20451
rect 31680 20448 31708 20488
rect 32398 20476 32404 20488
rect 32456 20476 32462 20528
rect 32582 20476 32588 20528
rect 32640 20516 32646 20528
rect 33137 20519 33195 20525
rect 32640 20488 32812 20516
rect 32640 20476 32646 20488
rect 31754 20448 31760 20460
rect 31680 20420 31760 20448
rect 30101 20411 30159 20417
rect 31754 20408 31760 20420
rect 31812 20408 31818 20460
rect 32030 20408 32036 20460
rect 32088 20448 32094 20460
rect 32490 20448 32496 20460
rect 32088 20420 32496 20448
rect 32088 20408 32094 20420
rect 32490 20408 32496 20420
rect 32548 20408 32554 20460
rect 32674 20448 32680 20460
rect 32635 20420 32680 20448
rect 32674 20408 32680 20420
rect 32732 20408 32738 20460
rect 32784 20457 32812 20488
rect 33137 20485 33149 20519
rect 33183 20516 33195 20519
rect 34710 20519 34768 20525
rect 34710 20516 34722 20519
rect 33183 20488 34722 20516
rect 33183 20485 33195 20488
rect 33137 20479 33195 20485
rect 34710 20485 34722 20488
rect 34756 20485 34768 20519
rect 40037 20519 40095 20525
rect 40037 20516 40049 20519
rect 34710 20479 34768 20485
rect 36096 20488 40049 20516
rect 32769 20451 32827 20457
rect 32769 20417 32781 20451
rect 32815 20417 32827 20451
rect 32769 20411 32827 20417
rect 32858 20408 32864 20460
rect 32916 20448 32922 20460
rect 36096 20448 36124 20488
rect 40037 20485 40049 20488
rect 40083 20516 40095 20519
rect 40678 20516 40684 20528
rect 40083 20488 40684 20516
rect 40083 20485 40095 20488
rect 40037 20479 40095 20485
rect 40678 20476 40684 20488
rect 40736 20516 40742 20528
rect 40736 20488 40816 20516
rect 40736 20476 40742 20488
rect 32916 20420 36124 20448
rect 36173 20451 36231 20457
rect 32916 20408 32922 20420
rect 36173 20417 36185 20451
rect 36219 20448 36231 20451
rect 36262 20448 36268 20460
rect 36219 20420 36268 20448
rect 36219 20417 36231 20420
rect 36173 20411 36231 20417
rect 36262 20408 36268 20420
rect 36320 20408 36326 20460
rect 40788 20457 40816 20488
rect 40880 20457 40908 20556
rect 40773 20451 40831 20457
rect 40773 20417 40785 20451
rect 40819 20417 40831 20451
rect 40773 20411 40831 20417
rect 40865 20451 40923 20457
rect 40865 20417 40877 20451
rect 40911 20417 40923 20451
rect 40865 20411 40923 20417
rect 40954 20408 40960 20460
rect 41012 20448 41018 20460
rect 41141 20451 41199 20457
rect 41012 20420 41057 20448
rect 41012 20408 41018 20420
rect 41141 20417 41153 20451
rect 41187 20448 41199 20451
rect 41230 20448 41236 20460
rect 41187 20420 41236 20448
rect 41187 20417 41199 20420
rect 41141 20411 41199 20417
rect 41230 20408 41236 20420
rect 41288 20408 41294 20460
rect 28442 20380 28448 20392
rect 24912 20352 28448 20380
rect 24912 20340 24918 20352
rect 28442 20340 28448 20352
rect 28500 20340 28506 20392
rect 28994 20340 29000 20392
rect 29052 20380 29058 20392
rect 29825 20383 29883 20389
rect 29825 20380 29837 20383
rect 29052 20352 29837 20380
rect 29052 20340 29058 20352
rect 29825 20349 29837 20352
rect 29871 20380 29883 20383
rect 29914 20380 29920 20392
rect 29871 20352 29920 20380
rect 29871 20349 29883 20352
rect 29825 20343 29883 20349
rect 29914 20340 29920 20352
rect 29972 20340 29978 20392
rect 34977 20383 35035 20389
rect 34977 20349 34989 20383
rect 35023 20349 35035 20383
rect 34977 20343 35035 20349
rect 35897 20383 35955 20389
rect 35897 20349 35909 20383
rect 35943 20380 35955 20383
rect 37182 20380 37188 20392
rect 35943 20352 37188 20380
rect 35943 20349 35955 20352
rect 35897 20343 35955 20349
rect 27614 20272 27620 20324
rect 27672 20312 27678 20324
rect 27709 20315 27767 20321
rect 27709 20312 27721 20315
rect 27672 20284 27721 20312
rect 27672 20272 27678 20284
rect 27709 20281 27721 20284
rect 27755 20312 27767 20315
rect 32858 20312 32864 20324
rect 27755 20284 32864 20312
rect 27755 20281 27767 20284
rect 27709 20275 27767 20281
rect 32858 20272 32864 20284
rect 32916 20272 32922 20324
rect 9401 20247 9459 20253
rect 9401 20213 9413 20247
rect 9447 20213 9459 20247
rect 9401 20207 9459 20213
rect 10137 20247 10195 20253
rect 10137 20213 10149 20247
rect 10183 20244 10195 20247
rect 11054 20244 11060 20256
rect 10183 20216 11060 20244
rect 10183 20213 10195 20216
rect 10137 20207 10195 20213
rect 11054 20204 11060 20216
rect 11112 20204 11118 20256
rect 11422 20204 11428 20256
rect 11480 20244 11486 20256
rect 11609 20247 11667 20253
rect 11609 20244 11621 20247
rect 11480 20216 11621 20244
rect 11480 20204 11486 20216
rect 11609 20213 11621 20216
rect 11655 20244 11667 20247
rect 16758 20244 16764 20256
rect 11655 20216 16764 20244
rect 11655 20213 11667 20216
rect 11609 20207 11667 20213
rect 16758 20204 16764 20216
rect 16816 20204 16822 20256
rect 16850 20204 16856 20256
rect 16908 20244 16914 20256
rect 17405 20247 17463 20253
rect 17405 20244 17417 20247
rect 16908 20216 17417 20244
rect 16908 20204 16914 20216
rect 17405 20213 17417 20216
rect 17451 20213 17463 20247
rect 17586 20244 17592 20256
rect 17547 20216 17592 20244
rect 17405 20207 17463 20213
rect 17586 20204 17592 20216
rect 17644 20204 17650 20256
rect 19889 20247 19947 20253
rect 19889 20213 19901 20247
rect 19935 20244 19947 20247
rect 19978 20244 19984 20256
rect 19935 20216 19984 20244
rect 19935 20213 19947 20216
rect 19889 20207 19947 20213
rect 19978 20204 19984 20216
rect 20036 20204 20042 20256
rect 24394 20244 24400 20256
rect 24355 20216 24400 20244
rect 24394 20204 24400 20216
rect 24452 20204 24458 20256
rect 25777 20247 25835 20253
rect 25777 20213 25789 20247
rect 25823 20244 25835 20247
rect 25866 20244 25872 20256
rect 25823 20216 25872 20244
rect 25823 20213 25835 20216
rect 25777 20207 25835 20213
rect 25866 20204 25872 20216
rect 25924 20204 25930 20256
rect 26142 20204 26148 20256
rect 26200 20244 26206 20256
rect 28994 20244 29000 20256
rect 26200 20216 29000 20244
rect 26200 20204 26206 20216
rect 28994 20204 29000 20216
rect 29052 20204 29058 20256
rect 29273 20247 29331 20253
rect 29273 20213 29285 20247
rect 29319 20244 29331 20247
rect 29362 20244 29368 20256
rect 29319 20216 29368 20244
rect 29319 20213 29331 20216
rect 29273 20207 29331 20213
rect 29362 20204 29368 20216
rect 29420 20204 29426 20256
rect 30190 20204 30196 20256
rect 30248 20244 30254 20256
rect 32214 20244 32220 20256
rect 30248 20216 32220 20244
rect 30248 20204 30254 20216
rect 32214 20204 32220 20216
rect 32272 20204 32278 20256
rect 33594 20204 33600 20256
rect 33652 20244 33658 20256
rect 34992 20244 35020 20343
rect 37182 20340 37188 20352
rect 37240 20340 37246 20392
rect 33652 20216 35020 20244
rect 33652 20204 33658 20216
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 5718 20000 5724 20052
rect 5776 20040 5782 20052
rect 11977 20043 12035 20049
rect 11977 20040 11989 20043
rect 5776 20012 11989 20040
rect 5776 20000 5782 20012
rect 11977 20009 11989 20012
rect 12023 20040 12035 20043
rect 12526 20040 12532 20052
rect 12023 20012 12434 20040
rect 12487 20012 12532 20040
rect 12023 20009 12035 20012
rect 11977 20003 12035 20009
rect 8389 19839 8447 19845
rect 8389 19805 8401 19839
rect 8435 19836 8447 19839
rect 9582 19836 9588 19848
rect 8435 19808 9588 19836
rect 8435 19805 8447 19808
rect 8389 19799 8447 19805
rect 9582 19796 9588 19808
rect 9640 19796 9646 19848
rect 12406 19836 12434 20012
rect 12526 20000 12532 20012
rect 12584 20000 12590 20052
rect 14921 20043 14979 20049
rect 14921 20009 14933 20043
rect 14967 20040 14979 20043
rect 15010 20040 15016 20052
rect 14967 20012 15016 20040
rect 14967 20009 14979 20012
rect 14921 20003 14979 20009
rect 15010 20000 15016 20012
rect 15068 20000 15074 20052
rect 19518 20040 19524 20052
rect 19479 20012 19524 20040
rect 19518 20000 19524 20012
rect 19576 20000 19582 20052
rect 22830 20000 22836 20052
rect 22888 20040 22894 20052
rect 23293 20043 23351 20049
rect 23293 20040 23305 20043
rect 22888 20012 23305 20040
rect 22888 20000 22894 20012
rect 23293 20009 23305 20012
rect 23339 20009 23351 20043
rect 25774 20040 25780 20052
rect 23293 20003 23351 20009
rect 25056 20012 25780 20040
rect 25056 19972 25084 20012
rect 25774 20000 25780 20012
rect 25832 20040 25838 20052
rect 26973 20043 27031 20049
rect 26973 20040 26985 20043
rect 25832 20012 26985 20040
rect 25832 20000 25838 20012
rect 26973 20009 26985 20012
rect 27019 20009 27031 20043
rect 26973 20003 27031 20009
rect 28736 20012 29684 20040
rect 22066 19944 25084 19972
rect 12710 19864 12716 19916
rect 12768 19904 12774 19916
rect 13262 19904 13268 19916
rect 12768 19876 13268 19904
rect 12768 19864 12774 19876
rect 12912 19845 12940 19876
rect 13262 19864 13268 19876
rect 13320 19864 13326 19916
rect 19886 19904 19892 19916
rect 19799 19876 19892 19904
rect 19886 19864 19892 19876
rect 19944 19904 19950 19916
rect 20530 19904 20536 19916
rect 19944 19876 20536 19904
rect 19944 19864 19950 19876
rect 20530 19864 20536 19876
rect 20588 19864 20594 19916
rect 12805 19839 12863 19845
rect 12805 19836 12817 19839
rect 12406 19808 12817 19836
rect 12805 19805 12817 19808
rect 12851 19805 12863 19839
rect 12805 19799 12863 19805
rect 12897 19839 12955 19845
rect 12897 19805 12909 19839
rect 12943 19805 12955 19839
rect 12897 19799 12955 19805
rect 12989 19839 13047 19845
rect 12989 19805 13001 19839
rect 13035 19836 13047 19839
rect 13078 19836 13084 19848
rect 13035 19808 13084 19836
rect 13035 19805 13047 19808
rect 12989 19799 13047 19805
rect 4798 19728 4804 19780
rect 4856 19768 4862 19780
rect 6457 19771 6515 19777
rect 6457 19768 6469 19771
rect 4856 19740 6469 19768
rect 4856 19728 4862 19740
rect 6457 19737 6469 19740
rect 6503 19737 6515 19771
rect 6457 19731 6515 19737
rect 4614 19700 4620 19712
rect 4575 19672 4620 19700
rect 4614 19660 4620 19672
rect 4672 19700 4678 19712
rect 5350 19700 5356 19712
rect 4672 19672 5356 19700
rect 4672 19660 4678 19672
rect 5350 19660 5356 19672
rect 5408 19700 5414 19712
rect 5905 19703 5963 19709
rect 5905 19700 5917 19703
rect 5408 19672 5917 19700
rect 5408 19660 5414 19672
rect 5905 19669 5917 19672
rect 5951 19669 5963 19703
rect 6472 19700 6500 19731
rect 7834 19728 7840 19780
rect 7892 19768 7898 19780
rect 8122 19771 8180 19777
rect 8122 19768 8134 19771
rect 7892 19740 8134 19768
rect 7892 19728 7898 19740
rect 8122 19737 8134 19740
rect 8168 19737 8180 19771
rect 12820 19768 12848 19799
rect 13078 19796 13084 19808
rect 13136 19796 13142 19848
rect 13170 19796 13176 19848
rect 13228 19836 13234 19848
rect 14826 19836 14832 19848
rect 13228 19808 13273 19836
rect 14787 19808 14832 19836
rect 13228 19796 13234 19808
rect 14826 19796 14832 19808
rect 14884 19796 14890 19848
rect 14921 19839 14979 19845
rect 14921 19805 14933 19839
rect 14967 19836 14979 19839
rect 17954 19836 17960 19848
rect 14967 19808 17960 19836
rect 14967 19805 14979 19808
rect 14921 19799 14979 19805
rect 17954 19796 17960 19808
rect 18012 19796 18018 19848
rect 19700 19839 19758 19845
rect 19700 19805 19712 19839
rect 19746 19836 19758 19839
rect 19904 19836 19932 19864
rect 20070 19836 20076 19848
rect 19746 19808 19932 19836
rect 20031 19808 20076 19836
rect 19746 19805 19758 19808
rect 19700 19799 19758 19805
rect 20070 19796 20076 19808
rect 20128 19796 20134 19848
rect 20165 19839 20223 19845
rect 20165 19805 20177 19839
rect 20211 19836 20223 19839
rect 21174 19836 21180 19848
rect 20211 19808 21180 19836
rect 20211 19805 20223 19808
rect 20165 19799 20223 19805
rect 21174 19796 21180 19808
rect 21232 19796 21238 19848
rect 13722 19768 13728 19780
rect 12820 19740 13728 19768
rect 8122 19731 8180 19737
rect 13722 19728 13728 19740
rect 13780 19728 13786 19780
rect 19797 19771 19855 19777
rect 19797 19737 19809 19771
rect 19843 19737 19855 19771
rect 19797 19731 19855 19737
rect 7009 19703 7067 19709
rect 7009 19700 7021 19703
rect 6472 19672 7021 19700
rect 5905 19663 5963 19669
rect 7009 19669 7021 19672
rect 7055 19700 7067 19703
rect 7650 19700 7656 19712
rect 7055 19672 7656 19700
rect 7055 19669 7067 19672
rect 7009 19663 7067 19669
rect 7650 19660 7656 19672
rect 7708 19660 7714 19712
rect 14553 19703 14611 19709
rect 14553 19669 14565 19703
rect 14599 19700 14611 19703
rect 15010 19700 15016 19712
rect 14599 19672 15016 19700
rect 14599 19669 14611 19672
rect 14553 19663 14611 19669
rect 15010 19660 15016 19672
rect 15068 19660 15074 19712
rect 19812 19700 19840 19731
rect 19886 19728 19892 19780
rect 19944 19768 19950 19780
rect 22066 19768 22094 19944
rect 26970 19864 26976 19916
rect 27028 19864 27034 19916
rect 23477 19839 23535 19845
rect 23477 19805 23489 19839
rect 23523 19836 23535 19839
rect 24394 19836 24400 19848
rect 23523 19808 24400 19836
rect 23523 19805 23535 19808
rect 23477 19799 23535 19805
rect 24394 19796 24400 19808
rect 24452 19796 24458 19848
rect 25593 19839 25651 19845
rect 25593 19805 25605 19839
rect 25639 19836 25651 19839
rect 25682 19836 25688 19848
rect 25639 19808 25688 19836
rect 25639 19805 25651 19808
rect 25593 19799 25651 19805
rect 25682 19796 25688 19808
rect 25740 19796 25746 19848
rect 25866 19845 25872 19848
rect 25860 19836 25872 19845
rect 25827 19808 25872 19836
rect 25860 19799 25872 19808
rect 25866 19796 25872 19799
rect 25924 19796 25930 19848
rect 26988 19836 27016 19864
rect 28736 19845 28764 20012
rect 29656 19972 29684 20012
rect 29730 20000 29736 20052
rect 29788 20040 29794 20052
rect 29871 20043 29929 20049
rect 29871 20040 29883 20043
rect 29788 20012 29883 20040
rect 29788 20000 29794 20012
rect 29871 20009 29883 20012
rect 29917 20040 29929 20043
rect 32122 20040 32128 20052
rect 29917 20012 32128 20040
rect 29917 20009 29929 20012
rect 29871 20003 29929 20009
rect 32122 20000 32128 20012
rect 32180 20000 32186 20052
rect 32674 20000 32680 20052
rect 32732 20040 32738 20052
rect 33137 20043 33195 20049
rect 33137 20040 33149 20043
rect 32732 20012 33149 20040
rect 32732 20000 32738 20012
rect 33137 20009 33149 20012
rect 33183 20009 33195 20043
rect 33137 20003 33195 20009
rect 35342 20000 35348 20052
rect 35400 20040 35406 20052
rect 36078 20040 36084 20052
rect 35400 20012 36084 20040
rect 35400 20000 35406 20012
rect 36078 20000 36084 20012
rect 36136 20040 36142 20052
rect 36403 20043 36461 20049
rect 36403 20040 36415 20043
rect 36136 20012 36415 20040
rect 36136 20000 36142 20012
rect 36403 20009 36415 20012
rect 36449 20009 36461 20043
rect 36403 20003 36461 20009
rect 40589 20043 40647 20049
rect 40589 20009 40601 20043
rect 40635 20040 40647 20043
rect 40954 20040 40960 20052
rect 40635 20012 40960 20040
rect 40635 20009 40647 20012
rect 40589 20003 40647 20009
rect 40954 20000 40960 20012
rect 41012 20000 41018 20052
rect 30190 19972 30196 19984
rect 29656 19944 30196 19972
rect 30190 19932 30196 19944
rect 30248 19932 30254 19984
rect 31110 19972 31116 19984
rect 30300 19944 31116 19972
rect 28445 19839 28503 19845
rect 28445 19836 28457 19839
rect 26988 19808 28457 19836
rect 28445 19805 28457 19808
rect 28491 19805 28503 19839
rect 28445 19799 28503 19805
rect 28721 19839 28779 19845
rect 28721 19805 28733 19839
rect 28767 19805 28779 19839
rect 28721 19799 28779 19805
rect 28813 19839 28871 19845
rect 28813 19805 28825 19839
rect 28859 19836 28871 19839
rect 28994 19836 29000 19848
rect 28859 19808 29000 19836
rect 28859 19805 28871 19808
rect 28813 19799 28871 19805
rect 28994 19796 29000 19808
rect 29052 19796 29058 19848
rect 29638 19836 29644 19848
rect 29551 19808 29644 19836
rect 29638 19796 29644 19808
rect 29696 19796 29702 19848
rect 23658 19768 23664 19780
rect 19944 19740 19989 19768
rect 20916 19740 22094 19768
rect 23619 19740 23664 19768
rect 19944 19728 19950 19740
rect 20916 19700 20944 19740
rect 23658 19728 23664 19740
rect 23716 19728 23722 19780
rect 24670 19728 24676 19780
rect 24728 19768 24734 19780
rect 28629 19771 28687 19777
rect 28629 19768 28641 19771
rect 24728 19740 28641 19768
rect 24728 19728 24734 19740
rect 28629 19737 28641 19740
rect 28675 19768 28687 19771
rect 29656 19768 29684 19796
rect 28675 19740 29684 19768
rect 28675 19737 28687 19740
rect 28629 19731 28687 19737
rect 19812 19672 20944 19700
rect 21082 19660 21088 19712
rect 21140 19700 21146 19712
rect 25866 19700 25872 19712
rect 21140 19672 25872 19700
rect 21140 19660 21146 19672
rect 25866 19660 25872 19672
rect 25924 19660 25930 19712
rect 26418 19660 26424 19712
rect 26476 19700 26482 19712
rect 27433 19703 27491 19709
rect 27433 19700 27445 19703
rect 26476 19672 27445 19700
rect 26476 19660 26482 19672
rect 27433 19669 27445 19672
rect 27479 19700 27491 19703
rect 27614 19700 27620 19712
rect 27479 19672 27620 19700
rect 27479 19669 27491 19672
rect 27433 19663 27491 19669
rect 27614 19660 27620 19672
rect 27672 19660 27678 19712
rect 28997 19703 29055 19709
rect 28997 19669 29009 19703
rect 29043 19700 29055 19703
rect 30300 19700 30328 19944
rect 31110 19932 31116 19944
rect 31168 19932 31174 19984
rect 37826 19972 37832 19984
rect 35728 19944 37832 19972
rect 31754 19904 31760 19916
rect 31128 19876 31760 19904
rect 30466 19796 30472 19848
rect 30524 19836 30530 19848
rect 31128 19845 31156 19876
rect 31754 19864 31760 19876
rect 31812 19864 31818 19916
rect 31113 19839 31171 19845
rect 31113 19836 31125 19839
rect 30524 19808 31125 19836
rect 30524 19796 30530 19808
rect 31113 19805 31125 19808
rect 31159 19805 31171 19839
rect 31478 19836 31484 19848
rect 31439 19808 31484 19836
rect 31113 19799 31171 19805
rect 31478 19796 31484 19808
rect 31536 19796 31542 19848
rect 31662 19796 31668 19848
rect 31720 19836 31726 19848
rect 32953 19839 33011 19845
rect 32953 19836 32965 19839
rect 31720 19808 32965 19836
rect 31720 19796 31726 19808
rect 32953 19805 32965 19808
rect 32999 19805 33011 19839
rect 35342 19836 35348 19848
rect 35303 19808 35348 19836
rect 32953 19799 33011 19805
rect 35342 19796 35348 19808
rect 35400 19796 35406 19848
rect 35728 19845 35756 19944
rect 37826 19932 37832 19944
rect 37884 19932 37890 19984
rect 35713 19839 35771 19845
rect 35713 19805 35725 19839
rect 35759 19805 35771 19839
rect 35713 19799 35771 19805
rect 36173 19839 36231 19845
rect 36173 19805 36185 19839
rect 36219 19836 36231 19839
rect 36998 19836 37004 19848
rect 36219 19808 37004 19836
rect 36219 19805 36231 19808
rect 36173 19799 36231 19805
rect 36998 19796 37004 19808
rect 37056 19796 37062 19848
rect 39298 19836 39304 19848
rect 39259 19808 39304 19836
rect 39298 19796 39304 19808
rect 39356 19796 39362 19848
rect 39850 19796 39856 19848
rect 39908 19836 39914 19848
rect 40221 19839 40279 19845
rect 40221 19836 40233 19839
rect 39908 19808 40233 19836
rect 39908 19796 39914 19808
rect 40221 19805 40233 19808
rect 40267 19805 40279 19839
rect 40402 19836 40408 19848
rect 40363 19808 40408 19836
rect 40221 19799 40279 19805
rect 40402 19796 40408 19808
rect 40460 19796 40466 19848
rect 58158 19836 58164 19848
rect 58119 19808 58164 19836
rect 58158 19796 58164 19808
rect 58216 19796 58222 19848
rect 31202 19768 31208 19780
rect 31163 19740 31208 19768
rect 31202 19728 31208 19740
rect 31260 19728 31266 19780
rect 31297 19771 31355 19777
rect 31297 19737 31309 19771
rect 31343 19768 31355 19771
rect 32122 19768 32128 19780
rect 31343 19740 32128 19768
rect 31343 19737 31355 19740
rect 31297 19731 31355 19737
rect 32122 19728 32128 19740
rect 32180 19728 32186 19780
rect 32766 19768 32772 19780
rect 32727 19740 32772 19768
rect 32766 19728 32772 19740
rect 32824 19728 32830 19780
rect 35437 19771 35495 19777
rect 35437 19737 35449 19771
rect 35483 19737 35495 19771
rect 35437 19731 35495 19737
rect 35529 19771 35587 19777
rect 35529 19737 35541 19771
rect 35575 19768 35587 19771
rect 36262 19768 36268 19780
rect 35575 19740 36268 19768
rect 35575 19737 35587 19740
rect 35529 19731 35587 19737
rect 30926 19700 30932 19712
rect 29043 19672 30328 19700
rect 30887 19672 30932 19700
rect 29043 19669 29055 19672
rect 28997 19663 29055 19669
rect 30926 19660 30932 19672
rect 30984 19660 30990 19712
rect 34514 19660 34520 19712
rect 34572 19700 34578 19712
rect 35161 19703 35219 19709
rect 35161 19700 35173 19703
rect 34572 19672 35173 19700
rect 34572 19660 34578 19672
rect 35161 19669 35173 19672
rect 35207 19669 35219 19703
rect 35452 19700 35480 19731
rect 36262 19728 36268 19740
rect 36320 19728 36326 19780
rect 39056 19771 39114 19777
rect 39056 19737 39068 19771
rect 39102 19768 39114 19771
rect 40126 19768 40132 19780
rect 39102 19740 40132 19768
rect 39102 19737 39114 19740
rect 39056 19731 39114 19737
rect 40126 19728 40132 19740
rect 40184 19728 40190 19780
rect 37366 19700 37372 19712
rect 35452 19672 37372 19700
rect 35161 19663 35219 19669
rect 37366 19660 37372 19672
rect 37424 19660 37430 19712
rect 37918 19700 37924 19712
rect 37879 19672 37924 19700
rect 37918 19660 37924 19672
rect 37976 19660 37982 19712
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 5718 19456 5724 19508
rect 5776 19496 5782 19508
rect 6549 19499 6607 19505
rect 6549 19496 6561 19499
rect 5776 19468 6561 19496
rect 5776 19456 5782 19468
rect 6549 19465 6561 19468
rect 6595 19465 6607 19499
rect 7834 19496 7840 19508
rect 7795 19468 7840 19496
rect 6549 19459 6607 19465
rect 7834 19456 7840 19468
rect 7892 19456 7898 19508
rect 14090 19496 14096 19508
rect 14051 19468 14096 19496
rect 14090 19456 14096 19468
rect 14148 19456 14154 19508
rect 16758 19456 16764 19508
rect 16816 19496 16822 19508
rect 17586 19496 17592 19508
rect 16816 19468 17592 19496
rect 16816 19456 16822 19468
rect 17586 19456 17592 19468
rect 17644 19456 17650 19508
rect 18046 19496 18052 19508
rect 17959 19468 18052 19496
rect 18046 19456 18052 19468
rect 18104 19496 18110 19508
rect 21082 19496 21088 19508
rect 18104 19468 21088 19496
rect 18104 19456 18110 19468
rect 21082 19456 21088 19468
rect 21140 19456 21146 19508
rect 21910 19456 21916 19508
rect 21968 19496 21974 19508
rect 22005 19499 22063 19505
rect 22005 19496 22017 19499
rect 21968 19468 22017 19496
rect 21968 19456 21974 19468
rect 22005 19465 22017 19468
rect 22051 19496 22063 19499
rect 23014 19496 23020 19508
rect 22051 19468 23020 19496
rect 22051 19465 22063 19468
rect 22005 19459 22063 19465
rect 23014 19456 23020 19468
rect 23072 19456 23078 19508
rect 25961 19499 26019 19505
rect 25961 19465 25973 19499
rect 26007 19496 26019 19499
rect 26694 19496 26700 19508
rect 26007 19468 26700 19496
rect 26007 19465 26019 19468
rect 25961 19459 26019 19465
rect 26694 19456 26700 19468
rect 26752 19456 26758 19508
rect 26970 19496 26976 19508
rect 26931 19468 26976 19496
rect 26970 19456 26976 19468
rect 27028 19456 27034 19508
rect 35897 19499 35955 19505
rect 35897 19496 35909 19499
rect 30852 19468 35909 19496
rect 5350 19388 5356 19440
rect 5408 19428 5414 19440
rect 6457 19431 6515 19437
rect 6457 19428 6469 19431
rect 5408 19400 6469 19428
rect 5408 19388 5414 19400
rect 6457 19397 6469 19400
rect 6503 19397 6515 19431
rect 9214 19428 9220 19440
rect 6457 19391 6515 19397
rect 7300 19400 9220 19428
rect 2406 19360 2412 19372
rect 2367 19332 2412 19360
rect 2406 19320 2412 19332
rect 2464 19320 2470 19372
rect 4617 19363 4675 19369
rect 4617 19329 4629 19363
rect 4663 19360 4675 19363
rect 4706 19360 4712 19372
rect 4663 19332 4712 19360
rect 4663 19329 4675 19332
rect 4617 19323 4675 19329
rect 4706 19320 4712 19332
rect 4764 19360 4770 19372
rect 5445 19363 5503 19369
rect 5445 19360 5457 19363
rect 4764 19332 5457 19360
rect 4764 19320 4770 19332
rect 5445 19329 5457 19332
rect 5491 19329 5503 19363
rect 5445 19323 5503 19329
rect 6914 19320 6920 19372
rect 6972 19360 6978 19372
rect 7300 19369 7328 19400
rect 9214 19388 9220 19400
rect 9272 19388 9278 19440
rect 13814 19388 13820 19440
rect 13872 19428 13878 19440
rect 14645 19431 14703 19437
rect 14645 19428 14657 19431
rect 13872 19400 14657 19428
rect 13872 19388 13878 19400
rect 7101 19363 7159 19369
rect 7101 19360 7113 19363
rect 6972 19332 7113 19360
rect 6972 19320 6978 19332
rect 7101 19329 7113 19332
rect 7147 19329 7159 19363
rect 7101 19323 7159 19329
rect 7285 19363 7343 19369
rect 7285 19329 7297 19363
rect 7331 19329 7343 19363
rect 7650 19360 7656 19372
rect 7611 19332 7656 19360
rect 7285 19323 7343 19329
rect 7650 19320 7656 19332
rect 7708 19320 7714 19372
rect 8665 19363 8723 19369
rect 8665 19329 8677 19363
rect 8711 19360 8723 19363
rect 11974 19360 11980 19372
rect 8711 19332 11980 19360
rect 8711 19329 8723 19332
rect 8665 19323 8723 19329
rect 11974 19320 11980 19332
rect 12032 19320 12038 19372
rect 14200 19369 14228 19400
rect 14645 19397 14657 19400
rect 14691 19428 14703 19431
rect 14691 19400 21956 19428
rect 14691 19397 14703 19400
rect 14645 19391 14703 19397
rect 14001 19363 14059 19369
rect 14001 19329 14013 19363
rect 14047 19329 14059 19363
rect 14001 19323 14059 19329
rect 14185 19363 14243 19369
rect 14185 19329 14197 19363
rect 14231 19329 14243 19363
rect 16666 19360 16672 19372
rect 16627 19332 16672 19360
rect 14185 19323 14243 19329
rect 5626 19252 5632 19304
rect 5684 19292 5690 19304
rect 7377 19295 7435 19301
rect 7377 19292 7389 19295
rect 5684 19264 7389 19292
rect 5684 19252 5690 19264
rect 7377 19261 7389 19264
rect 7423 19261 7435 19295
rect 7377 19255 7435 19261
rect 7469 19295 7527 19301
rect 7469 19261 7481 19295
rect 7515 19261 7527 19295
rect 8573 19295 8631 19301
rect 7469 19255 7527 19261
rect 7944 19264 8524 19292
rect 4890 19184 4896 19236
rect 4948 19224 4954 19236
rect 4948 19196 7236 19224
rect 4948 19184 4954 19196
rect 2130 19116 2136 19168
rect 2188 19156 2194 19168
rect 2225 19159 2283 19165
rect 2225 19156 2237 19159
rect 2188 19128 2237 19156
rect 2188 19116 2194 19128
rect 2225 19125 2237 19128
rect 2271 19125 2283 19159
rect 2225 19119 2283 19125
rect 5353 19159 5411 19165
rect 5353 19125 5365 19159
rect 5399 19156 5411 19159
rect 5442 19156 5448 19168
rect 5399 19128 5448 19156
rect 5399 19125 5411 19128
rect 5353 19119 5411 19125
rect 5442 19116 5448 19128
rect 5500 19116 5506 19168
rect 7208 19156 7236 19196
rect 7282 19184 7288 19236
rect 7340 19224 7346 19236
rect 7484 19224 7512 19255
rect 7340 19196 7512 19224
rect 7340 19184 7346 19196
rect 7944 19156 7972 19264
rect 8202 19184 8208 19236
rect 8260 19224 8266 19236
rect 8496 19224 8524 19264
rect 8573 19261 8585 19295
rect 8619 19292 8631 19295
rect 9217 19295 9275 19301
rect 9217 19292 9229 19295
rect 8619 19264 9229 19292
rect 8619 19261 8631 19264
rect 8573 19255 8631 19261
rect 9217 19261 9229 19264
rect 9263 19292 9275 19295
rect 13906 19292 13912 19304
rect 9263 19264 13912 19292
rect 9263 19261 9275 19264
rect 9217 19255 9275 19261
rect 13906 19252 13912 19264
rect 13964 19252 13970 19304
rect 14016 19292 14044 19323
rect 16666 19320 16672 19332
rect 16724 19320 16730 19372
rect 16758 19320 16764 19372
rect 16816 19360 16822 19372
rect 21928 19369 21956 19400
rect 24670 19388 24676 19440
rect 24728 19428 24734 19440
rect 25593 19431 25651 19437
rect 25593 19428 25605 19431
rect 24728 19400 25605 19428
rect 24728 19388 24734 19400
rect 25593 19397 25605 19400
rect 25639 19397 25651 19431
rect 25593 19391 25651 19397
rect 25866 19388 25872 19440
rect 25924 19428 25930 19440
rect 27433 19431 27491 19437
rect 25924 19400 27384 19428
rect 25924 19388 25930 19400
rect 16925 19363 16983 19369
rect 16925 19360 16937 19363
rect 16816 19332 16937 19360
rect 16816 19320 16822 19332
rect 16925 19329 16937 19332
rect 16971 19329 16983 19363
rect 16925 19323 16983 19329
rect 21913 19363 21971 19369
rect 21913 19329 21925 19363
rect 21959 19329 21971 19363
rect 21913 19323 21971 19329
rect 14550 19292 14556 19304
rect 14016 19264 14556 19292
rect 14550 19252 14556 19264
rect 14608 19252 14614 19304
rect 21928 19292 21956 19323
rect 22094 19320 22100 19372
rect 22152 19360 22158 19372
rect 22152 19332 22197 19360
rect 22152 19320 22158 19332
rect 24394 19320 24400 19372
rect 24452 19360 24458 19372
rect 25409 19363 25467 19369
rect 25409 19360 25421 19363
rect 24452 19332 25421 19360
rect 24452 19320 24458 19332
rect 25409 19329 25421 19332
rect 25455 19329 25467 19363
rect 25682 19360 25688 19372
rect 25643 19332 25688 19360
rect 25409 19323 25467 19329
rect 25682 19320 25688 19332
rect 25740 19320 25746 19372
rect 25777 19363 25835 19369
rect 25777 19329 25789 19363
rect 25823 19360 25835 19363
rect 26142 19360 26148 19372
rect 25823 19332 26148 19360
rect 25823 19329 25835 19332
rect 25777 19323 25835 19329
rect 22370 19292 22376 19304
rect 21928 19264 22376 19292
rect 22370 19252 22376 19264
rect 22428 19292 22434 19304
rect 22557 19295 22615 19301
rect 22557 19292 22569 19295
rect 22428 19264 22569 19292
rect 22428 19252 22434 19264
rect 22557 19261 22569 19264
rect 22603 19261 22615 19295
rect 22557 19255 22615 19261
rect 24946 19252 24952 19304
rect 25004 19292 25010 19304
rect 25792 19292 25820 19323
rect 26142 19320 26148 19332
rect 26200 19320 26206 19372
rect 26418 19320 26424 19372
rect 26476 19360 26482 19372
rect 26476 19332 27108 19360
rect 26476 19320 26482 19332
rect 25004 19264 25820 19292
rect 27080 19292 27108 19332
rect 27154 19320 27160 19372
rect 27212 19360 27218 19372
rect 27356 19360 27384 19400
rect 27433 19397 27445 19431
rect 27479 19428 27491 19431
rect 27522 19428 27528 19440
rect 27479 19400 27528 19428
rect 27479 19397 27491 19400
rect 27433 19391 27491 19397
rect 27522 19388 27528 19400
rect 27580 19388 27586 19440
rect 29730 19428 29736 19440
rect 29691 19400 29736 19428
rect 29730 19388 29736 19400
rect 29788 19388 29794 19440
rect 30374 19388 30380 19440
rect 30432 19428 30438 19440
rect 30852 19428 30880 19468
rect 35897 19465 35909 19468
rect 35943 19465 35955 19499
rect 39298 19496 39304 19508
rect 35897 19459 35955 19465
rect 36004 19468 39304 19496
rect 31018 19428 31024 19440
rect 30432 19400 30880 19428
rect 30979 19400 31024 19428
rect 30432 19388 30438 19400
rect 31018 19388 31024 19400
rect 31076 19388 31082 19440
rect 34422 19428 34428 19440
rect 31726 19400 34428 19428
rect 29549 19363 29607 19369
rect 29549 19360 29561 19363
rect 27212 19332 27257 19360
rect 27356 19332 29561 19360
rect 27212 19320 27218 19332
rect 29549 19329 29561 19332
rect 29595 19329 29607 19363
rect 29822 19360 29828 19372
rect 29783 19332 29828 19360
rect 29549 19323 29607 19329
rect 29822 19320 29828 19332
rect 29880 19320 29886 19372
rect 29917 19363 29975 19369
rect 29917 19329 29929 19363
rect 29963 19360 29975 19363
rect 30466 19360 30472 19372
rect 29963 19332 30472 19360
rect 29963 19329 29975 19332
rect 29917 19323 29975 19329
rect 30466 19320 30472 19332
rect 30524 19320 30530 19372
rect 30745 19363 30803 19369
rect 30745 19329 30757 19363
rect 30791 19360 30803 19363
rect 31726 19360 31754 19400
rect 34422 19388 34428 19400
rect 34480 19388 34486 19440
rect 36004 19428 36032 19468
rect 39298 19456 39304 19468
rect 39356 19456 39362 19508
rect 40126 19456 40132 19508
rect 40184 19496 40190 19508
rect 40589 19499 40647 19505
rect 40589 19496 40601 19499
rect 40184 19468 40601 19496
rect 40184 19456 40190 19468
rect 40589 19465 40601 19468
rect 40635 19465 40647 19499
rect 40589 19459 40647 19465
rect 36262 19428 36268 19440
rect 35912 19400 36032 19428
rect 36223 19400 36268 19428
rect 35912 19372 35940 19400
rect 36262 19388 36268 19400
rect 36320 19388 36326 19440
rect 38102 19428 38108 19440
rect 36372 19400 38108 19428
rect 33318 19360 33324 19372
rect 33376 19369 33382 19372
rect 30791 19332 31754 19360
rect 33288 19332 33324 19360
rect 30791 19329 30803 19332
rect 30745 19323 30803 19329
rect 33318 19320 33324 19332
rect 33376 19323 33388 19369
rect 33594 19360 33600 19372
rect 33555 19332 33600 19360
rect 33376 19320 33382 19323
rect 33594 19320 33600 19332
rect 33652 19360 33658 19372
rect 35894 19360 35900 19372
rect 33652 19332 35900 19360
rect 33652 19320 33658 19332
rect 35894 19320 35900 19332
rect 35952 19320 35958 19372
rect 36078 19360 36084 19372
rect 36039 19332 36084 19360
rect 36078 19320 36084 19332
rect 36136 19320 36142 19372
rect 36173 19363 36231 19369
rect 36173 19329 36185 19363
rect 36219 19360 36231 19363
rect 36372 19360 36400 19400
rect 38102 19388 38108 19400
rect 38160 19388 38166 19440
rect 40678 19388 40684 19440
rect 40736 19428 40742 19440
rect 40736 19400 41000 19428
rect 40736 19388 40742 19400
rect 36219 19332 36400 19360
rect 36449 19363 36507 19369
rect 36219 19329 36231 19332
rect 36173 19323 36231 19329
rect 36449 19329 36461 19363
rect 36495 19360 36507 19363
rect 37274 19360 37280 19372
rect 36495 19332 37280 19360
rect 36495 19329 36507 19332
rect 36449 19323 36507 19329
rect 37274 19320 37280 19332
rect 37332 19320 37338 19372
rect 37553 19363 37611 19369
rect 37553 19329 37565 19363
rect 37599 19360 37611 19363
rect 37642 19360 37648 19372
rect 37599 19332 37648 19360
rect 37599 19329 37611 19332
rect 37553 19323 37611 19329
rect 37642 19320 37648 19332
rect 37700 19360 37706 19372
rect 38013 19363 38071 19369
rect 38013 19360 38025 19363
rect 37700 19332 38025 19360
rect 37700 19320 37706 19332
rect 38013 19329 38025 19332
rect 38059 19329 38071 19363
rect 40862 19360 40868 19372
rect 40823 19332 40868 19360
rect 38013 19323 38071 19329
rect 40862 19320 40868 19332
rect 40920 19320 40926 19372
rect 40972 19369 41000 19400
rect 40957 19363 41015 19369
rect 40957 19329 40969 19363
rect 41003 19329 41015 19363
rect 40957 19323 41015 19329
rect 41046 19320 41052 19372
rect 41104 19360 41110 19372
rect 41104 19332 41149 19360
rect 41104 19320 41110 19332
rect 41230 19320 41236 19372
rect 41288 19360 41294 19372
rect 41288 19332 41333 19360
rect 41288 19320 41294 19332
rect 27249 19295 27307 19301
rect 27249 19292 27261 19295
rect 27080 19264 27261 19292
rect 25004 19252 25010 19264
rect 27249 19261 27261 19264
rect 27295 19261 27307 19295
rect 30834 19292 30840 19304
rect 27249 19255 27307 19261
rect 30484 19264 30696 19292
rect 30795 19264 30840 19292
rect 8260 19196 8432 19224
rect 8496 19196 8800 19224
rect 8260 19184 8266 19196
rect 8294 19156 8300 19168
rect 7208 19128 7972 19156
rect 8255 19128 8300 19156
rect 8294 19116 8300 19128
rect 8352 19116 8358 19168
rect 8404 19156 8432 19196
rect 8481 19159 8539 19165
rect 8481 19156 8493 19159
rect 8404 19128 8493 19156
rect 8481 19125 8493 19128
rect 8527 19125 8539 19159
rect 8772 19156 8800 19196
rect 10778 19184 10784 19236
rect 10836 19224 10842 19236
rect 10836 19196 11008 19224
rect 10836 19184 10842 19196
rect 10686 19156 10692 19168
rect 8772 19128 10692 19156
rect 8481 19119 8539 19125
rect 10686 19116 10692 19128
rect 10744 19156 10750 19168
rect 10873 19159 10931 19165
rect 10873 19156 10885 19159
rect 10744 19128 10885 19156
rect 10744 19116 10750 19128
rect 10873 19125 10885 19128
rect 10919 19125 10931 19159
rect 10980 19156 11008 19196
rect 11054 19184 11060 19236
rect 11112 19224 11118 19236
rect 11112 19196 16712 19224
rect 11112 19184 11118 19196
rect 11517 19159 11575 19165
rect 11517 19156 11529 19159
rect 10980 19128 11529 19156
rect 10873 19119 10931 19125
rect 11517 19125 11529 19128
rect 11563 19125 11575 19159
rect 11517 19119 11575 19125
rect 11606 19116 11612 19168
rect 11664 19156 11670 19168
rect 12710 19156 12716 19168
rect 11664 19128 12716 19156
rect 11664 19116 11670 19128
rect 12710 19116 12716 19128
rect 12768 19116 12774 19168
rect 16684 19156 16712 19196
rect 20622 19184 20628 19236
rect 20680 19224 20686 19236
rect 30484 19224 30512 19264
rect 20680 19196 30512 19224
rect 30668 19224 30696 19264
rect 30834 19252 30840 19264
rect 30892 19252 30898 19304
rect 31478 19224 31484 19236
rect 30668 19196 31484 19224
rect 20680 19184 20686 19196
rect 31478 19184 31484 19196
rect 31536 19184 31542 19236
rect 32214 19224 32220 19236
rect 32175 19196 32220 19224
rect 32214 19184 32220 19196
rect 32272 19184 32278 19236
rect 19242 19156 19248 19168
rect 16684 19128 19248 19156
rect 19242 19116 19248 19128
rect 19300 19116 19306 19168
rect 27338 19156 27344 19168
rect 27299 19128 27344 19156
rect 27338 19116 27344 19128
rect 27396 19116 27402 19168
rect 30101 19159 30159 19165
rect 30101 19125 30113 19159
rect 30147 19156 30159 19159
rect 30466 19156 30472 19168
rect 30147 19128 30472 19156
rect 30147 19125 30159 19128
rect 30101 19119 30159 19125
rect 30466 19116 30472 19128
rect 30524 19116 30530 19168
rect 30561 19159 30619 19165
rect 30561 19125 30573 19159
rect 30607 19156 30619 19159
rect 30650 19156 30656 19168
rect 30607 19128 30656 19156
rect 30607 19125 30619 19128
rect 30561 19119 30619 19125
rect 30650 19116 30656 19128
rect 30708 19116 30714 19168
rect 31021 19159 31079 19165
rect 31021 19125 31033 19159
rect 31067 19156 31079 19159
rect 31110 19156 31116 19168
rect 31067 19128 31116 19156
rect 31067 19125 31079 19128
rect 31021 19119 31079 19125
rect 31110 19116 31116 19128
rect 31168 19116 31174 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 5626 18952 5632 18964
rect 5587 18924 5632 18952
rect 5626 18912 5632 18924
rect 5684 18912 5690 18964
rect 6365 18955 6423 18961
rect 6365 18921 6377 18955
rect 6411 18952 6423 18955
rect 6822 18952 6828 18964
rect 6411 18924 6828 18952
rect 6411 18921 6423 18924
rect 6365 18915 6423 18921
rect 6822 18912 6828 18924
rect 6880 18952 6886 18964
rect 12526 18952 12532 18964
rect 6880 18924 12532 18952
rect 6880 18912 6886 18924
rect 12526 18912 12532 18924
rect 12584 18952 12590 18964
rect 13630 18952 13636 18964
rect 12584 18924 13636 18952
rect 12584 18912 12590 18924
rect 13630 18912 13636 18924
rect 13688 18952 13694 18964
rect 15838 18952 15844 18964
rect 13688 18924 15844 18952
rect 13688 18912 13694 18924
rect 15838 18912 15844 18924
rect 15896 18912 15902 18964
rect 16393 18955 16451 18961
rect 16393 18921 16405 18955
rect 16439 18952 16451 18955
rect 16758 18952 16764 18964
rect 16439 18924 16764 18952
rect 16439 18921 16451 18924
rect 16393 18915 16451 18921
rect 16758 18912 16764 18924
rect 16816 18912 16822 18964
rect 20622 18952 20628 18964
rect 20583 18924 20628 18952
rect 20622 18912 20628 18924
rect 20680 18912 20686 18964
rect 26694 18912 26700 18964
rect 26752 18952 26758 18964
rect 27338 18952 27344 18964
rect 26752 18924 27344 18952
rect 26752 18912 26758 18924
rect 27338 18912 27344 18924
rect 27396 18912 27402 18964
rect 30101 18955 30159 18961
rect 30101 18921 30113 18955
rect 30147 18921 30159 18955
rect 30101 18915 30159 18921
rect 3237 18887 3295 18893
rect 3237 18853 3249 18887
rect 3283 18884 3295 18887
rect 3283 18856 4292 18884
rect 3283 18853 3295 18856
rect 3237 18847 3295 18853
rect 4264 18825 4292 18856
rect 6730 18844 6736 18896
rect 6788 18884 6794 18896
rect 6788 18856 7512 18884
rect 6788 18844 6794 18856
rect 4249 18819 4307 18825
rect 4249 18785 4261 18819
rect 4295 18785 4307 18819
rect 4249 18779 4307 18785
rect 4433 18819 4491 18825
rect 4433 18785 4445 18819
rect 4479 18816 4491 18819
rect 4614 18816 4620 18828
rect 4479 18788 4620 18816
rect 4479 18785 4491 18788
rect 4433 18779 4491 18785
rect 1854 18748 1860 18760
rect 1815 18720 1860 18748
rect 1854 18708 1860 18720
rect 1912 18708 1918 18760
rect 2130 18757 2136 18760
rect 2124 18748 2136 18757
rect 2091 18720 2136 18748
rect 2124 18711 2136 18720
rect 2130 18708 2136 18711
rect 2188 18708 2194 18760
rect 4264 18748 4292 18779
rect 4614 18776 4620 18788
rect 4672 18776 4678 18828
rect 7374 18816 7380 18828
rect 6932 18788 7380 18816
rect 6932 18760 6960 18788
rect 7374 18776 7380 18788
rect 7432 18776 7438 18828
rect 5353 18751 5411 18757
rect 5353 18748 5365 18751
rect 4264 18720 5365 18748
rect 5353 18717 5365 18720
rect 5399 18717 5411 18751
rect 5353 18711 5411 18717
rect 5445 18751 5503 18757
rect 5445 18717 5457 18751
rect 5491 18748 5503 18751
rect 5534 18748 5540 18760
rect 5491 18720 5540 18748
rect 5491 18717 5503 18720
rect 5445 18711 5503 18717
rect 5534 18708 5540 18720
rect 5592 18708 5598 18760
rect 6914 18748 6920 18760
rect 6875 18720 6920 18748
rect 6914 18708 6920 18720
rect 6972 18708 6978 18760
rect 7006 18708 7012 18760
rect 7064 18748 7070 18760
rect 7101 18751 7159 18757
rect 7101 18748 7113 18751
rect 7064 18720 7113 18748
rect 7064 18708 7070 18720
rect 7101 18717 7113 18720
rect 7147 18717 7159 18751
rect 7101 18711 7159 18717
rect 7193 18751 7251 18757
rect 7193 18717 7205 18751
rect 7239 18717 7251 18751
rect 7193 18711 7251 18717
rect 4062 18640 4068 18692
rect 4120 18680 4126 18692
rect 4890 18680 4896 18692
rect 4120 18652 4896 18680
rect 4120 18640 4126 18652
rect 4890 18640 4896 18652
rect 4948 18640 4954 18692
rect 6273 18683 6331 18689
rect 6273 18649 6285 18683
rect 6319 18649 6331 18683
rect 6273 18643 6331 18649
rect 3326 18572 3332 18624
rect 3384 18612 3390 18624
rect 3789 18615 3847 18621
rect 3789 18612 3801 18615
rect 3384 18584 3801 18612
rect 3384 18572 3390 18584
rect 3789 18581 3801 18584
rect 3835 18581 3847 18615
rect 4154 18612 4160 18624
rect 4115 18584 4160 18612
rect 3789 18575 3847 18581
rect 4154 18572 4160 18584
rect 4212 18572 4218 18624
rect 4985 18615 5043 18621
rect 4985 18581 4997 18615
rect 5031 18612 5043 18615
rect 5626 18612 5632 18624
rect 5031 18584 5632 18612
rect 5031 18581 5043 18584
rect 4985 18575 5043 18581
rect 5626 18572 5632 18584
rect 5684 18572 5690 18624
rect 6288 18612 6316 18643
rect 7208 18624 7236 18711
rect 7282 18708 7288 18760
rect 7340 18748 7346 18760
rect 7484 18757 7512 18856
rect 10870 18844 10876 18896
rect 10928 18884 10934 18896
rect 10928 18856 12020 18884
rect 10928 18844 10934 18856
rect 11425 18819 11483 18825
rect 11425 18816 11437 18819
rect 11164 18788 11437 18816
rect 7469 18751 7527 18757
rect 7340 18720 7385 18748
rect 7340 18708 7346 18720
rect 7469 18717 7481 18751
rect 7515 18748 7527 18751
rect 8113 18751 8171 18757
rect 8113 18748 8125 18751
rect 7515 18720 8125 18748
rect 7515 18717 7527 18720
rect 7469 18711 7527 18717
rect 8113 18717 8125 18720
rect 8159 18717 8171 18751
rect 9582 18748 9588 18760
rect 9543 18720 9588 18748
rect 8113 18711 8171 18717
rect 9582 18708 9588 18720
rect 9640 18708 9646 18760
rect 9852 18751 9910 18757
rect 9852 18717 9864 18751
rect 9898 18748 9910 18751
rect 11164 18748 11192 18788
rect 11425 18785 11437 18788
rect 11471 18785 11483 18819
rect 11425 18779 11483 18785
rect 11606 18776 11612 18828
rect 11664 18816 11670 18828
rect 11992 18816 12020 18856
rect 23014 18844 23020 18896
rect 23072 18884 23078 18896
rect 27614 18884 27620 18896
rect 23072 18856 27620 18884
rect 23072 18844 23078 18856
rect 27614 18844 27620 18856
rect 27672 18844 27678 18896
rect 30116 18884 30144 18915
rect 30466 18912 30472 18964
rect 30524 18952 30530 18964
rect 30745 18955 30803 18961
rect 30745 18952 30757 18955
rect 30524 18924 30757 18952
rect 30524 18912 30530 18924
rect 30745 18921 30757 18924
rect 30791 18921 30803 18955
rect 32769 18955 32827 18961
rect 30745 18915 30803 18921
rect 32140 18924 32720 18952
rect 30926 18884 30932 18896
rect 30116 18856 30932 18884
rect 30926 18844 30932 18856
rect 30984 18844 30990 18896
rect 11664 18788 11836 18816
rect 11992 18788 12112 18816
rect 11664 18776 11670 18788
rect 11698 18748 11704 18760
rect 9898 18720 11192 18748
rect 11659 18720 11704 18748
rect 9898 18717 9910 18720
rect 9852 18711 9910 18717
rect 11698 18708 11704 18720
rect 11756 18708 11762 18760
rect 11808 18757 11836 18788
rect 11793 18751 11851 18757
rect 11793 18717 11805 18751
rect 11839 18717 11851 18751
rect 11793 18711 11851 18717
rect 11882 18708 11888 18760
rect 11940 18748 11946 18760
rect 12084 18757 12112 18788
rect 13722 18776 13728 18828
rect 13780 18816 13786 18828
rect 17589 18819 17647 18825
rect 17589 18816 17601 18819
rect 13780 18788 17601 18816
rect 13780 18776 13786 18788
rect 17589 18785 17601 18788
rect 17635 18816 17647 18819
rect 17635 18788 18460 18816
rect 17635 18785 17647 18788
rect 17589 18779 17647 18785
rect 12069 18751 12127 18757
rect 11940 18720 11985 18748
rect 11940 18708 11946 18720
rect 12069 18717 12081 18751
rect 12115 18717 12127 18751
rect 12069 18711 12127 18717
rect 15838 18708 15844 18760
rect 15896 18748 15902 18760
rect 16669 18751 16727 18757
rect 16669 18748 16681 18751
rect 15896 18720 16681 18748
rect 15896 18708 15902 18720
rect 16669 18717 16681 18720
rect 16715 18717 16727 18751
rect 16669 18711 16727 18717
rect 16761 18751 16819 18757
rect 16761 18717 16773 18751
rect 16807 18717 16819 18751
rect 16761 18711 16819 18717
rect 10594 18640 10600 18692
rect 10652 18680 10658 18692
rect 12529 18683 12587 18689
rect 12529 18680 12541 18683
rect 10652 18652 12541 18680
rect 10652 18640 10658 18652
rect 12529 18649 12541 18652
rect 12575 18649 12587 18683
rect 16776 18680 16804 18711
rect 16850 18708 16856 18760
rect 16908 18748 16914 18760
rect 17037 18751 17095 18757
rect 16908 18720 16953 18748
rect 16908 18708 16914 18720
rect 17037 18717 17049 18751
rect 17083 18748 17095 18751
rect 17310 18748 17316 18760
rect 17083 18720 17316 18748
rect 17083 18717 17095 18720
rect 17037 18711 17095 18717
rect 17310 18708 17316 18720
rect 17368 18748 17374 18760
rect 18049 18751 18107 18757
rect 18049 18748 18061 18751
rect 17368 18720 18061 18748
rect 17368 18708 17374 18720
rect 18049 18717 18061 18720
rect 18095 18717 18107 18751
rect 18230 18748 18236 18760
rect 18191 18720 18236 18748
rect 18049 18711 18107 18717
rect 18230 18708 18236 18720
rect 18288 18708 18294 18760
rect 18432 18757 18460 18788
rect 18524 18788 19380 18816
rect 18325 18751 18383 18757
rect 18325 18717 18337 18751
rect 18371 18717 18383 18751
rect 18325 18711 18383 18717
rect 18417 18751 18475 18757
rect 18417 18717 18429 18751
rect 18463 18717 18475 18751
rect 18417 18711 18475 18717
rect 17126 18680 17132 18692
rect 16776 18652 17132 18680
rect 12529 18643 12587 18649
rect 17126 18640 17132 18652
rect 17184 18680 17190 18692
rect 18340 18680 18368 18711
rect 18524 18680 18552 18788
rect 18690 18708 18696 18760
rect 18748 18748 18754 18760
rect 19245 18751 19303 18757
rect 19245 18748 19257 18751
rect 18748 18720 19257 18748
rect 18748 18708 18754 18720
rect 19245 18717 19257 18720
rect 19291 18717 19303 18751
rect 19352 18748 19380 18788
rect 20898 18776 20904 18828
rect 20956 18816 20962 18828
rect 21910 18816 21916 18828
rect 20956 18788 21772 18816
rect 21871 18788 21916 18816
rect 20956 18776 20962 18788
rect 21637 18751 21695 18757
rect 21637 18748 21649 18751
rect 19352 18720 21649 18748
rect 19245 18711 19303 18717
rect 21637 18717 21649 18720
rect 21683 18717 21695 18751
rect 21744 18748 21772 18788
rect 21910 18776 21916 18788
rect 21968 18776 21974 18828
rect 23293 18819 23351 18825
rect 23293 18785 23305 18819
rect 23339 18816 23351 18819
rect 23382 18816 23388 18828
rect 23339 18788 23388 18816
rect 23339 18785 23351 18788
rect 23293 18779 23351 18785
rect 23382 18776 23388 18788
rect 23440 18776 23446 18828
rect 30374 18816 30380 18828
rect 29840 18788 30380 18816
rect 29840 18757 29868 18788
rect 30374 18776 30380 18788
rect 30432 18776 30438 18828
rect 32140 18816 32168 18924
rect 32490 18884 32496 18896
rect 30760 18788 32168 18816
rect 32232 18856 32496 18884
rect 23017 18751 23075 18757
rect 23017 18748 23029 18751
rect 21744 18720 23029 18748
rect 21637 18711 21695 18717
rect 23017 18717 23029 18720
rect 23063 18717 23075 18751
rect 23017 18711 23075 18717
rect 29825 18751 29883 18757
rect 29825 18717 29837 18751
rect 29871 18717 29883 18751
rect 29825 18711 29883 18717
rect 29917 18751 29975 18757
rect 29917 18717 29929 18751
rect 29963 18717 29975 18751
rect 30098 18748 30104 18760
rect 30059 18720 30104 18748
rect 29917 18711 29975 18717
rect 19490 18683 19548 18689
rect 19490 18680 19502 18683
rect 17184 18652 18552 18680
rect 18708 18652 19502 18680
rect 17184 18640 17190 18652
rect 6914 18612 6920 18624
rect 6288 18584 6920 18612
rect 6914 18572 6920 18584
rect 6972 18572 6978 18624
rect 7190 18572 7196 18624
rect 7248 18572 7254 18624
rect 7650 18612 7656 18624
rect 7611 18584 7656 18612
rect 7650 18572 7656 18584
rect 7708 18572 7714 18624
rect 10965 18615 11023 18621
rect 10965 18581 10977 18615
rect 11011 18612 11023 18615
rect 11054 18612 11060 18624
rect 11011 18584 11060 18612
rect 11011 18581 11023 18584
rect 10965 18575 11023 18581
rect 11054 18572 11060 18584
rect 11112 18572 11118 18624
rect 18708 18621 18736 18652
rect 19490 18649 19502 18652
rect 19536 18649 19548 18683
rect 19490 18643 19548 18649
rect 20806 18640 20812 18692
rect 20864 18680 20870 18692
rect 26786 18680 26792 18692
rect 20864 18652 26792 18680
rect 20864 18640 20870 18652
rect 26786 18640 26792 18652
rect 26844 18640 26850 18692
rect 27341 18683 27399 18689
rect 27341 18649 27353 18683
rect 27387 18649 27399 18683
rect 27341 18643 27399 18649
rect 18693 18615 18751 18621
rect 18693 18581 18705 18615
rect 18739 18581 18751 18615
rect 18693 18575 18751 18581
rect 25498 18572 25504 18624
rect 25556 18612 25562 18624
rect 26510 18612 26516 18624
rect 25556 18584 26516 18612
rect 25556 18572 25562 18584
rect 26510 18572 26516 18584
rect 26568 18612 26574 18624
rect 26697 18615 26755 18621
rect 26697 18612 26709 18615
rect 26568 18584 26709 18612
rect 26568 18572 26574 18584
rect 26697 18581 26709 18584
rect 26743 18612 26755 18615
rect 27356 18612 27384 18643
rect 27982 18640 27988 18692
rect 28040 18680 28046 18692
rect 29932 18680 29960 18711
rect 30098 18708 30104 18720
rect 30156 18708 30162 18760
rect 30558 18708 30564 18760
rect 30616 18708 30622 18760
rect 30760 18757 30788 18788
rect 30745 18751 30803 18757
rect 30745 18717 30757 18751
rect 30791 18717 30803 18751
rect 30745 18711 30803 18717
rect 30837 18751 30895 18757
rect 30837 18717 30849 18751
rect 30883 18748 30895 18751
rect 30926 18748 30932 18760
rect 30883 18720 30932 18748
rect 30883 18717 30895 18720
rect 30837 18711 30895 18717
rect 30926 18708 30932 18720
rect 30984 18708 30990 18760
rect 31938 18708 31944 18760
rect 31996 18748 32002 18760
rect 32113 18751 32171 18757
rect 32113 18748 32125 18751
rect 31996 18720 32125 18748
rect 31996 18708 32002 18720
rect 32113 18717 32125 18720
rect 32159 18717 32171 18751
rect 32232 18748 32260 18856
rect 32490 18844 32496 18856
rect 32548 18844 32554 18896
rect 32692 18884 32720 18924
rect 32769 18921 32781 18955
rect 32815 18952 32827 18955
rect 33318 18952 33324 18964
rect 32815 18924 33324 18952
rect 32815 18921 32827 18924
rect 32769 18915 32827 18921
rect 33318 18912 33324 18924
rect 33376 18912 33382 18964
rect 34422 18912 34428 18964
rect 34480 18952 34486 18964
rect 37277 18955 37335 18961
rect 37277 18952 37289 18955
rect 34480 18924 37289 18952
rect 34480 18912 34486 18924
rect 37277 18921 37289 18924
rect 37323 18921 37335 18955
rect 37277 18915 37335 18921
rect 40221 18955 40279 18961
rect 40221 18921 40233 18955
rect 40267 18952 40279 18955
rect 41046 18952 41052 18964
rect 40267 18924 41052 18952
rect 40267 18921 40279 18924
rect 40221 18915 40279 18921
rect 41046 18912 41052 18924
rect 41104 18912 41110 18964
rect 34514 18884 34520 18896
rect 32692 18856 34520 18884
rect 34514 18844 34520 18856
rect 34572 18844 34578 18896
rect 32674 18816 32680 18828
rect 32416 18788 32680 18816
rect 32416 18757 32444 18788
rect 32674 18776 32680 18788
rect 32732 18776 32738 18828
rect 37918 18816 37924 18828
rect 37568 18788 37924 18816
rect 32288 18751 32346 18757
rect 32288 18748 32300 18751
rect 32232 18720 32300 18748
rect 32113 18711 32171 18717
rect 32288 18717 32300 18720
rect 32334 18717 32346 18751
rect 32288 18711 32346 18717
rect 32404 18751 32462 18757
rect 32404 18717 32416 18751
rect 32450 18717 32462 18751
rect 32404 18711 32462 18717
rect 32493 18751 32551 18757
rect 32493 18717 32505 18751
rect 32539 18717 32551 18751
rect 32493 18711 32551 18717
rect 28040 18652 29960 18680
rect 30576 18680 30604 18708
rect 31021 18683 31079 18689
rect 31021 18680 31033 18683
rect 30576 18652 31033 18680
rect 28040 18640 28046 18652
rect 31021 18649 31033 18652
rect 31067 18649 31079 18683
rect 31021 18643 31079 18649
rect 26743 18584 27384 18612
rect 26743 18581 26755 18584
rect 26697 18575 26755 18581
rect 27430 18572 27436 18624
rect 27488 18612 27494 18624
rect 28810 18612 28816 18624
rect 27488 18584 28816 18612
rect 27488 18572 27494 18584
rect 28810 18572 28816 18584
rect 28868 18572 28874 18624
rect 29638 18612 29644 18624
rect 29599 18584 29644 18612
rect 29638 18572 29644 18584
rect 29696 18572 29702 18624
rect 30558 18612 30564 18624
rect 30519 18584 30564 18612
rect 30558 18572 30564 18584
rect 30616 18572 30622 18624
rect 31662 18612 31668 18624
rect 31575 18584 31668 18612
rect 31662 18572 31668 18584
rect 31720 18612 31726 18624
rect 32508 18612 32536 18711
rect 36998 18708 37004 18760
rect 37056 18748 37062 18760
rect 37568 18757 37596 18788
rect 37918 18776 37924 18788
rect 37976 18816 37982 18828
rect 37976 18788 40080 18816
rect 37976 18776 37982 18788
rect 37461 18751 37519 18757
rect 37461 18748 37473 18751
rect 37056 18720 37473 18748
rect 37056 18708 37062 18720
rect 37461 18717 37473 18720
rect 37507 18717 37519 18751
rect 37461 18711 37519 18717
rect 37553 18751 37611 18757
rect 37553 18717 37565 18751
rect 37599 18717 37611 18751
rect 37553 18711 37611 18717
rect 37829 18751 37887 18757
rect 37829 18717 37841 18751
rect 37875 18748 37887 18751
rect 38930 18748 38936 18760
rect 37875 18720 38936 18748
rect 37875 18717 37887 18720
rect 37829 18711 37887 18717
rect 38930 18708 38936 18720
rect 38988 18708 38994 18760
rect 40052 18757 40080 18788
rect 40037 18751 40095 18757
rect 40037 18717 40049 18751
rect 40083 18717 40095 18751
rect 58158 18748 58164 18760
rect 58119 18720 58164 18748
rect 40037 18711 40095 18717
rect 58158 18708 58164 18720
rect 58216 18708 58222 18760
rect 37182 18640 37188 18692
rect 37240 18680 37246 18692
rect 37645 18683 37703 18689
rect 37645 18680 37657 18683
rect 37240 18652 37657 18680
rect 37240 18640 37246 18652
rect 37645 18649 37657 18652
rect 37691 18649 37703 18683
rect 37645 18643 37703 18649
rect 38746 18640 38752 18692
rect 38804 18680 38810 18692
rect 39850 18680 39856 18692
rect 38804 18652 39856 18680
rect 38804 18640 38810 18652
rect 39850 18640 39856 18652
rect 39908 18640 39914 18692
rect 40681 18615 40739 18621
rect 40681 18612 40693 18615
rect 31720 18584 40693 18612
rect 31720 18572 31726 18584
rect 40681 18581 40693 18584
rect 40727 18612 40739 18615
rect 40862 18612 40868 18624
rect 40727 18584 40868 18612
rect 40727 18581 40739 18584
rect 40681 18575 40739 18581
rect 40862 18572 40868 18584
rect 40920 18612 40926 18624
rect 41046 18612 41052 18624
rect 40920 18584 41052 18612
rect 40920 18572 40926 18584
rect 41046 18572 41052 18584
rect 41104 18572 41110 18624
rect 41322 18572 41328 18624
rect 41380 18612 41386 18624
rect 41509 18615 41567 18621
rect 41509 18612 41521 18615
rect 41380 18584 41521 18612
rect 41380 18572 41386 18584
rect 41509 18581 41521 18584
rect 41555 18581 41567 18615
rect 41509 18575 41567 18581
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 2317 18411 2375 18417
rect 2317 18377 2329 18411
rect 2363 18408 2375 18411
rect 2406 18408 2412 18420
rect 2363 18380 2412 18408
rect 2363 18377 2375 18380
rect 2317 18371 2375 18377
rect 2406 18368 2412 18380
rect 2464 18368 2470 18420
rect 5169 18411 5227 18417
rect 5169 18377 5181 18411
rect 5215 18408 5227 18411
rect 7190 18408 7196 18420
rect 5215 18380 7196 18408
rect 5215 18377 5227 18380
rect 5169 18371 5227 18377
rect 7190 18368 7196 18380
rect 7248 18368 7254 18420
rect 8294 18408 8300 18420
rect 7300 18380 8300 18408
rect 3697 18343 3755 18349
rect 3697 18309 3709 18343
rect 3743 18340 3755 18343
rect 4062 18340 4068 18352
rect 3743 18312 4068 18340
rect 3743 18309 3755 18312
rect 3697 18303 3755 18309
rect 4062 18300 4068 18312
rect 4120 18300 4126 18352
rect 4525 18343 4583 18349
rect 4525 18309 4537 18343
rect 4571 18340 4583 18343
rect 5626 18340 5632 18352
rect 4571 18312 5632 18340
rect 4571 18309 4583 18312
rect 4525 18303 4583 18309
rect 5626 18300 5632 18312
rect 5684 18300 5690 18352
rect 7006 18300 7012 18352
rect 7064 18340 7070 18352
rect 7300 18340 7328 18380
rect 8294 18368 8300 18380
rect 8352 18368 8358 18420
rect 11606 18408 11612 18420
rect 10704 18380 11612 18408
rect 7064 18312 7328 18340
rect 7064 18300 7070 18312
rect 7650 18300 7656 18352
rect 7708 18340 7714 18352
rect 7846 18343 7904 18349
rect 7846 18340 7858 18343
rect 7708 18312 7858 18340
rect 7708 18300 7714 18312
rect 7846 18309 7858 18312
rect 7892 18309 7904 18343
rect 7846 18303 7904 18309
rect 1670 18272 1676 18284
rect 1631 18244 1676 18272
rect 1670 18232 1676 18244
rect 1728 18232 1734 18284
rect 2501 18275 2559 18281
rect 2501 18241 2513 18275
rect 2547 18272 2559 18275
rect 3326 18272 3332 18284
rect 2547 18244 3332 18272
rect 2547 18241 2559 18244
rect 2501 18235 2559 18241
rect 3326 18232 3332 18244
rect 3384 18232 3390 18284
rect 4893 18275 4951 18281
rect 4893 18272 4905 18275
rect 3804 18244 4905 18272
rect 2406 18164 2412 18216
rect 2464 18204 2470 18216
rect 2685 18207 2743 18213
rect 2685 18204 2697 18207
rect 2464 18176 2697 18204
rect 2464 18164 2470 18176
rect 2685 18173 2697 18176
rect 2731 18173 2743 18207
rect 2685 18167 2743 18173
rect 3234 18164 3240 18216
rect 3292 18204 3298 18216
rect 3804 18213 3832 18244
rect 4893 18241 4905 18244
rect 4939 18241 4951 18275
rect 4893 18235 4951 18241
rect 7374 18232 7380 18284
rect 7432 18272 7438 18284
rect 8202 18272 8208 18284
rect 7432 18244 8208 18272
rect 7432 18232 7438 18244
rect 8202 18232 8208 18244
rect 8260 18232 8266 18284
rect 9214 18232 9220 18284
rect 9272 18272 9278 18284
rect 10704 18281 10732 18380
rect 11606 18368 11612 18380
rect 11664 18368 11670 18420
rect 11882 18408 11888 18420
rect 11843 18380 11888 18408
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 11974 18368 11980 18420
rect 12032 18408 12038 18420
rect 14921 18411 14979 18417
rect 14921 18408 14933 18411
rect 12032 18380 14933 18408
rect 12032 18368 12038 18380
rect 14921 18377 14933 18380
rect 14967 18377 14979 18411
rect 14921 18371 14979 18377
rect 16850 18368 16856 18420
rect 16908 18408 16914 18420
rect 17037 18411 17095 18417
rect 17037 18408 17049 18411
rect 16908 18380 17049 18408
rect 16908 18368 16914 18380
rect 17037 18377 17049 18380
rect 17083 18377 17095 18411
rect 17037 18371 17095 18377
rect 18230 18368 18236 18420
rect 18288 18408 18294 18420
rect 18969 18411 19027 18417
rect 18969 18408 18981 18411
rect 18288 18380 18981 18408
rect 18288 18368 18294 18380
rect 18969 18377 18981 18380
rect 19015 18377 19027 18411
rect 18969 18371 19027 18377
rect 19242 18368 19248 18420
rect 19300 18408 19306 18420
rect 29638 18408 29644 18420
rect 19300 18380 29644 18408
rect 19300 18368 19306 18380
rect 29638 18368 29644 18380
rect 29696 18368 29702 18420
rect 32490 18408 32496 18420
rect 32451 18380 32496 18408
rect 32490 18368 32496 18380
rect 32548 18368 32554 18420
rect 38013 18411 38071 18417
rect 38013 18377 38025 18411
rect 38059 18408 38071 18411
rect 40586 18408 40592 18420
rect 38059 18380 40592 18408
rect 38059 18377 38071 18380
rect 38013 18371 38071 18377
rect 40586 18368 40592 18380
rect 40644 18408 40650 18420
rect 40644 18380 41092 18408
rect 40644 18368 40650 18380
rect 11054 18300 11060 18352
rect 11112 18340 11118 18352
rect 11701 18343 11759 18349
rect 11701 18340 11713 18343
rect 11112 18312 11713 18340
rect 11112 18300 11118 18312
rect 11701 18309 11713 18312
rect 11747 18309 11759 18343
rect 11701 18303 11759 18309
rect 12710 18300 12716 18352
rect 12768 18340 12774 18352
rect 12768 18312 13492 18340
rect 12768 18300 12774 18312
rect 10597 18275 10655 18281
rect 10597 18272 10609 18275
rect 9272 18244 10609 18272
rect 9272 18232 9278 18244
rect 10597 18241 10609 18244
rect 10643 18241 10655 18275
rect 10597 18235 10655 18241
rect 10689 18275 10747 18281
rect 10689 18241 10701 18275
rect 10735 18241 10747 18275
rect 10689 18235 10747 18241
rect 10781 18275 10839 18281
rect 10781 18241 10793 18275
rect 10827 18241 10839 18275
rect 10781 18235 10839 18241
rect 3789 18207 3847 18213
rect 3789 18204 3801 18207
rect 3292 18176 3801 18204
rect 3292 18164 3298 18176
rect 3789 18173 3801 18176
rect 3835 18173 3847 18207
rect 3789 18167 3847 18173
rect 3973 18207 4031 18213
rect 3973 18173 3985 18207
rect 4019 18204 4031 18207
rect 4614 18204 4620 18216
rect 4019 18176 4620 18204
rect 4019 18173 4031 18176
rect 3973 18167 4031 18173
rect 4614 18164 4620 18176
rect 4672 18164 4678 18216
rect 4985 18207 5043 18213
rect 4985 18173 4997 18207
rect 5031 18204 5043 18207
rect 5534 18204 5540 18216
rect 5031 18176 5540 18204
rect 5031 18173 5043 18176
rect 4985 18167 5043 18173
rect 5534 18164 5540 18176
rect 5592 18204 5598 18216
rect 6086 18204 6092 18216
rect 5592 18176 6092 18204
rect 5592 18164 5598 18176
rect 6086 18164 6092 18176
rect 6144 18164 6150 18216
rect 8113 18207 8171 18213
rect 8113 18173 8125 18207
rect 8159 18204 8171 18207
rect 9582 18204 9588 18216
rect 8159 18176 9588 18204
rect 8159 18173 8171 18176
rect 8113 18167 8171 18173
rect 9582 18164 9588 18176
rect 9640 18164 9646 18216
rect 10796 18204 10824 18235
rect 10870 18232 10876 18284
rect 10928 18272 10934 18284
rect 10965 18275 11023 18281
rect 10965 18272 10977 18275
rect 10928 18244 10977 18272
rect 10928 18232 10934 18244
rect 10965 18241 10977 18244
rect 11011 18241 11023 18275
rect 10965 18235 11023 18241
rect 11517 18275 11575 18281
rect 11517 18241 11529 18275
rect 11563 18272 11575 18275
rect 12342 18272 12348 18284
rect 11563 18244 12348 18272
rect 11563 18241 11575 18244
rect 11517 18235 11575 18241
rect 12342 18232 12348 18244
rect 12400 18232 12406 18284
rect 12526 18232 12532 18284
rect 12584 18272 12590 18284
rect 12621 18275 12679 18281
rect 12621 18272 12633 18275
rect 12584 18244 12633 18272
rect 12584 18232 12590 18244
rect 12621 18241 12633 18244
rect 12667 18241 12679 18275
rect 13170 18272 13176 18284
rect 13131 18244 13176 18272
rect 12621 18235 12679 18241
rect 13170 18232 13176 18244
rect 13228 18232 13234 18284
rect 13464 18281 13492 18312
rect 13906 18300 13912 18352
rect 13964 18340 13970 18352
rect 30558 18340 30564 18352
rect 13964 18312 30564 18340
rect 13964 18300 13970 18312
rect 30558 18300 30564 18312
rect 30616 18300 30622 18352
rect 31938 18300 31944 18352
rect 31996 18340 32002 18352
rect 32125 18343 32183 18349
rect 32125 18340 32137 18343
rect 31996 18312 32137 18340
rect 31996 18300 32002 18312
rect 32125 18309 32137 18312
rect 32171 18340 32183 18343
rect 32766 18340 32772 18352
rect 32171 18312 32772 18340
rect 32171 18309 32183 18312
rect 32125 18303 32183 18309
rect 32766 18300 32772 18312
rect 32824 18340 32830 18352
rect 32953 18343 33011 18349
rect 32953 18340 32965 18343
rect 32824 18312 32965 18340
rect 32824 18300 32830 18312
rect 32953 18309 32965 18312
rect 32999 18309 33011 18343
rect 32953 18303 33011 18309
rect 33137 18343 33195 18349
rect 33137 18309 33149 18343
rect 33183 18340 33195 18343
rect 33410 18340 33416 18352
rect 33183 18312 33416 18340
rect 33183 18309 33195 18312
rect 33137 18303 33195 18309
rect 33410 18300 33416 18312
rect 33468 18340 33474 18352
rect 34422 18340 34428 18352
rect 33468 18312 34428 18340
rect 33468 18300 33474 18312
rect 34422 18300 34428 18312
rect 34480 18300 34486 18352
rect 36541 18343 36599 18349
rect 36541 18309 36553 18343
rect 36587 18340 36599 18343
rect 37182 18340 37188 18352
rect 36587 18312 37188 18340
rect 36587 18309 36599 18312
rect 36541 18303 36599 18309
rect 37182 18300 37188 18312
rect 37240 18300 37246 18352
rect 37550 18300 37556 18352
rect 37608 18340 37614 18352
rect 38105 18343 38163 18349
rect 38105 18340 38117 18343
rect 37608 18312 38117 18340
rect 37608 18300 37614 18312
rect 38105 18309 38117 18312
rect 38151 18309 38163 18343
rect 38105 18303 38163 18309
rect 39298 18300 39304 18352
rect 39356 18340 39362 18352
rect 41064 18340 41092 18380
rect 39356 18312 40356 18340
rect 41064 18312 41184 18340
rect 39356 18300 39362 18312
rect 13357 18275 13415 18281
rect 13357 18241 13369 18275
rect 13403 18241 13415 18275
rect 13357 18235 13415 18241
rect 13449 18275 13507 18281
rect 13449 18241 13461 18275
rect 13495 18241 13507 18275
rect 13449 18235 13507 18241
rect 13541 18275 13599 18281
rect 13541 18241 13553 18275
rect 13587 18272 13599 18275
rect 13630 18272 13636 18284
rect 13587 18244 13636 18272
rect 13587 18241 13599 18244
rect 13541 18235 13599 18241
rect 11422 18204 11428 18216
rect 10796 18176 11428 18204
rect 11422 18164 11428 18176
rect 11480 18164 11486 18216
rect 13372 18204 13400 18235
rect 13630 18232 13636 18244
rect 13688 18232 13694 18284
rect 14274 18272 14280 18284
rect 14235 18244 14280 18272
rect 14274 18232 14280 18244
rect 14332 18232 14338 18284
rect 14366 18232 14372 18284
rect 14424 18272 14430 18284
rect 14550 18272 14556 18284
rect 14424 18244 14469 18272
rect 14511 18244 14556 18272
rect 14424 18232 14430 18244
rect 14550 18232 14556 18244
rect 14608 18232 14614 18284
rect 14645 18275 14703 18281
rect 14645 18241 14657 18275
rect 14691 18241 14703 18275
rect 14645 18235 14703 18241
rect 14660 18204 14688 18235
rect 14734 18232 14740 18284
rect 14792 18281 14798 18284
rect 14792 18272 14800 18281
rect 17221 18275 17279 18281
rect 14792 18244 14837 18272
rect 14792 18235 14800 18244
rect 17221 18241 17233 18275
rect 17267 18241 17279 18275
rect 17221 18235 17279 18241
rect 17405 18275 17463 18281
rect 17405 18241 17417 18275
rect 17451 18272 17463 18275
rect 17954 18272 17960 18284
rect 17451 18244 17960 18272
rect 17451 18241 17463 18244
rect 17405 18235 17463 18241
rect 14792 18232 14798 18235
rect 16942 18204 16948 18216
rect 13372 18176 13492 18204
rect 14660 18176 16948 18204
rect 5810 18136 5816 18148
rect 5723 18108 5816 18136
rect 5810 18096 5816 18108
rect 5868 18136 5874 18148
rect 9861 18139 9919 18145
rect 5868 18108 6868 18136
rect 5868 18096 5874 18108
rect 1857 18071 1915 18077
rect 1857 18037 1869 18071
rect 1903 18068 1915 18071
rect 1946 18068 1952 18080
rect 1903 18040 1952 18068
rect 1903 18037 1915 18040
rect 1857 18031 1915 18037
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 3326 18068 3332 18080
rect 3287 18040 3332 18068
rect 3326 18028 3332 18040
rect 3384 18028 3390 18080
rect 6730 18068 6736 18080
rect 6691 18040 6736 18068
rect 6730 18028 6736 18040
rect 6788 18028 6794 18080
rect 6840 18068 6868 18108
rect 9861 18105 9873 18139
rect 9907 18136 9919 18139
rect 10870 18136 10876 18148
rect 9907 18108 10876 18136
rect 9907 18105 9919 18108
rect 9861 18099 9919 18105
rect 10870 18096 10876 18108
rect 10928 18096 10934 18148
rect 13464 18136 13492 18176
rect 16942 18164 16948 18176
rect 17000 18164 17006 18216
rect 17236 18204 17264 18235
rect 17954 18232 17960 18244
rect 18012 18272 18018 18284
rect 19153 18275 19211 18281
rect 18012 18244 18215 18272
rect 18012 18232 18018 18244
rect 18046 18204 18052 18216
rect 17236 18176 18052 18204
rect 18046 18164 18052 18176
rect 18104 18164 18110 18216
rect 13906 18136 13912 18148
rect 13464 18108 13912 18136
rect 13906 18096 13912 18108
rect 13964 18096 13970 18148
rect 18187 18136 18215 18244
rect 19153 18241 19165 18275
rect 19199 18241 19211 18275
rect 19153 18235 19211 18241
rect 19169 18204 19197 18235
rect 19242 18232 19248 18284
rect 19300 18272 19306 18284
rect 19337 18275 19395 18281
rect 19337 18272 19349 18275
rect 19300 18244 19349 18272
rect 19300 18232 19306 18244
rect 19337 18241 19349 18244
rect 19383 18272 19395 18275
rect 21177 18275 21235 18281
rect 19383 18244 21036 18272
rect 19383 18241 19395 18244
rect 19337 18235 19395 18241
rect 20622 18204 20628 18216
rect 19169 18176 20628 18204
rect 20622 18164 20628 18176
rect 20680 18164 20686 18216
rect 19242 18136 19248 18148
rect 18187 18108 19248 18136
rect 19242 18096 19248 18108
rect 19300 18096 19306 18148
rect 21008 18145 21036 18244
rect 21177 18241 21189 18275
rect 21223 18272 21235 18275
rect 22005 18275 22063 18281
rect 21223 18244 21864 18272
rect 21223 18241 21235 18244
rect 21177 18235 21235 18241
rect 21836 18145 21864 18244
rect 22005 18241 22017 18275
rect 22051 18272 22063 18275
rect 22094 18272 22100 18284
rect 22051 18244 22100 18272
rect 22051 18241 22063 18244
rect 22005 18235 22063 18241
rect 22094 18232 22100 18244
rect 22152 18232 22158 18284
rect 23382 18272 23388 18284
rect 23343 18244 23388 18272
rect 23382 18232 23388 18244
rect 23440 18232 23446 18284
rect 24486 18272 24492 18284
rect 24447 18244 24492 18272
rect 24486 18232 24492 18244
rect 24544 18232 24550 18284
rect 24670 18272 24676 18284
rect 24583 18244 24676 18272
rect 24670 18232 24676 18244
rect 24728 18232 24734 18284
rect 24765 18275 24823 18281
rect 24765 18241 24777 18275
rect 24811 18241 24823 18275
rect 24765 18235 24823 18241
rect 24857 18275 24915 18281
rect 24857 18241 24869 18275
rect 24903 18272 24915 18275
rect 24946 18272 24952 18284
rect 24903 18244 24952 18272
rect 24903 18241 24915 18244
rect 24857 18235 24915 18241
rect 21910 18164 21916 18216
rect 21968 18204 21974 18216
rect 22189 18207 22247 18213
rect 22189 18204 22201 18207
rect 21968 18176 22201 18204
rect 21968 18164 21974 18176
rect 22189 18173 22201 18176
rect 22235 18204 22247 18207
rect 22649 18207 22707 18213
rect 22649 18204 22661 18207
rect 22235 18176 22661 18204
rect 22235 18173 22247 18176
rect 22189 18167 22247 18173
rect 22649 18173 22661 18176
rect 22695 18173 22707 18207
rect 22649 18167 22707 18173
rect 24394 18164 24400 18216
rect 24452 18204 24458 18216
rect 24688 18204 24716 18232
rect 24452 18176 24716 18204
rect 24780 18204 24808 18235
rect 24946 18232 24952 18244
rect 25004 18232 25010 18284
rect 25774 18232 25780 18284
rect 25832 18272 25838 18284
rect 26970 18272 26976 18284
rect 25832 18244 26976 18272
rect 25832 18232 25838 18244
rect 26970 18232 26976 18244
rect 27028 18232 27034 18284
rect 29089 18275 29147 18281
rect 29089 18241 29101 18275
rect 29135 18272 29147 18275
rect 29270 18272 29276 18284
rect 29135 18244 29276 18272
rect 29135 18241 29147 18244
rect 29089 18235 29147 18241
rect 29270 18232 29276 18244
rect 29328 18272 29334 18284
rect 29641 18275 29699 18281
rect 29641 18272 29653 18275
rect 29328 18244 29653 18272
rect 29328 18232 29334 18244
rect 29641 18241 29653 18244
rect 29687 18241 29699 18275
rect 29641 18235 29699 18241
rect 32214 18232 32220 18284
rect 32272 18272 32278 18284
rect 32309 18275 32367 18281
rect 32309 18272 32321 18275
rect 32272 18244 32321 18272
rect 32272 18232 32278 18244
rect 32309 18241 32321 18244
rect 32355 18241 32367 18275
rect 32309 18235 32367 18241
rect 36357 18275 36415 18281
rect 36357 18241 36369 18275
rect 36403 18241 36415 18275
rect 36357 18235 36415 18241
rect 26234 18204 26240 18216
rect 24780 18176 26240 18204
rect 24452 18164 24458 18176
rect 26234 18164 26240 18176
rect 26292 18164 26298 18216
rect 28810 18164 28816 18216
rect 28868 18204 28874 18216
rect 31662 18204 31668 18216
rect 28868 18176 31668 18204
rect 28868 18164 28874 18176
rect 31662 18164 31668 18176
rect 31720 18164 31726 18216
rect 36372 18204 36400 18235
rect 36446 18232 36452 18284
rect 36504 18272 36510 18284
rect 36725 18275 36783 18281
rect 36504 18244 36549 18272
rect 36504 18232 36510 18244
rect 36725 18241 36737 18275
rect 36771 18272 36783 18275
rect 37458 18272 37464 18284
rect 36771 18244 37464 18272
rect 36771 18241 36783 18244
rect 36725 18235 36783 18241
rect 37458 18232 37464 18244
rect 37516 18232 37522 18284
rect 40328 18281 40356 18312
rect 40057 18275 40115 18281
rect 40057 18241 40069 18275
rect 40103 18272 40115 18275
rect 40313 18275 40371 18281
rect 40103 18244 40264 18272
rect 40103 18241 40115 18244
rect 40057 18235 40115 18241
rect 36998 18204 37004 18216
rect 36372 18176 37004 18204
rect 36998 18164 37004 18176
rect 37056 18164 37062 18216
rect 40236 18204 40264 18244
rect 40313 18241 40325 18275
rect 40359 18241 40371 18275
rect 41046 18272 41052 18284
rect 41007 18244 41052 18272
rect 40313 18235 40371 18241
rect 41046 18232 41052 18244
rect 41104 18232 41110 18284
rect 41156 18281 41184 18312
rect 41141 18275 41199 18281
rect 41141 18241 41153 18275
rect 41187 18241 41199 18275
rect 41141 18235 41199 18241
rect 41230 18232 41236 18284
rect 41288 18272 41294 18284
rect 41417 18275 41475 18281
rect 41288 18244 41333 18272
rect 41288 18232 41294 18244
rect 41417 18241 41429 18275
rect 41463 18241 41475 18275
rect 41417 18235 41475 18241
rect 40773 18207 40831 18213
rect 40773 18204 40785 18207
rect 40236 18176 40785 18204
rect 40773 18173 40785 18176
rect 40819 18173 40831 18207
rect 40773 18167 40831 18173
rect 41322 18164 41328 18216
rect 41380 18204 41386 18216
rect 41432 18204 41460 18235
rect 41380 18176 41460 18204
rect 41380 18164 41386 18176
rect 20993 18139 21051 18145
rect 20993 18105 21005 18139
rect 21039 18105 21051 18139
rect 20993 18099 21051 18105
rect 21821 18139 21879 18145
rect 21821 18105 21833 18139
rect 21867 18136 21879 18139
rect 23658 18136 23664 18148
rect 21867 18108 22140 18136
rect 21867 18105 21879 18108
rect 21821 18099 21879 18105
rect 6914 18068 6920 18080
rect 6840 18040 6920 18068
rect 6914 18028 6920 18040
rect 6972 18068 6978 18080
rect 7742 18068 7748 18080
rect 6972 18040 7748 18068
rect 6972 18028 6978 18040
rect 7742 18028 7748 18040
rect 7800 18028 7806 18080
rect 9214 18068 9220 18080
rect 9175 18040 9220 18068
rect 9214 18028 9220 18040
rect 9272 18028 9278 18080
rect 10318 18068 10324 18080
rect 10279 18040 10324 18068
rect 10318 18028 10324 18040
rect 10376 18028 10382 18080
rect 13814 18068 13820 18080
rect 13775 18040 13820 18068
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 14918 18028 14924 18080
rect 14976 18068 14982 18080
rect 21910 18068 21916 18080
rect 14976 18040 21916 18068
rect 14976 18028 14982 18040
rect 21910 18028 21916 18040
rect 21968 18028 21974 18080
rect 22112 18068 22140 18108
rect 22296 18108 23664 18136
rect 22296 18068 22324 18108
rect 23658 18096 23664 18108
rect 23716 18096 23722 18148
rect 27154 18096 27160 18148
rect 27212 18136 27218 18148
rect 36173 18139 36231 18145
rect 36173 18136 36185 18139
rect 27212 18108 36185 18136
rect 27212 18096 27218 18108
rect 36173 18105 36185 18108
rect 36219 18105 36231 18139
rect 36173 18099 36231 18105
rect 22112 18040 22324 18068
rect 23477 18071 23535 18077
rect 23477 18037 23489 18071
rect 23523 18068 23535 18071
rect 24854 18068 24860 18080
rect 23523 18040 24860 18068
rect 23523 18037 23535 18040
rect 23477 18031 23535 18037
rect 24854 18028 24860 18040
rect 24912 18028 24918 18080
rect 25038 18068 25044 18080
rect 24999 18040 25044 18068
rect 25038 18028 25044 18040
rect 25096 18028 25102 18080
rect 29730 18068 29736 18080
rect 29691 18040 29736 18068
rect 29730 18028 29736 18040
rect 29788 18068 29794 18080
rect 30006 18068 30012 18080
rect 29788 18040 30012 18068
rect 29788 18028 29794 18040
rect 30006 18028 30012 18040
rect 30064 18028 30070 18080
rect 32582 18028 32588 18080
rect 32640 18068 32646 18080
rect 33321 18071 33379 18077
rect 33321 18068 33333 18071
rect 32640 18040 33333 18068
rect 32640 18028 32646 18040
rect 33321 18037 33333 18040
rect 33367 18037 33379 18071
rect 38930 18068 38936 18080
rect 38891 18040 38936 18068
rect 33321 18031 33379 18037
rect 38930 18028 38936 18040
rect 38988 18028 38994 18080
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 1670 17824 1676 17876
rect 1728 17864 1734 17876
rect 2133 17867 2191 17873
rect 2133 17864 2145 17867
rect 1728 17836 2145 17864
rect 1728 17824 1734 17836
rect 2133 17833 2145 17836
rect 2179 17833 2191 17867
rect 2133 17827 2191 17833
rect 4062 17824 4068 17876
rect 4120 17864 4126 17876
rect 4157 17867 4215 17873
rect 4157 17864 4169 17867
rect 4120 17836 4169 17864
rect 4120 17824 4126 17836
rect 4157 17833 4169 17836
rect 4203 17864 4215 17867
rect 5810 17864 5816 17876
rect 4203 17836 5816 17864
rect 4203 17833 4215 17836
rect 4157 17827 4215 17833
rect 5810 17824 5816 17836
rect 5868 17824 5874 17876
rect 6178 17824 6184 17876
rect 6236 17864 6242 17876
rect 6733 17867 6791 17873
rect 6733 17864 6745 17867
rect 6236 17836 6745 17864
rect 6236 17824 6242 17836
rect 6733 17833 6745 17836
rect 6779 17864 6791 17867
rect 9858 17864 9864 17876
rect 6779 17836 9864 17864
rect 6779 17833 6791 17836
rect 6733 17827 6791 17833
rect 9858 17824 9864 17836
rect 9916 17824 9922 17876
rect 12710 17824 12716 17876
rect 12768 17864 12774 17876
rect 19705 17867 19763 17873
rect 12768 17836 13124 17864
rect 12768 17824 12774 17836
rect 4890 17796 4896 17808
rect 4851 17768 4896 17796
rect 4890 17756 4896 17768
rect 4948 17756 4954 17808
rect 5074 17756 5080 17808
rect 5132 17796 5138 17808
rect 5721 17799 5779 17805
rect 5721 17796 5733 17799
rect 5132 17768 5733 17796
rect 5132 17756 5138 17768
rect 5721 17765 5733 17768
rect 5767 17796 5779 17799
rect 9214 17796 9220 17808
rect 5767 17768 9220 17796
rect 5767 17765 5779 17768
rect 5721 17759 5779 17765
rect 9214 17756 9220 17768
rect 9272 17796 9278 17808
rect 12986 17796 12992 17808
rect 9272 17768 12992 17796
rect 9272 17756 9278 17768
rect 12986 17756 12992 17768
rect 13044 17756 13050 17808
rect 13096 17796 13124 17836
rect 19705 17833 19717 17867
rect 19751 17833 19763 17867
rect 24854 17864 24860 17876
rect 19705 17827 19763 17833
rect 20916 17836 24860 17864
rect 13096 17768 13170 17796
rect 3326 17728 3332 17740
rect 2332 17700 3332 17728
rect 2332 17669 2360 17700
rect 3326 17688 3332 17700
rect 3384 17688 3390 17740
rect 2317 17663 2375 17669
rect 2317 17629 2329 17663
rect 2363 17629 2375 17663
rect 2317 17623 2375 17629
rect 2406 17620 2412 17672
rect 2464 17660 2470 17672
rect 3237 17663 3295 17669
rect 2464 17632 2509 17660
rect 2464 17620 2470 17632
rect 3237 17629 3249 17663
rect 3283 17660 3295 17663
rect 4706 17660 4712 17672
rect 3283 17632 4712 17660
rect 3283 17629 3295 17632
rect 3237 17623 3295 17629
rect 4706 17620 4712 17632
rect 4764 17620 4770 17672
rect 5166 17620 5172 17672
rect 5224 17660 5230 17672
rect 5537 17663 5595 17669
rect 5537 17660 5549 17663
rect 5224 17632 5549 17660
rect 5224 17620 5230 17632
rect 5537 17629 5549 17632
rect 5583 17660 5595 17663
rect 7009 17663 7067 17669
rect 7009 17660 7021 17663
rect 5583 17632 7021 17660
rect 5583 17629 5595 17632
rect 5537 17623 5595 17629
rect 7009 17629 7021 17632
rect 7055 17660 7067 17663
rect 7561 17663 7619 17669
rect 7561 17660 7573 17663
rect 7055 17632 7573 17660
rect 7055 17629 7067 17632
rect 7009 17623 7067 17629
rect 7561 17629 7573 17632
rect 7607 17629 7619 17663
rect 7561 17623 7619 17629
rect 9674 17620 9680 17672
rect 9732 17660 9738 17672
rect 10594 17660 10600 17672
rect 9732 17632 10600 17660
rect 9732 17620 9738 17632
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 13142 17669 13170 17768
rect 13630 17688 13636 17740
rect 13688 17728 13694 17740
rect 14093 17731 14151 17737
rect 14093 17728 14105 17731
rect 13688 17700 14105 17728
rect 13688 17688 13694 17700
rect 14093 17697 14105 17700
rect 14139 17697 14151 17731
rect 14093 17691 14151 17697
rect 16022 17688 16028 17740
rect 16080 17728 16086 17740
rect 19720 17728 19748 17827
rect 16080 17700 19748 17728
rect 19797 17731 19855 17737
rect 16080 17688 16086 17700
rect 19797 17697 19809 17731
rect 19843 17728 19855 17731
rect 20916 17728 20944 17836
rect 24854 17824 24860 17836
rect 24912 17824 24918 17876
rect 25682 17824 25688 17876
rect 25740 17864 25746 17876
rect 25961 17867 26019 17873
rect 25961 17864 25973 17867
rect 25740 17836 25973 17864
rect 25740 17824 25746 17836
rect 25961 17833 25973 17836
rect 26007 17833 26019 17867
rect 25961 17827 26019 17833
rect 21177 17799 21235 17805
rect 21177 17765 21189 17799
rect 21223 17765 21235 17799
rect 21177 17759 21235 17765
rect 19843 17700 20944 17728
rect 19843 17697 19855 17700
rect 19797 17691 19855 17697
rect 13035 17663 13093 17669
rect 13035 17660 13047 17663
rect 12728 17632 13047 17660
rect 12728 17604 12756 17632
rect 13035 17629 13047 17632
rect 13081 17629 13093 17663
rect 13142 17663 13212 17669
rect 13142 17632 13166 17663
rect 13035 17623 13093 17629
rect 13154 17629 13166 17632
rect 13200 17629 13212 17663
rect 13154 17623 13212 17629
rect 13262 17620 13268 17672
rect 13320 17657 13326 17672
rect 13446 17660 13452 17672
rect 13320 17629 13362 17657
rect 13407 17632 13452 17660
rect 13320 17620 13326 17629
rect 13446 17620 13452 17632
rect 13504 17620 13510 17672
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 14349 17663 14407 17669
rect 14349 17660 14361 17663
rect 13872 17632 14361 17660
rect 13872 17620 13878 17632
rect 14349 17629 14361 17632
rect 14395 17629 14407 17663
rect 14349 17623 14407 17629
rect 19889 17663 19947 17669
rect 19889 17629 19901 17663
rect 19935 17660 19947 17663
rect 19978 17660 19984 17672
rect 19935 17632 19984 17660
rect 19935 17629 19947 17632
rect 19889 17623 19947 17629
rect 19978 17620 19984 17632
rect 20036 17620 20042 17672
rect 20254 17620 20260 17672
rect 20312 17660 20318 17672
rect 20533 17663 20591 17669
rect 20533 17660 20545 17663
rect 20312 17632 20545 17660
rect 20312 17620 20318 17632
rect 20533 17629 20545 17632
rect 20579 17660 20591 17663
rect 21192 17660 21220 17759
rect 22557 17731 22615 17737
rect 22557 17697 22569 17731
rect 22603 17728 22615 17731
rect 24581 17731 24639 17737
rect 24581 17728 24593 17731
rect 22603 17700 24593 17728
rect 22603 17697 22615 17700
rect 22557 17691 22615 17697
rect 24581 17697 24593 17700
rect 24627 17697 24639 17731
rect 24581 17691 24639 17697
rect 20579 17632 21220 17660
rect 23017 17663 23075 17669
rect 20579 17629 20591 17632
rect 20533 17623 20591 17629
rect 23017 17629 23029 17663
rect 23063 17660 23075 17663
rect 23106 17660 23112 17672
rect 23063 17632 23112 17660
rect 23063 17629 23075 17632
rect 23017 17623 23075 17629
rect 23106 17620 23112 17632
rect 23164 17620 23170 17672
rect 23293 17663 23351 17669
rect 23293 17629 23305 17663
rect 23339 17660 23351 17663
rect 24394 17660 24400 17672
rect 23339 17632 24400 17660
rect 23339 17629 23351 17632
rect 23293 17623 23351 17629
rect 24394 17620 24400 17632
rect 24452 17620 24458 17672
rect 24596 17660 24624 17691
rect 25406 17660 25412 17672
rect 24596 17632 25412 17660
rect 25406 17620 25412 17632
rect 25464 17620 25470 17672
rect 25976 17660 26004 17827
rect 29362 17824 29368 17876
rect 29420 17864 29426 17876
rect 30374 17864 30380 17876
rect 29420 17836 30380 17864
rect 29420 17824 29426 17836
rect 30374 17824 30380 17836
rect 30432 17864 30438 17876
rect 33873 17867 33931 17873
rect 33873 17864 33885 17867
rect 30432 17836 33885 17864
rect 30432 17824 30438 17836
rect 31389 17799 31447 17805
rect 31389 17765 31401 17799
rect 31435 17796 31447 17799
rect 31938 17796 31944 17808
rect 31435 17768 31944 17796
rect 31435 17765 31447 17768
rect 31389 17759 31447 17765
rect 31938 17756 31944 17768
rect 31996 17756 32002 17808
rect 32766 17756 32772 17808
rect 32824 17796 32830 17808
rect 32824 17768 33088 17796
rect 32824 17756 32830 17768
rect 32309 17731 32367 17737
rect 32309 17697 32321 17731
rect 32355 17728 32367 17731
rect 32355 17700 32904 17728
rect 32355 17697 32367 17700
rect 32309 17691 32367 17697
rect 26605 17663 26663 17669
rect 26605 17660 26617 17663
rect 25976 17632 26617 17660
rect 26605 17629 26617 17632
rect 26651 17629 26663 17663
rect 29086 17660 29092 17672
rect 26605 17623 26663 17629
rect 26712 17632 29092 17660
rect 4890 17552 4896 17604
rect 4948 17592 4954 17604
rect 12710 17592 12716 17604
rect 4948 17564 12716 17592
rect 4948 17552 4954 17564
rect 12710 17552 12716 17564
rect 12768 17552 12774 17604
rect 20349 17595 20407 17601
rect 20349 17561 20361 17595
rect 20395 17592 20407 17595
rect 20717 17595 20775 17601
rect 20395 17564 20668 17592
rect 20395 17561 20407 17564
rect 20349 17555 20407 17561
rect 12066 17524 12072 17536
rect 12027 17496 12072 17524
rect 12066 17484 12072 17496
rect 12124 17484 12130 17536
rect 12802 17524 12808 17536
rect 12763 17496 12808 17524
rect 12802 17484 12808 17496
rect 12860 17484 12866 17536
rect 12986 17484 12992 17536
rect 13044 17524 13050 17536
rect 14090 17524 14096 17536
rect 13044 17496 14096 17524
rect 13044 17484 13050 17496
rect 14090 17484 14096 17496
rect 14148 17484 14154 17536
rect 14366 17484 14372 17536
rect 14424 17524 14430 17536
rect 15473 17527 15531 17533
rect 15473 17524 15485 17527
rect 14424 17496 15485 17524
rect 14424 17484 14430 17496
rect 15473 17493 15485 17496
rect 15519 17493 15531 17527
rect 15473 17487 15531 17493
rect 19521 17527 19579 17533
rect 19521 17493 19533 17527
rect 19567 17524 19579 17527
rect 20438 17524 20444 17536
rect 19567 17496 20444 17524
rect 19567 17493 19579 17496
rect 19521 17487 19579 17493
rect 20438 17484 20444 17496
rect 20496 17484 20502 17536
rect 20640 17524 20668 17564
rect 20717 17561 20729 17595
rect 20763 17592 20775 17595
rect 20763 17564 21772 17592
rect 20763 17561 20775 17564
rect 20717 17555 20775 17561
rect 20898 17524 20904 17536
rect 20640 17496 20904 17524
rect 20898 17484 20904 17496
rect 20956 17484 20962 17536
rect 21744 17524 21772 17564
rect 21818 17552 21824 17604
rect 21876 17592 21882 17604
rect 22290 17595 22348 17601
rect 22290 17592 22302 17595
rect 21876 17564 22302 17592
rect 21876 17552 21882 17564
rect 22290 17561 22302 17564
rect 22336 17561 22348 17595
rect 22290 17555 22348 17561
rect 24848 17595 24906 17601
rect 24848 17561 24860 17595
rect 24894 17592 24906 17595
rect 25682 17592 25688 17604
rect 24894 17564 25688 17592
rect 24894 17561 24906 17564
rect 24848 17555 24906 17561
rect 25682 17552 25688 17564
rect 25740 17552 25746 17604
rect 26712 17592 26740 17632
rect 29086 17620 29092 17632
rect 29144 17620 29150 17672
rect 31205 17663 31263 17669
rect 31205 17629 31217 17663
rect 31251 17660 31263 17663
rect 31294 17660 31300 17672
rect 31251 17632 31300 17660
rect 31251 17629 31263 17632
rect 31205 17623 31263 17629
rect 31294 17620 31300 17632
rect 31352 17620 31358 17672
rect 31938 17660 31944 17672
rect 31899 17632 31944 17660
rect 31938 17620 31944 17632
rect 31996 17620 32002 17672
rect 32398 17620 32404 17672
rect 32456 17660 32462 17672
rect 32769 17663 32827 17669
rect 32769 17660 32781 17663
rect 32456 17632 32781 17660
rect 32456 17620 32462 17632
rect 32769 17629 32781 17632
rect 32815 17629 32827 17663
rect 32876 17660 32904 17700
rect 33060 17669 33088 17768
rect 33152 17669 33180 17836
rect 33873 17833 33885 17836
rect 33919 17833 33931 17867
rect 37458 17864 37464 17876
rect 37419 17836 37464 17864
rect 33873 17827 33931 17833
rect 37458 17824 37464 17836
rect 37516 17824 37522 17876
rect 40773 17867 40831 17873
rect 40773 17833 40785 17867
rect 40819 17864 40831 17867
rect 41230 17864 41236 17876
rect 40819 17836 41236 17864
rect 40819 17833 40831 17836
rect 40773 17827 40831 17833
rect 41230 17824 41236 17836
rect 41288 17824 41294 17876
rect 35894 17688 35900 17740
rect 35952 17728 35958 17740
rect 36081 17731 36139 17737
rect 36081 17728 36093 17731
rect 35952 17700 36093 17728
rect 35952 17688 35958 17700
rect 36081 17697 36093 17700
rect 36127 17697 36139 17731
rect 38194 17728 38200 17740
rect 38155 17700 38200 17728
rect 36081 17691 36139 17697
rect 38194 17688 38200 17700
rect 38252 17688 38258 17740
rect 41046 17688 41052 17740
rect 41104 17728 41110 17740
rect 41233 17731 41291 17737
rect 41233 17728 41245 17731
rect 41104 17700 41245 17728
rect 41104 17688 41110 17700
rect 41233 17697 41245 17700
rect 41279 17697 41291 17731
rect 41233 17691 41291 17697
rect 32932 17663 32990 17669
rect 32932 17660 32944 17663
rect 32876 17632 32944 17660
rect 32769 17623 32827 17629
rect 32932 17629 32944 17632
rect 32978 17629 32990 17663
rect 32932 17623 32990 17629
rect 33045 17663 33103 17669
rect 33045 17629 33057 17663
rect 33091 17629 33103 17663
rect 33152 17663 33215 17669
rect 33152 17632 33169 17663
rect 33045 17623 33103 17629
rect 33157 17629 33169 17632
rect 33203 17629 33215 17663
rect 37918 17660 37924 17672
rect 37879 17632 37924 17660
rect 33157 17623 33215 17629
rect 37918 17620 37924 17632
rect 37976 17620 37982 17672
rect 25792 17564 26740 17592
rect 26789 17595 26847 17601
rect 22186 17524 22192 17536
rect 21744 17496 22192 17524
rect 22186 17484 22192 17496
rect 22244 17484 22250 17536
rect 25498 17484 25504 17536
rect 25556 17524 25562 17536
rect 25792 17524 25820 17564
rect 26789 17561 26801 17595
rect 26835 17592 26847 17595
rect 27430 17592 27436 17604
rect 26835 17564 27436 17592
rect 26835 17561 26847 17564
rect 26789 17555 26847 17561
rect 27430 17552 27436 17564
rect 27488 17552 27494 17604
rect 32125 17595 32183 17601
rect 32125 17561 32137 17595
rect 32171 17592 32183 17595
rect 34054 17592 34060 17604
rect 32171 17564 34060 17592
rect 32171 17561 32183 17564
rect 32125 17555 32183 17561
rect 34054 17552 34060 17564
rect 34112 17552 34118 17604
rect 36354 17601 36360 17604
rect 36348 17555 36360 17601
rect 36412 17592 36418 17604
rect 38212 17592 38240 17688
rect 38930 17620 38936 17672
rect 38988 17660 38994 17672
rect 40589 17663 40647 17669
rect 40589 17660 40601 17663
rect 38988 17632 40601 17660
rect 38988 17620 38994 17632
rect 40589 17629 40601 17632
rect 40635 17629 40647 17663
rect 40589 17623 40647 17629
rect 40405 17595 40463 17601
rect 40405 17592 40417 17595
rect 36412 17564 36448 17592
rect 38212 17564 40417 17592
rect 36354 17552 36360 17555
rect 36412 17552 36418 17564
rect 40405 17561 40417 17564
rect 40451 17561 40463 17595
rect 40405 17555 40463 17561
rect 25556 17496 25820 17524
rect 25556 17484 25562 17496
rect 26142 17484 26148 17536
rect 26200 17524 26206 17536
rect 26421 17527 26479 17533
rect 26421 17524 26433 17527
rect 26200 17496 26433 17524
rect 26200 17484 26206 17496
rect 26421 17493 26433 17496
rect 26467 17493 26479 17527
rect 33410 17524 33416 17536
rect 33371 17496 33416 17524
rect 26421 17487 26479 17493
rect 33410 17484 33416 17496
rect 33468 17484 33474 17536
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 11422 17280 11428 17332
rect 11480 17320 11486 17332
rect 11517 17323 11575 17329
rect 11517 17320 11529 17323
rect 11480 17292 11529 17320
rect 11480 17280 11486 17292
rect 11517 17289 11529 17292
rect 11563 17289 11575 17323
rect 11517 17283 11575 17289
rect 12989 17323 13047 17329
rect 12989 17289 13001 17323
rect 13035 17320 13047 17323
rect 13262 17320 13268 17332
rect 13035 17292 13268 17320
rect 13035 17289 13047 17292
rect 12989 17283 13047 17289
rect 13262 17280 13268 17292
rect 13320 17280 13326 17332
rect 13906 17320 13912 17332
rect 13867 17292 13912 17320
rect 13906 17280 13912 17292
rect 13964 17280 13970 17332
rect 14090 17280 14096 17332
rect 14148 17320 14154 17332
rect 16669 17323 16727 17329
rect 16669 17320 16681 17323
rect 14148 17292 16681 17320
rect 14148 17280 14154 17292
rect 16669 17289 16681 17292
rect 16715 17320 16727 17323
rect 16850 17320 16856 17332
rect 16715 17292 16856 17320
rect 16715 17289 16727 17292
rect 16669 17283 16727 17289
rect 16850 17280 16856 17292
rect 16908 17280 16914 17332
rect 21818 17320 21824 17332
rect 21779 17292 21824 17320
rect 21818 17280 21824 17292
rect 21876 17280 21882 17332
rect 25498 17320 25504 17332
rect 21928 17292 25504 17320
rect 1854 17212 1860 17264
rect 1912 17252 1918 17264
rect 2685 17255 2743 17261
rect 2685 17252 2697 17255
rect 1912 17224 2697 17252
rect 1912 17212 1918 17224
rect 2685 17221 2697 17224
rect 2731 17252 2743 17255
rect 2774 17252 2780 17264
rect 2731 17224 2780 17252
rect 2731 17221 2743 17224
rect 2685 17215 2743 17221
rect 2774 17212 2780 17224
rect 2832 17212 2838 17264
rect 6546 17212 6552 17264
rect 6604 17252 6610 17264
rect 6733 17255 6791 17261
rect 6733 17252 6745 17255
rect 6604 17224 6745 17252
rect 6604 17212 6610 17224
rect 6733 17221 6745 17224
rect 6779 17221 6791 17255
rect 12066 17252 12072 17264
rect 6733 17215 6791 17221
rect 9646 17224 12072 17252
rect 9646 17196 9674 17224
rect 12066 17212 12072 17224
rect 12124 17212 12130 17264
rect 12342 17212 12348 17264
rect 12400 17252 12406 17264
rect 12621 17255 12679 17261
rect 12621 17252 12633 17255
rect 12400 17224 12633 17252
rect 12400 17212 12406 17224
rect 12621 17221 12633 17224
rect 12667 17252 12679 17255
rect 14277 17255 14335 17261
rect 14277 17252 14289 17255
rect 12667 17224 14289 17252
rect 12667 17221 12679 17224
rect 12621 17215 12679 17221
rect 14277 17221 14289 17224
rect 14323 17221 14335 17255
rect 14277 17215 14335 17221
rect 4433 17187 4491 17193
rect 4433 17153 4445 17187
rect 4479 17184 4491 17187
rect 4982 17184 4988 17196
rect 4479 17156 4988 17184
rect 4479 17153 4491 17156
rect 4433 17147 4491 17153
rect 4982 17144 4988 17156
rect 5040 17144 5046 17196
rect 5994 17144 6000 17196
rect 6052 17184 6058 17196
rect 7101 17187 7159 17193
rect 7101 17184 7113 17187
rect 6052 17156 7113 17184
rect 6052 17144 6058 17156
rect 7101 17153 7113 17156
rect 7147 17153 7159 17187
rect 9582 17184 9588 17196
rect 9495 17156 9588 17184
rect 7101 17147 7159 17153
rect 9582 17144 9588 17156
rect 9640 17156 9674 17196
rect 9852 17187 9910 17193
rect 9640 17144 9646 17156
rect 9852 17153 9864 17187
rect 9898 17184 9910 17187
rect 10318 17184 10324 17196
rect 9898 17156 10324 17184
rect 9898 17153 9910 17156
rect 9852 17147 9910 17153
rect 10318 17144 10324 17156
rect 10376 17144 10382 17196
rect 11606 17184 11612 17196
rect 10980 17156 11612 17184
rect 10980 17057 11008 17156
rect 11606 17144 11612 17156
rect 11664 17184 11670 17196
rect 11701 17187 11759 17193
rect 11701 17184 11713 17187
rect 11664 17156 11713 17184
rect 11664 17144 11670 17156
rect 11701 17153 11713 17156
rect 11747 17153 11759 17187
rect 11701 17147 11759 17153
rect 11885 17187 11943 17193
rect 11885 17153 11897 17187
rect 11931 17184 11943 17187
rect 12360 17184 12388 17212
rect 11931 17156 12388 17184
rect 11931 17153 11943 17156
rect 11885 17147 11943 17153
rect 12526 17144 12532 17196
rect 12584 17184 12590 17196
rect 12805 17187 12863 17193
rect 12805 17184 12817 17187
rect 12584 17156 12817 17184
rect 12584 17144 12590 17156
rect 12805 17153 12817 17156
rect 12851 17153 12863 17187
rect 12805 17147 12863 17153
rect 14093 17187 14151 17193
rect 14093 17153 14105 17187
rect 14139 17184 14151 17187
rect 14366 17184 14372 17196
rect 14139 17156 14372 17184
rect 14139 17153 14151 17156
rect 14093 17147 14151 17153
rect 14366 17144 14372 17156
rect 14424 17144 14430 17196
rect 15194 17184 15200 17196
rect 15155 17156 15200 17184
rect 15194 17144 15200 17156
rect 15252 17144 15258 17196
rect 15286 17144 15292 17196
rect 15344 17184 15350 17196
rect 21928 17184 21956 17292
rect 25498 17280 25504 17292
rect 25556 17280 25562 17332
rect 25682 17320 25688 17332
rect 25643 17292 25688 17320
rect 25682 17280 25688 17292
rect 25740 17280 25746 17332
rect 26694 17320 26700 17332
rect 26068 17292 26700 17320
rect 23382 17252 23388 17264
rect 22201 17224 23388 17252
rect 22201 17199 22229 17224
rect 23382 17212 23388 17224
rect 23440 17212 23446 17264
rect 26068 17199 26096 17292
rect 26694 17280 26700 17292
rect 26752 17280 26758 17332
rect 27246 17280 27252 17332
rect 27304 17320 27310 17332
rect 29178 17320 29184 17332
rect 27304 17292 29184 17320
rect 27304 17280 27310 17292
rect 29178 17280 29184 17292
rect 29236 17280 29242 17332
rect 33502 17280 33508 17332
rect 33560 17320 33566 17332
rect 34606 17320 34612 17332
rect 33560 17292 34612 17320
rect 33560 17280 33566 17292
rect 34606 17280 34612 17292
rect 34664 17280 34670 17332
rect 34977 17323 35035 17329
rect 34977 17289 34989 17323
rect 35023 17289 35035 17323
rect 36354 17320 36360 17332
rect 34977 17283 35035 17289
rect 35973 17292 36216 17320
rect 36315 17292 36360 17320
rect 26602 17212 26608 17264
rect 26660 17252 26666 17264
rect 30650 17252 30656 17264
rect 26660 17224 30656 17252
rect 26660 17212 26666 17224
rect 30650 17212 30656 17224
rect 30708 17212 30714 17264
rect 33137 17255 33195 17261
rect 33137 17221 33149 17255
rect 33183 17252 33195 17255
rect 33842 17255 33900 17261
rect 33842 17252 33854 17255
rect 33183 17224 33854 17252
rect 33183 17221 33195 17224
rect 33137 17215 33195 17221
rect 33842 17221 33854 17224
rect 33888 17221 33900 17255
rect 33842 17215 33900 17221
rect 34422 17212 34428 17264
rect 34480 17252 34486 17264
rect 34992 17252 35020 17283
rect 34480 17224 35020 17252
rect 34480 17212 34486 17224
rect 22170 17193 22229 17199
rect 15344 17156 21956 17184
rect 22051 17187 22109 17193
rect 15344 17144 15350 17156
rect 22051 17153 22063 17187
rect 22097 17153 22109 17187
rect 22170 17159 22182 17193
rect 22216 17159 22229 17193
rect 22170 17153 22229 17159
rect 22051 17147 22109 17153
rect 13262 17076 13268 17128
rect 13320 17116 13326 17128
rect 14458 17116 14464 17128
rect 13320 17088 14464 17116
rect 13320 17076 13326 17088
rect 14458 17076 14464 17088
rect 14516 17076 14522 17128
rect 14918 17116 14924 17128
rect 14879 17088 14924 17116
rect 14918 17076 14924 17088
rect 14976 17076 14982 17128
rect 16574 17076 16580 17128
rect 16632 17116 16638 17128
rect 21910 17116 21916 17128
rect 16632 17088 21916 17116
rect 16632 17076 16638 17088
rect 21910 17076 21916 17088
rect 21968 17076 21974 17128
rect 10965 17051 11023 17057
rect 10965 17017 10977 17051
rect 11011 17017 11023 17051
rect 10965 17011 11023 17017
rect 11698 17008 11704 17060
rect 11756 17048 11762 17060
rect 17497 17051 17555 17057
rect 17497 17048 17509 17051
rect 11756 17020 17509 17048
rect 11756 17008 11762 17020
rect 17497 17017 17509 17020
rect 17543 17048 17555 17051
rect 18138 17048 18144 17060
rect 17543 17020 18144 17048
rect 17543 17017 17555 17020
rect 17497 17011 17555 17017
rect 18138 17008 18144 17020
rect 18196 17008 18202 17060
rect 5166 16980 5172 16992
rect 5127 16952 5172 16980
rect 5166 16940 5172 16952
rect 5224 16940 5230 16992
rect 5813 16983 5871 16989
rect 5813 16949 5825 16983
rect 5859 16980 5871 16983
rect 5994 16980 6000 16992
rect 5859 16952 6000 16980
rect 5859 16949 5871 16952
rect 5813 16943 5871 16949
rect 5994 16940 6000 16952
rect 6052 16940 6058 16992
rect 10594 16940 10600 16992
rect 10652 16980 10658 16992
rect 19334 16980 19340 16992
rect 10652 16952 19340 16980
rect 10652 16940 10658 16952
rect 19334 16940 19340 16952
rect 19392 16940 19398 16992
rect 21266 16980 21272 16992
rect 21227 16952 21272 16980
rect 21266 16940 21272 16952
rect 21324 16980 21330 16992
rect 22066 16980 22094 17147
rect 22201 17048 22229 17153
rect 22278 17144 22284 17196
rect 22336 17187 22342 17196
rect 22465 17187 22523 17193
rect 22336 17159 22378 17187
rect 22336 17144 22342 17159
rect 22465 17153 22477 17187
rect 22511 17184 22523 17187
rect 22554 17184 22560 17196
rect 22511 17156 22560 17184
rect 22511 17153 22523 17156
rect 22465 17147 22523 17153
rect 22554 17144 22560 17156
rect 22612 17144 22618 17196
rect 26050 17193 26108 17199
rect 25961 17187 26019 17193
rect 25961 17184 25973 17187
rect 25148 17156 25973 17184
rect 23014 17116 23020 17128
rect 22975 17088 23020 17116
rect 23014 17076 23020 17088
rect 23072 17076 23078 17128
rect 23658 17116 23664 17128
rect 23619 17088 23664 17116
rect 23658 17076 23664 17088
rect 23716 17076 23722 17128
rect 23937 17119 23995 17125
rect 23937 17085 23949 17119
rect 23983 17116 23995 17119
rect 24946 17116 24952 17128
rect 23983 17088 24952 17116
rect 23983 17085 23995 17088
rect 23937 17079 23995 17085
rect 24946 17076 24952 17088
rect 25004 17076 25010 17128
rect 22278 17048 22284 17060
rect 22201 17020 22284 17048
rect 22278 17008 22284 17020
rect 22336 17008 22342 17060
rect 22554 17008 22560 17060
rect 22612 17048 22618 17060
rect 23032 17048 23060 17076
rect 22612 17020 23060 17048
rect 22612 17008 22618 17020
rect 25148 16989 25176 17156
rect 25961 17153 25973 17156
rect 26007 17153 26019 17187
rect 26050 17159 26062 17193
rect 26096 17159 26108 17193
rect 26050 17153 26108 17159
rect 25961 17147 26019 17153
rect 26142 17144 26148 17196
rect 26200 17184 26206 17196
rect 26329 17187 26387 17193
rect 26200 17156 26245 17184
rect 26200 17144 26206 17156
rect 26329 17153 26341 17187
rect 26375 17153 26387 17187
rect 26329 17147 26387 17153
rect 25314 17008 25320 17060
rect 25372 17048 25378 17060
rect 26142 17048 26148 17060
rect 25372 17020 26148 17048
rect 25372 17008 25378 17020
rect 26142 17008 26148 17020
rect 26200 17048 26206 17060
rect 26344 17048 26372 17147
rect 26786 17144 26792 17196
rect 26844 17184 26850 17196
rect 27229 17187 27287 17193
rect 27229 17184 27241 17187
rect 26844 17156 27241 17184
rect 26844 17144 26850 17156
rect 27229 17153 27241 17156
rect 27275 17153 27287 17187
rect 27229 17147 27287 17153
rect 29822 17144 29828 17196
rect 29880 17184 29886 17196
rect 30006 17184 30012 17196
rect 29880 17156 30012 17184
rect 29880 17144 29886 17156
rect 30006 17144 30012 17156
rect 30064 17144 30070 17196
rect 30193 17187 30251 17193
rect 30193 17153 30205 17187
rect 30239 17184 30251 17187
rect 31386 17184 31392 17196
rect 30239 17156 31392 17184
rect 30239 17153 30251 17156
rect 30193 17147 30251 17153
rect 31386 17144 31392 17156
rect 31444 17144 31450 17196
rect 32398 17144 32404 17196
rect 32456 17184 32462 17196
rect 32493 17187 32551 17193
rect 32493 17184 32505 17187
rect 32456 17156 32505 17184
rect 32456 17144 32462 17156
rect 32493 17153 32505 17156
rect 32539 17153 32551 17187
rect 32493 17147 32551 17153
rect 32582 17144 32588 17196
rect 32640 17184 32646 17196
rect 32677 17187 32735 17193
rect 32677 17184 32689 17187
rect 32640 17156 32689 17184
rect 32640 17144 32646 17156
rect 32677 17153 32689 17156
rect 32723 17153 32735 17187
rect 32677 17147 32735 17153
rect 32766 17144 32772 17196
rect 32824 17184 32830 17196
rect 32907 17187 32965 17193
rect 32824 17156 32869 17184
rect 32824 17144 32830 17156
rect 32907 17153 32919 17187
rect 32953 17184 32965 17187
rect 32953 17153 32975 17184
rect 32907 17147 32975 17153
rect 26970 17116 26976 17128
rect 26931 17088 26976 17116
rect 26970 17076 26976 17088
rect 27028 17076 27034 17128
rect 28718 17076 28724 17128
rect 28776 17116 28782 17128
rect 30926 17116 30932 17128
rect 28776 17088 30932 17116
rect 28776 17076 28782 17088
rect 30926 17076 30932 17088
rect 30984 17076 30990 17128
rect 31570 17076 31576 17128
rect 31628 17116 31634 17128
rect 32947 17116 32975 17147
rect 35618 17144 35624 17196
rect 35676 17184 35682 17196
rect 35973 17193 36001 17292
rect 35713 17187 35771 17193
rect 35713 17184 35725 17187
rect 35676 17156 35725 17184
rect 35676 17144 35682 17156
rect 35713 17153 35725 17156
rect 35759 17153 35771 17187
rect 35713 17147 35771 17153
rect 35876 17187 35934 17193
rect 35876 17153 35888 17187
rect 35922 17184 35934 17187
rect 35973 17187 36047 17193
rect 35922 17153 35940 17184
rect 35973 17156 36001 17187
rect 35876 17147 35940 17153
rect 35989 17153 36001 17156
rect 36035 17153 36047 17187
rect 35989 17147 36047 17153
rect 33594 17116 33600 17128
rect 31628 17088 32975 17116
rect 33555 17088 33600 17116
rect 31628 17076 31634 17088
rect 33594 17076 33600 17088
rect 33652 17076 33658 17128
rect 35912 17116 35940 17147
rect 36078 17144 36084 17196
rect 36136 17193 36142 17196
rect 36136 17187 36159 17193
rect 36147 17153 36159 17187
rect 36188 17184 36216 17292
rect 36354 17280 36360 17292
rect 36412 17280 36418 17332
rect 37458 17252 37464 17264
rect 37419 17224 37464 17252
rect 37458 17212 37464 17224
rect 37516 17212 37522 17264
rect 37645 17255 37703 17261
rect 37645 17221 37657 17255
rect 37691 17252 37703 17255
rect 37918 17252 37924 17264
rect 37691 17224 37924 17252
rect 37691 17221 37703 17224
rect 37645 17215 37703 17221
rect 37918 17212 37924 17224
rect 37976 17212 37982 17264
rect 37550 17184 37556 17196
rect 36188 17156 37556 17184
rect 36136 17147 36159 17153
rect 36136 17144 36142 17147
rect 37550 17144 37556 17156
rect 37608 17144 37614 17196
rect 38746 17184 38752 17196
rect 38707 17156 38752 17184
rect 38746 17144 38752 17156
rect 38804 17144 38810 17196
rect 37277 17119 37335 17125
rect 37277 17116 37289 17119
rect 35912 17088 37289 17116
rect 37277 17085 37289 17088
rect 37323 17085 37335 17119
rect 37277 17079 37335 17085
rect 39025 17119 39083 17125
rect 39025 17085 39037 17119
rect 39071 17116 39083 17119
rect 39850 17116 39856 17128
rect 39071 17088 39856 17116
rect 39071 17085 39083 17088
rect 39025 17079 39083 17085
rect 39850 17076 39856 17088
rect 39908 17076 39914 17128
rect 58158 17048 58164 17060
rect 26200 17020 26372 17048
rect 27908 17020 31754 17048
rect 58119 17020 58164 17048
rect 26200 17008 26206 17020
rect 25133 16983 25191 16989
rect 25133 16980 25145 16983
rect 21324 16952 25145 16980
rect 21324 16940 21330 16952
rect 25133 16949 25145 16952
rect 25179 16949 25191 16983
rect 25133 16943 25191 16949
rect 25498 16940 25504 16992
rect 25556 16980 25562 16992
rect 27908 16980 27936 17020
rect 28350 16980 28356 16992
rect 25556 16952 27936 16980
rect 28311 16952 28356 16980
rect 25556 16940 25562 16952
rect 28350 16940 28356 16952
rect 28408 16940 28414 16992
rect 29362 16940 29368 16992
rect 29420 16980 29426 16992
rect 29825 16983 29883 16989
rect 29825 16980 29837 16983
rect 29420 16952 29837 16980
rect 29420 16940 29426 16952
rect 29825 16949 29837 16952
rect 29871 16949 29883 16983
rect 31570 16980 31576 16992
rect 31531 16952 31576 16980
rect 29825 16943 29883 16949
rect 31570 16940 31576 16952
rect 31628 16940 31634 16992
rect 31726 16980 31754 17020
rect 58158 17008 58164 17020
rect 58216 17008 58222 17060
rect 33962 16980 33968 16992
rect 31726 16952 33968 16980
rect 33962 16940 33968 16952
rect 34020 16940 34026 16992
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 3234 16776 3240 16788
rect 3195 16748 3240 16776
rect 3234 16736 3240 16748
rect 3292 16736 3298 16788
rect 4982 16776 4988 16788
rect 4895 16748 4988 16776
rect 4982 16736 4988 16748
rect 5040 16776 5046 16788
rect 9674 16776 9680 16788
rect 5040 16748 9680 16776
rect 5040 16736 5046 16748
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 22462 16776 22468 16788
rect 9784 16748 22468 16776
rect 4341 16711 4399 16717
rect 4341 16677 4353 16711
rect 4387 16708 4399 16711
rect 4890 16708 4896 16720
rect 4387 16680 4896 16708
rect 4387 16677 4399 16680
rect 4341 16671 4399 16677
rect 4890 16668 4896 16680
rect 4948 16668 4954 16720
rect 1854 16640 1860 16652
rect 1815 16612 1860 16640
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 8389 16643 8447 16649
rect 8389 16609 8401 16643
rect 8435 16640 8447 16643
rect 9582 16640 9588 16652
rect 8435 16612 9588 16640
rect 8435 16609 8447 16612
rect 8389 16603 8447 16609
rect 9582 16600 9588 16612
rect 9640 16600 9646 16652
rect 1946 16532 1952 16584
rect 2004 16572 2010 16584
rect 2113 16575 2171 16581
rect 2113 16572 2125 16575
rect 2004 16544 2125 16572
rect 2004 16532 2010 16544
rect 2113 16541 2125 16544
rect 2159 16541 2171 16575
rect 2113 16535 2171 16541
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16572 4215 16575
rect 5994 16572 6000 16584
rect 4203 16544 6000 16572
rect 4203 16541 4215 16544
rect 4157 16535 4215 16541
rect 5994 16532 6000 16544
rect 6052 16532 6058 16584
rect 9398 16532 9404 16584
rect 9456 16572 9462 16584
rect 9784 16572 9812 16748
rect 22462 16736 22468 16748
rect 22520 16736 22526 16788
rect 24854 16776 24860 16788
rect 24815 16748 24860 16776
rect 24854 16736 24860 16748
rect 24912 16736 24918 16788
rect 25038 16776 25044 16788
rect 24999 16748 25044 16776
rect 25038 16736 25044 16748
rect 25096 16736 25102 16788
rect 26786 16776 26792 16788
rect 26747 16748 26792 16776
rect 26786 16736 26792 16748
rect 26844 16736 26850 16788
rect 27430 16776 27436 16788
rect 27343 16748 27436 16776
rect 27430 16736 27436 16748
rect 27488 16776 27494 16788
rect 31294 16776 31300 16788
rect 27488 16748 31300 16776
rect 27488 16736 27494 16748
rect 31294 16736 31300 16748
rect 31352 16736 31358 16788
rect 34054 16736 34060 16788
rect 34112 16776 34118 16788
rect 34149 16779 34207 16785
rect 34149 16776 34161 16779
rect 34112 16748 34161 16776
rect 34112 16736 34118 16748
rect 34149 16745 34161 16748
rect 34195 16745 34207 16779
rect 34149 16739 34207 16745
rect 35618 16736 35624 16788
rect 35676 16776 35682 16788
rect 36262 16776 36268 16788
rect 35676 16748 36268 16776
rect 35676 16736 35682 16748
rect 36262 16736 36268 16748
rect 36320 16736 36326 16788
rect 39117 16779 39175 16785
rect 39117 16745 39129 16779
rect 39163 16776 39175 16779
rect 40678 16776 40684 16788
rect 39163 16748 40684 16776
rect 39163 16745 39175 16748
rect 39117 16739 39175 16745
rect 40678 16736 40684 16748
rect 40736 16736 40742 16788
rect 9858 16668 9864 16720
rect 9916 16708 9922 16720
rect 11609 16711 11667 16717
rect 11609 16708 11621 16711
rect 9916 16680 11621 16708
rect 9916 16668 9922 16680
rect 11609 16677 11621 16680
rect 11655 16677 11667 16711
rect 11609 16671 11667 16677
rect 12161 16711 12219 16717
rect 12161 16677 12173 16711
rect 12207 16708 12219 16711
rect 12986 16708 12992 16720
rect 12207 16680 12992 16708
rect 12207 16677 12219 16680
rect 12161 16671 12219 16677
rect 10226 16600 10232 16652
rect 10284 16640 10290 16652
rect 12176 16640 12204 16671
rect 12986 16668 12992 16680
rect 13044 16668 13050 16720
rect 20349 16711 20407 16717
rect 16500 16680 17632 16708
rect 12710 16640 12716 16652
rect 10284 16612 12204 16640
rect 12671 16612 12716 16640
rect 10284 16600 10290 16612
rect 12710 16600 12716 16612
rect 12768 16640 12774 16652
rect 14829 16643 14887 16649
rect 14829 16640 14841 16643
rect 12768 16612 14841 16640
rect 12768 16600 12774 16612
rect 14829 16609 14841 16612
rect 14875 16640 14887 16643
rect 16500 16640 16528 16680
rect 17604 16640 17632 16680
rect 20349 16677 20361 16711
rect 20395 16708 20407 16711
rect 20714 16708 20720 16720
rect 20395 16680 20720 16708
rect 20395 16677 20407 16680
rect 20349 16671 20407 16677
rect 20714 16668 20720 16680
rect 20772 16668 20778 16720
rect 18598 16640 18604 16652
rect 14875 16612 15700 16640
rect 14875 16609 14887 16612
rect 14829 16603 14887 16609
rect 10962 16572 10968 16584
rect 9456 16544 9812 16572
rect 10923 16544 10968 16572
rect 9456 16532 9462 16544
rect 10962 16532 10968 16544
rect 11020 16532 11026 16584
rect 11054 16532 11060 16584
rect 11112 16572 11118 16584
rect 11471 16575 11529 16581
rect 11112 16544 11157 16572
rect 11112 16532 11118 16544
rect 11471 16541 11483 16575
rect 11517 16572 11529 16575
rect 11698 16572 11704 16584
rect 11517 16544 11704 16572
rect 11517 16541 11529 16544
rect 11471 16535 11529 16541
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 15672 16581 15700 16612
rect 16040 16612 16528 16640
rect 15657 16575 15715 16581
rect 15657 16541 15669 16575
rect 15703 16541 15715 16575
rect 15657 16535 15715 16541
rect 15749 16575 15807 16581
rect 15749 16541 15761 16575
rect 15795 16541 15807 16575
rect 15749 16535 15807 16541
rect 7558 16464 7564 16516
rect 7616 16504 7622 16516
rect 8122 16507 8180 16513
rect 8122 16504 8134 16507
rect 7616 16476 8134 16504
rect 7616 16464 7622 16476
rect 8122 16473 8134 16476
rect 8168 16473 8180 16507
rect 11238 16504 11244 16516
rect 11199 16476 11244 16504
rect 8122 16467 8180 16473
rect 11238 16464 11244 16476
rect 11296 16464 11302 16516
rect 11333 16507 11391 16513
rect 11333 16473 11345 16507
rect 11379 16504 11391 16507
rect 13906 16504 13912 16516
rect 11379 16476 13912 16504
rect 11379 16473 11391 16476
rect 11333 16467 11391 16473
rect 13906 16464 13912 16476
rect 13964 16464 13970 16516
rect 15764 16504 15792 16535
rect 15838 16532 15844 16584
rect 15896 16572 15902 16584
rect 16040 16581 16068 16612
rect 16500 16581 16528 16612
rect 16592 16612 17080 16640
rect 16025 16575 16083 16581
rect 15896 16544 15941 16572
rect 15896 16532 15902 16544
rect 16025 16541 16037 16575
rect 16071 16541 16083 16575
rect 16025 16535 16083 16541
rect 16485 16575 16543 16581
rect 16485 16541 16497 16575
rect 16531 16541 16543 16575
rect 16485 16535 16543 16541
rect 16592 16504 16620 16612
rect 16776 16581 16804 16612
rect 16669 16575 16727 16581
rect 16669 16541 16681 16575
rect 16715 16541 16727 16575
rect 16669 16535 16727 16541
rect 16761 16575 16819 16581
rect 16761 16541 16773 16575
rect 16807 16541 16819 16575
rect 16761 16535 16819 16541
rect 15764 16476 16620 16504
rect 16684 16504 16712 16535
rect 16850 16532 16856 16584
rect 16908 16572 16914 16584
rect 17052 16572 17080 16612
rect 17604 16612 18604 16640
rect 17126 16572 17132 16584
rect 16908 16544 16953 16572
rect 17052 16544 17132 16572
rect 16908 16532 16914 16544
rect 17126 16532 17132 16544
rect 17184 16572 17190 16584
rect 17604 16581 17632 16612
rect 18598 16600 18604 16612
rect 18656 16600 18662 16652
rect 20254 16600 20260 16652
rect 20312 16640 20318 16652
rect 20809 16643 20867 16649
rect 20809 16640 20821 16643
rect 20312 16612 20821 16640
rect 20312 16600 20318 16612
rect 20809 16609 20821 16612
rect 20855 16609 20867 16643
rect 20809 16603 20867 16609
rect 22094 16600 22100 16652
rect 22152 16640 22158 16652
rect 22738 16640 22744 16652
rect 22152 16612 22744 16640
rect 22152 16600 22158 16612
rect 22738 16600 22744 16612
rect 22796 16640 22802 16652
rect 22833 16643 22891 16649
rect 22833 16640 22845 16643
rect 22796 16612 22845 16640
rect 22796 16600 22802 16612
rect 22833 16609 22845 16612
rect 22879 16609 22891 16643
rect 22833 16603 22891 16609
rect 22922 16600 22928 16652
rect 22980 16640 22986 16652
rect 25133 16643 25191 16649
rect 25133 16640 25145 16643
rect 22980 16612 25145 16640
rect 22980 16600 22986 16612
rect 25133 16609 25145 16612
rect 25179 16609 25191 16643
rect 26694 16640 26700 16652
rect 25133 16603 25191 16609
rect 26436 16612 26700 16640
rect 17589 16575 17647 16581
rect 17184 16544 17540 16572
rect 17184 16532 17190 16544
rect 17310 16504 17316 16516
rect 16684 16476 17316 16504
rect 17310 16464 17316 16476
rect 17368 16464 17374 16516
rect 17512 16504 17540 16544
rect 17589 16541 17601 16575
rect 17635 16541 17647 16575
rect 17770 16572 17776 16584
rect 17731 16544 17776 16572
rect 17589 16535 17647 16541
rect 17770 16532 17776 16544
rect 17828 16532 17834 16584
rect 17865 16575 17923 16581
rect 17865 16541 17877 16575
rect 17911 16541 17923 16575
rect 17865 16535 17923 16541
rect 17957 16575 18015 16581
rect 17957 16541 17969 16575
rect 18003 16572 18015 16575
rect 18138 16572 18144 16584
rect 18003 16544 18144 16572
rect 18003 16541 18015 16544
rect 17957 16535 18015 16541
rect 17880 16504 17908 16535
rect 18138 16532 18144 16544
rect 18196 16532 18202 16584
rect 23106 16572 23112 16584
rect 23067 16544 23112 16572
rect 23106 16532 23112 16544
rect 23164 16532 23170 16584
rect 25038 16572 25044 16584
rect 24999 16544 25044 16572
rect 25038 16532 25044 16544
rect 25096 16532 25102 16584
rect 25317 16575 25375 16581
rect 25317 16541 25329 16575
rect 25363 16572 25375 16575
rect 25498 16572 25504 16584
rect 25363 16544 25504 16572
rect 25363 16541 25375 16544
rect 25317 16535 25375 16541
rect 25498 16532 25504 16544
rect 25556 16532 25562 16584
rect 26142 16532 26148 16584
rect 26200 16581 26206 16584
rect 26200 16572 26209 16581
rect 26326 16572 26332 16584
rect 26200 16544 26245 16572
rect 26287 16544 26332 16572
rect 26200 16535 26209 16544
rect 26200 16532 26206 16535
rect 26326 16532 26332 16544
rect 26384 16532 26390 16584
rect 26436 16581 26464 16612
rect 26694 16600 26700 16612
rect 26752 16600 26758 16652
rect 27246 16600 27252 16652
rect 27304 16640 27310 16652
rect 27801 16643 27859 16649
rect 27801 16640 27813 16643
rect 27304 16612 27813 16640
rect 27304 16600 27310 16612
rect 27801 16609 27813 16612
rect 27847 16609 27859 16643
rect 32769 16643 32827 16649
rect 32769 16640 32781 16643
rect 27801 16603 27859 16609
rect 30668 16612 32781 16640
rect 26421 16575 26479 16581
rect 26421 16541 26433 16575
rect 26467 16541 26479 16575
rect 26421 16535 26479 16541
rect 26513 16575 26571 16581
rect 26513 16541 26525 16575
rect 26559 16572 26571 16575
rect 26602 16572 26608 16584
rect 26559 16544 26608 16572
rect 26559 16541 26571 16544
rect 26513 16535 26571 16541
rect 26602 16532 26608 16544
rect 26660 16532 26666 16584
rect 27522 16532 27528 16584
rect 27580 16572 27586 16584
rect 27617 16575 27675 16581
rect 27617 16572 27629 16575
rect 27580 16544 27629 16572
rect 27580 16532 27586 16544
rect 27617 16541 27629 16544
rect 27663 16541 27675 16575
rect 27617 16535 27675 16541
rect 29546 16532 29552 16584
rect 29604 16572 29610 16584
rect 29641 16575 29699 16581
rect 29641 16572 29653 16575
rect 29604 16544 29653 16572
rect 29604 16532 29610 16544
rect 29641 16541 29653 16544
rect 29687 16572 29699 16575
rect 30668 16572 30696 16612
rect 32769 16609 32781 16612
rect 32815 16640 32827 16643
rect 32815 16612 32904 16640
rect 32815 16609 32827 16612
rect 32769 16603 32827 16609
rect 29687 16544 30696 16572
rect 31481 16575 31539 16581
rect 29687 16541 29699 16544
rect 29641 16535 29699 16541
rect 31481 16541 31493 16575
rect 31527 16541 31539 16575
rect 31481 16535 31539 16541
rect 31757 16575 31815 16581
rect 31757 16541 31769 16575
rect 31803 16572 31815 16575
rect 32674 16572 32680 16584
rect 31803 16544 32680 16572
rect 31803 16541 31815 16544
rect 31757 16535 31815 16541
rect 17512 16476 17908 16504
rect 26234 16464 26240 16516
rect 26292 16504 26298 16516
rect 28350 16504 28356 16516
rect 26292 16476 28356 16504
rect 26292 16464 26298 16476
rect 28350 16464 28356 16476
rect 28408 16464 28414 16516
rect 28902 16464 28908 16516
rect 28960 16504 28966 16516
rect 29886 16507 29944 16513
rect 29886 16504 29898 16507
rect 28960 16476 29898 16504
rect 28960 16464 28966 16476
rect 29886 16473 29898 16476
rect 29932 16473 29944 16507
rect 29886 16467 29944 16473
rect 30098 16464 30104 16516
rect 30156 16504 30162 16516
rect 31496 16504 31524 16535
rect 32674 16532 32680 16544
rect 32732 16532 32738 16584
rect 32876 16572 32904 16612
rect 33594 16572 33600 16584
rect 32876 16544 33600 16572
rect 33594 16532 33600 16544
rect 33652 16532 33658 16584
rect 36998 16572 37004 16584
rect 36959 16544 37004 16572
rect 36998 16532 37004 16544
rect 37056 16532 37062 16584
rect 37093 16575 37151 16581
rect 37093 16541 37105 16575
rect 37139 16572 37151 16575
rect 37369 16575 37427 16581
rect 37139 16544 37320 16572
rect 37139 16541 37151 16544
rect 37093 16535 37151 16541
rect 30156 16476 31524 16504
rect 33036 16507 33094 16513
rect 30156 16464 30162 16476
rect 33036 16473 33048 16507
rect 33082 16504 33094 16507
rect 33410 16504 33416 16516
rect 33082 16476 33416 16504
rect 33082 16473 33094 16476
rect 33036 16467 33094 16473
rect 33410 16464 33416 16476
rect 33468 16464 33474 16516
rect 37182 16504 37188 16516
rect 37143 16476 37188 16504
rect 37182 16464 37188 16476
rect 37240 16464 37246 16516
rect 37292 16504 37320 16544
rect 37369 16541 37381 16575
rect 37415 16572 37427 16575
rect 38654 16572 38660 16584
rect 37415 16544 38660 16572
rect 37415 16541 37427 16544
rect 37369 16535 37427 16541
rect 38654 16532 38660 16544
rect 38712 16532 38718 16584
rect 40037 16575 40095 16581
rect 40037 16572 40049 16575
rect 39132 16544 40049 16572
rect 39132 16504 39160 16544
rect 40037 16541 40049 16544
rect 40083 16572 40095 16575
rect 40218 16572 40224 16584
rect 40083 16544 40224 16572
rect 40083 16541 40095 16544
rect 40037 16535 40095 16541
rect 40218 16532 40224 16544
rect 40276 16532 40282 16584
rect 37292 16476 39160 16504
rect 39206 16464 39212 16516
rect 39264 16504 39270 16516
rect 39850 16504 39856 16516
rect 39264 16476 39309 16504
rect 39811 16476 39856 16504
rect 39264 16464 39270 16476
rect 39850 16464 39856 16476
rect 39908 16464 39914 16516
rect 7009 16439 7067 16445
rect 7009 16405 7021 16439
rect 7055 16436 7067 16439
rect 7374 16436 7380 16448
rect 7055 16408 7380 16436
rect 7055 16405 7067 16408
rect 7009 16399 7067 16405
rect 7374 16396 7380 16408
rect 7432 16396 7438 16448
rect 10410 16436 10416 16448
rect 10371 16408 10416 16436
rect 10410 16396 10416 16408
rect 10468 16396 10474 16448
rect 12710 16396 12716 16448
rect 12768 16436 12774 16448
rect 13173 16439 13231 16445
rect 13173 16436 13185 16439
rect 12768 16408 13185 16436
rect 12768 16396 12774 16408
rect 13173 16405 13185 16408
rect 13219 16405 13231 16439
rect 15378 16436 15384 16448
rect 15339 16408 15384 16436
rect 13173 16399 13231 16405
rect 15378 16396 15384 16408
rect 15436 16396 15442 16448
rect 17126 16436 17132 16448
rect 17087 16408 17132 16436
rect 17126 16396 17132 16408
rect 17184 16396 17190 16448
rect 18233 16439 18291 16445
rect 18233 16405 18245 16439
rect 18279 16436 18291 16439
rect 18414 16436 18420 16448
rect 18279 16408 18420 16436
rect 18279 16405 18291 16408
rect 18233 16399 18291 16405
rect 18414 16396 18420 16408
rect 18472 16396 18478 16448
rect 19245 16439 19303 16445
rect 19245 16405 19257 16439
rect 19291 16436 19303 16439
rect 19426 16436 19432 16448
rect 19291 16408 19432 16436
rect 19291 16405 19303 16408
rect 19245 16399 19303 16405
rect 19426 16396 19432 16408
rect 19484 16396 19490 16448
rect 30006 16396 30012 16448
rect 30064 16436 30070 16448
rect 31021 16439 31079 16445
rect 31021 16436 31033 16439
rect 30064 16408 31033 16436
rect 30064 16396 30070 16408
rect 31021 16405 31033 16408
rect 31067 16405 31079 16439
rect 31021 16399 31079 16405
rect 35621 16439 35679 16445
rect 35621 16405 35633 16439
rect 35667 16436 35679 16439
rect 35894 16436 35900 16448
rect 35667 16408 35900 16436
rect 35667 16405 35679 16408
rect 35621 16399 35679 16405
rect 35894 16396 35900 16408
rect 35952 16396 35958 16448
rect 36814 16436 36820 16448
rect 36775 16408 36820 16436
rect 36814 16396 36820 16408
rect 36872 16396 36878 16448
rect 38194 16396 38200 16448
rect 38252 16436 38258 16448
rect 39868 16436 39896 16464
rect 38252 16408 39896 16436
rect 40221 16439 40279 16445
rect 38252 16396 38258 16408
rect 40221 16405 40233 16439
rect 40267 16436 40279 16439
rect 40310 16436 40316 16448
rect 40267 16408 40316 16436
rect 40267 16405 40279 16408
rect 40221 16399 40279 16405
rect 40310 16396 40316 16408
rect 40368 16396 40374 16448
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 10045 16235 10103 16241
rect 10045 16201 10057 16235
rect 10091 16232 10103 16235
rect 10134 16232 10140 16244
rect 10091 16204 10140 16232
rect 10091 16201 10103 16204
rect 10045 16195 10103 16201
rect 10134 16192 10140 16204
rect 10192 16192 10198 16244
rect 10689 16235 10747 16241
rect 10689 16201 10701 16235
rect 10735 16232 10747 16235
rect 11146 16232 11152 16244
rect 10735 16204 11152 16232
rect 10735 16201 10747 16204
rect 10689 16195 10747 16201
rect 11146 16192 11152 16204
rect 11204 16192 11210 16244
rect 12158 16232 12164 16244
rect 12119 16204 12164 16232
rect 12158 16192 12164 16204
rect 12216 16192 12222 16244
rect 12434 16192 12440 16244
rect 12492 16232 12498 16244
rect 12713 16235 12771 16241
rect 12713 16232 12725 16235
rect 12492 16204 12725 16232
rect 12492 16192 12498 16204
rect 12713 16201 12725 16204
rect 12759 16201 12771 16235
rect 12713 16195 12771 16201
rect 15838 16192 15844 16244
rect 15896 16232 15902 16244
rect 16761 16235 16819 16241
rect 16761 16232 16773 16235
rect 15896 16204 16773 16232
rect 15896 16192 15902 16204
rect 16761 16201 16773 16204
rect 16807 16201 16819 16235
rect 16761 16195 16819 16201
rect 17310 16192 17316 16244
rect 17368 16232 17374 16244
rect 17589 16235 17647 16241
rect 17589 16232 17601 16235
rect 17368 16204 17601 16232
rect 17368 16192 17374 16204
rect 17589 16201 17601 16204
rect 17635 16201 17647 16235
rect 17589 16195 17647 16201
rect 17770 16192 17776 16244
rect 17828 16232 17834 16244
rect 18785 16235 18843 16241
rect 18785 16232 18797 16235
rect 17828 16204 18797 16232
rect 17828 16192 17834 16204
rect 18785 16201 18797 16204
rect 18831 16201 18843 16235
rect 18785 16195 18843 16201
rect 20717 16235 20775 16241
rect 20717 16201 20729 16235
rect 20763 16232 20775 16235
rect 20806 16232 20812 16244
rect 20763 16204 20812 16232
rect 20763 16201 20775 16204
rect 20717 16195 20775 16201
rect 20806 16192 20812 16204
rect 20864 16192 20870 16244
rect 22465 16235 22523 16241
rect 22465 16201 22477 16235
rect 22511 16232 22523 16235
rect 23106 16232 23112 16244
rect 22511 16204 23112 16232
rect 22511 16201 22523 16204
rect 22465 16195 22523 16201
rect 23106 16192 23112 16204
rect 23164 16192 23170 16244
rect 23382 16192 23388 16244
rect 23440 16232 23446 16244
rect 25041 16235 25099 16241
rect 23440 16204 23612 16232
rect 23440 16192 23446 16204
rect 3697 16167 3755 16173
rect 3697 16133 3709 16167
rect 3743 16164 3755 16167
rect 3786 16164 3792 16176
rect 3743 16136 3792 16164
rect 3743 16133 3755 16136
rect 3697 16127 3755 16133
rect 3786 16124 3792 16136
rect 3844 16124 3850 16176
rect 10410 16164 10416 16176
rect 9968 16136 10416 16164
rect 2130 16056 2136 16108
rect 2188 16096 2194 16108
rect 9968 16105 9996 16136
rect 10410 16124 10416 16136
rect 10468 16164 10474 16176
rect 10468 16136 10640 16164
rect 10468 16124 10474 16136
rect 2225 16099 2283 16105
rect 2225 16096 2237 16099
rect 2188 16068 2237 16096
rect 2188 16056 2194 16068
rect 2225 16065 2237 16068
rect 2271 16065 2283 16099
rect 2225 16059 2283 16065
rect 3605 16099 3663 16105
rect 3605 16065 3617 16099
rect 3651 16065 3663 16099
rect 9953 16099 10011 16105
rect 9953 16096 9965 16099
rect 3605 16059 3663 16065
rect 9416 16068 9965 16096
rect 1765 15963 1823 15969
rect 1765 15929 1777 15963
rect 1811 15960 1823 15963
rect 3620 15960 3648 16059
rect 3881 16031 3939 16037
rect 3881 15997 3893 16031
rect 3927 16028 3939 16031
rect 4614 16028 4620 16040
rect 3927 16000 4620 16028
rect 3927 15997 3939 16000
rect 3881 15991 3939 15997
rect 4614 15988 4620 16000
rect 4672 16028 4678 16040
rect 5350 16028 5356 16040
rect 4672 16000 5356 16028
rect 4672 15988 4678 16000
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 1811 15932 3648 15960
rect 1811 15929 1823 15932
rect 1765 15923 1823 15929
rect 2409 15895 2467 15901
rect 2409 15861 2421 15895
rect 2455 15892 2467 15895
rect 2498 15892 2504 15904
rect 2455 15864 2504 15892
rect 2455 15861 2467 15864
rect 2409 15855 2467 15861
rect 2498 15852 2504 15864
rect 2556 15852 2562 15904
rect 2590 15852 2596 15904
rect 2648 15892 2654 15904
rect 3237 15895 3295 15901
rect 3237 15892 3249 15895
rect 2648 15864 3249 15892
rect 2648 15852 2654 15864
rect 3237 15861 3249 15864
rect 3283 15861 3295 15895
rect 3620 15892 3648 15932
rect 4525 15895 4583 15901
rect 4525 15892 4537 15895
rect 3620 15864 4537 15892
rect 3237 15855 3295 15861
rect 4525 15861 4537 15864
rect 4571 15892 4583 15895
rect 5994 15892 6000 15904
rect 4571 15864 6000 15892
rect 4571 15861 4583 15864
rect 4525 15855 4583 15861
rect 5994 15852 6000 15864
rect 6052 15852 6058 15904
rect 6546 15852 6552 15904
rect 6604 15892 6610 15904
rect 7653 15895 7711 15901
rect 7653 15892 7665 15895
rect 6604 15864 7665 15892
rect 6604 15852 6610 15864
rect 7653 15861 7665 15864
rect 7699 15861 7711 15895
rect 7653 15855 7711 15861
rect 8662 15852 8668 15904
rect 8720 15892 8726 15904
rect 9416 15901 9444 16068
rect 9953 16065 9965 16068
rect 9999 16065 10011 16099
rect 9953 16059 10011 16065
rect 10137 16099 10195 16105
rect 10137 16065 10149 16099
rect 10183 16096 10195 16099
rect 10226 16096 10232 16108
rect 10183 16068 10232 16096
rect 10183 16065 10195 16068
rect 10137 16059 10195 16065
rect 10226 16056 10232 16068
rect 10284 16056 10290 16108
rect 10612 16105 10640 16136
rect 11238 16124 11244 16176
rect 11296 16164 11302 16176
rect 11793 16167 11851 16173
rect 11793 16164 11805 16167
rect 11296 16136 11805 16164
rect 11296 16124 11302 16136
rect 11793 16133 11805 16136
rect 11839 16133 11851 16167
rect 11793 16127 11851 16133
rect 11885 16167 11943 16173
rect 11885 16133 11897 16167
rect 11931 16164 11943 16167
rect 13354 16164 13360 16176
rect 11931 16136 13360 16164
rect 11931 16133 11943 16136
rect 11885 16127 11943 16133
rect 10597 16099 10655 16105
rect 10597 16065 10609 16099
rect 10643 16065 10655 16099
rect 10597 16059 10655 16065
rect 10781 16099 10839 16105
rect 10781 16065 10793 16099
rect 10827 16096 10839 16099
rect 10962 16096 10968 16108
rect 10827 16068 10968 16096
rect 10827 16065 10839 16068
rect 10781 16059 10839 16065
rect 9401 15895 9459 15901
rect 9401 15892 9413 15895
rect 8720 15864 9413 15892
rect 8720 15852 8726 15864
rect 9401 15861 9413 15864
rect 9447 15861 9459 15895
rect 10612 15892 10640 16059
rect 10962 16056 10968 16068
rect 11020 16056 11026 16108
rect 11514 16096 11520 16108
rect 11475 16068 11520 16096
rect 11514 16056 11520 16068
rect 11572 16056 11578 16108
rect 11606 16056 11612 16108
rect 11664 16096 11670 16108
rect 11664 16068 11709 16096
rect 11664 16056 11670 16068
rect 11808 16028 11836 16127
rect 13354 16124 13360 16136
rect 13412 16124 13418 16176
rect 17129 16167 17187 16173
rect 17129 16133 17141 16167
rect 17175 16164 17187 16167
rect 17954 16164 17960 16176
rect 17175 16136 17960 16164
rect 17175 16133 17187 16136
rect 17129 16127 17187 16133
rect 17954 16124 17960 16136
rect 18012 16124 18018 16176
rect 18969 16167 19027 16173
rect 18969 16133 18981 16167
rect 19015 16164 19027 16167
rect 23474 16164 23480 16176
rect 19015 16136 19334 16164
rect 19015 16133 19027 16136
rect 18969 16127 19027 16133
rect 11974 16056 11980 16108
rect 12032 16105 12038 16108
rect 12032 16096 12040 16105
rect 12621 16099 12679 16105
rect 12032 16068 12077 16096
rect 12406 16068 12572 16096
rect 12032 16059 12040 16068
rect 12032 16056 12038 16059
rect 12406 16028 12434 16068
rect 11808 16000 12434 16028
rect 12544 16028 12572 16068
rect 12621 16065 12633 16099
rect 12667 16096 12679 16099
rect 12710 16096 12716 16108
rect 12667 16068 12716 16096
rect 12667 16065 12679 16068
rect 12621 16059 12679 16065
rect 12710 16056 12716 16068
rect 12768 16056 12774 16108
rect 12805 16099 12863 16105
rect 12805 16065 12817 16099
rect 12851 16096 12863 16099
rect 12986 16096 12992 16108
rect 12851 16068 12992 16096
rect 12851 16065 12863 16068
rect 12805 16059 12863 16065
rect 12986 16056 12992 16068
rect 13044 16056 13050 16108
rect 14274 16096 14280 16108
rect 14187 16068 14280 16096
rect 14274 16056 14280 16068
rect 14332 16096 14338 16108
rect 14918 16096 14924 16108
rect 14332 16068 14924 16096
rect 14332 16056 14338 16068
rect 14918 16056 14924 16068
rect 14976 16056 14982 16108
rect 16850 16056 16856 16108
rect 16908 16096 16914 16108
rect 16945 16099 17003 16105
rect 16945 16096 16957 16099
rect 16908 16068 16957 16096
rect 16908 16056 16914 16068
rect 16945 16065 16957 16068
rect 16991 16065 17003 16099
rect 16945 16059 17003 16065
rect 17773 16099 17831 16105
rect 17773 16065 17785 16099
rect 17819 16065 17831 16099
rect 17972 16096 18000 16124
rect 19153 16099 19211 16105
rect 19153 16096 19165 16099
rect 17972 16068 19165 16096
rect 17773 16059 17831 16065
rect 19153 16065 19165 16068
rect 19199 16065 19211 16099
rect 19306 16096 19334 16136
rect 22572 16136 23480 16164
rect 19426 16096 19432 16108
rect 19306 16068 19432 16096
rect 19153 16059 19211 16065
rect 12894 16028 12900 16040
rect 12544 16000 12900 16028
rect 12894 15988 12900 16000
rect 12952 16028 12958 16040
rect 14550 16028 14556 16040
rect 12952 16000 14556 16028
rect 12952 15988 12958 16000
rect 14550 15988 14556 16000
rect 14608 15988 14614 16040
rect 17788 16028 17816 16059
rect 19426 16056 19432 16068
rect 19484 16056 19490 16108
rect 20625 16099 20683 16105
rect 20625 16096 20637 16099
rect 20088 16068 20637 16096
rect 18230 16028 18236 16040
rect 17788 16000 18236 16028
rect 18230 15988 18236 16000
rect 18288 15988 18294 16040
rect 12710 15920 12716 15972
rect 12768 15960 12774 15972
rect 19886 15960 19892 15972
rect 12768 15932 19892 15960
rect 12768 15920 12774 15932
rect 19886 15920 19892 15932
rect 19944 15960 19950 15972
rect 20088 15969 20116 16068
rect 20625 16065 20637 16068
rect 20671 16065 20683 16099
rect 20806 16096 20812 16108
rect 20767 16068 20812 16096
rect 20625 16059 20683 16065
rect 20806 16056 20812 16068
rect 20864 16056 20870 16108
rect 22094 16056 22100 16108
rect 22152 16096 22158 16108
rect 22572 16105 22600 16136
rect 23474 16124 23480 16136
rect 23532 16124 23538 16176
rect 23584 16164 23612 16204
rect 25041 16201 25053 16235
rect 25087 16232 25099 16235
rect 25498 16232 25504 16244
rect 25087 16204 25504 16232
rect 25087 16201 25099 16204
rect 25041 16195 25099 16201
rect 25498 16192 25504 16204
rect 25556 16192 25562 16244
rect 26053 16235 26111 16241
rect 26053 16201 26065 16235
rect 26099 16232 26111 16235
rect 26326 16232 26332 16244
rect 26099 16204 26332 16232
rect 26099 16201 26111 16204
rect 26053 16195 26111 16201
rect 26326 16192 26332 16204
rect 26384 16192 26390 16244
rect 26602 16192 26608 16244
rect 26660 16232 26666 16244
rect 28902 16232 28908 16244
rect 26660 16204 27568 16232
rect 28863 16204 28908 16232
rect 26660 16192 26666 16204
rect 26234 16164 26240 16176
rect 23584 16136 25636 16164
rect 26195 16136 26240 16164
rect 22373 16099 22431 16105
rect 22373 16096 22385 16099
rect 22152 16068 22385 16096
rect 22152 16056 22158 16068
rect 22373 16065 22385 16068
rect 22419 16065 22431 16099
rect 22373 16059 22431 16065
rect 22557 16099 22615 16105
rect 22557 16065 22569 16099
rect 22603 16065 22615 16099
rect 22557 16059 22615 16065
rect 23201 16099 23259 16105
rect 23201 16065 23213 16099
rect 23247 16096 23259 16099
rect 23658 16096 23664 16108
rect 23247 16068 23664 16096
rect 23247 16065 23259 16068
rect 23201 16059 23259 16065
rect 20073 15963 20131 15969
rect 20073 15960 20085 15963
rect 19944 15932 20085 15960
rect 19944 15920 19950 15932
rect 20073 15929 20085 15932
rect 20119 15929 20131 15963
rect 20073 15923 20131 15929
rect 13814 15892 13820 15904
rect 10612 15864 13820 15892
rect 9401 15855 9459 15861
rect 13814 15852 13820 15864
rect 13872 15852 13878 15904
rect 20346 15852 20352 15904
rect 20404 15892 20410 15904
rect 21821 15895 21879 15901
rect 21821 15892 21833 15895
rect 20404 15864 21833 15892
rect 20404 15852 20410 15864
rect 21821 15861 21833 15864
rect 21867 15892 21879 15895
rect 22572 15892 22600 16059
rect 23658 16056 23664 16068
rect 23716 16056 23722 16108
rect 25608 16105 25636 16136
rect 26234 16124 26240 16136
rect 26292 16124 26298 16176
rect 26421 16167 26479 16173
rect 26421 16133 26433 16167
rect 26467 16164 26479 16167
rect 27430 16164 27436 16176
rect 26467 16136 27436 16164
rect 26467 16133 26479 16136
rect 26421 16127 26479 16133
rect 27430 16124 27436 16136
rect 27488 16124 27494 16176
rect 27540 16164 27568 16204
rect 28902 16192 28908 16204
rect 28960 16192 28966 16244
rect 33594 16192 33600 16244
rect 33652 16232 33658 16244
rect 33781 16235 33839 16241
rect 33781 16232 33793 16235
rect 33652 16204 33793 16232
rect 33652 16192 33658 16204
rect 33781 16201 33793 16204
rect 33827 16201 33839 16235
rect 40218 16232 40224 16244
rect 40179 16204 40224 16232
rect 33781 16195 33839 16201
rect 40218 16192 40224 16204
rect 40276 16192 40282 16244
rect 38286 16164 38292 16176
rect 27540 16136 38292 16164
rect 38286 16124 38292 16136
rect 38344 16124 38350 16176
rect 39298 16164 39304 16176
rect 38856 16136 39304 16164
rect 25593 16099 25651 16105
rect 25593 16065 25605 16099
rect 25639 16096 25651 16099
rect 26602 16096 26608 16108
rect 25639 16068 26608 16096
rect 25639 16065 25651 16068
rect 25593 16059 25651 16065
rect 26602 16056 26608 16068
rect 26660 16056 26666 16108
rect 29181 16099 29239 16105
rect 29181 16096 29193 16099
rect 28368 16068 29193 16096
rect 23477 16031 23535 16037
rect 23477 15997 23489 16031
rect 23523 16028 23535 16031
rect 23566 16028 23572 16040
rect 23523 16000 23572 16028
rect 23523 15997 23535 16000
rect 23477 15991 23535 15997
rect 23566 15988 23572 16000
rect 23624 16028 23630 16040
rect 27522 16028 27528 16040
rect 23624 16000 27528 16028
rect 23624 15988 23630 16000
rect 27522 15988 27528 16000
rect 27580 15988 27586 16040
rect 27246 15892 27252 15904
rect 21867 15864 22600 15892
rect 27207 15864 27252 15892
rect 21867 15861 21879 15864
rect 21821 15855 21879 15861
rect 27246 15852 27252 15864
rect 27304 15852 27310 15904
rect 27890 15852 27896 15904
rect 27948 15892 27954 15904
rect 28368 15901 28396 16068
rect 29181 16065 29193 16068
rect 29227 16065 29239 16099
rect 29181 16059 29239 16065
rect 29273 16099 29331 16105
rect 29273 16065 29285 16099
rect 29319 16065 29331 16099
rect 29273 16059 29331 16065
rect 29288 15960 29316 16059
rect 29362 16056 29368 16108
rect 29420 16096 29426 16108
rect 29549 16099 29607 16105
rect 29420 16068 29465 16096
rect 29420 16056 29426 16068
rect 29549 16065 29561 16099
rect 29595 16096 29607 16099
rect 30190 16096 30196 16108
rect 29595 16068 30196 16096
rect 29595 16065 29607 16068
rect 29549 16059 29607 16065
rect 30190 16056 30196 16068
rect 30248 16056 30254 16108
rect 31294 16096 31300 16108
rect 31255 16068 31300 16096
rect 31294 16056 31300 16068
rect 31352 16056 31358 16108
rect 32490 16096 32496 16108
rect 32451 16068 32496 16096
rect 32490 16056 32496 16068
rect 32548 16056 32554 16108
rect 35529 16099 35587 16105
rect 35529 16065 35541 16099
rect 35575 16096 35587 16099
rect 37182 16096 37188 16108
rect 35575 16068 37188 16096
rect 35575 16065 35587 16068
rect 35529 16059 35587 16065
rect 37182 16056 37188 16068
rect 37240 16056 37246 16108
rect 38856 16105 38884 16136
rect 39298 16124 39304 16136
rect 39356 16124 39362 16176
rect 38841 16099 38899 16105
rect 38841 16065 38853 16099
rect 38887 16065 38899 16099
rect 38841 16059 38899 16065
rect 39108 16099 39166 16105
rect 39108 16065 39120 16099
rect 39154 16096 39166 16099
rect 39850 16096 39856 16108
rect 39154 16068 39856 16096
rect 39154 16065 39166 16068
rect 39108 16059 39166 16065
rect 39850 16056 39856 16068
rect 39908 16056 39914 16108
rect 40957 16099 41015 16105
rect 40957 16065 40969 16099
rect 41003 16096 41015 16099
rect 41138 16096 41144 16108
rect 41003 16068 41144 16096
rect 41003 16065 41015 16068
rect 40957 16059 41015 16065
rect 41138 16056 41144 16068
rect 41196 16056 41202 16108
rect 30006 16028 30012 16040
rect 29967 16000 30012 16028
rect 30006 15988 30012 16000
rect 30064 15988 30070 16040
rect 30098 15988 30104 16040
rect 30156 16028 30162 16040
rect 30285 16031 30343 16037
rect 30285 16028 30297 16031
rect 30156 16000 30297 16028
rect 30156 15988 30162 16000
rect 30285 15997 30297 16000
rect 30331 15997 30343 16031
rect 30285 15991 30343 15997
rect 35253 16031 35311 16037
rect 35253 15997 35265 16031
rect 35299 16028 35311 16031
rect 35342 16028 35348 16040
rect 35299 16000 35348 16028
rect 35299 15997 35311 16000
rect 35253 15991 35311 15997
rect 35342 15988 35348 16000
rect 35400 15988 35406 16040
rect 40678 16028 40684 16040
rect 40639 16000 40684 16028
rect 40678 15988 40684 16000
rect 40736 15988 40742 16040
rect 30116 15960 30144 15988
rect 29288 15932 30144 15960
rect 28353 15895 28411 15901
rect 28353 15892 28365 15895
rect 27948 15864 28365 15892
rect 27948 15852 27954 15864
rect 28353 15861 28365 15864
rect 28399 15861 28411 15895
rect 28353 15855 28411 15861
rect 31386 15852 31392 15904
rect 31444 15892 31450 15904
rect 31481 15895 31539 15901
rect 31481 15892 31493 15895
rect 31444 15864 31493 15892
rect 31444 15852 31450 15864
rect 31481 15861 31493 15864
rect 31527 15861 31539 15895
rect 58158 15892 58164 15904
rect 58119 15864 58164 15892
rect 31481 15855 31539 15861
rect 58158 15852 58164 15864
rect 58216 15852 58222 15904
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 2130 15688 2136 15700
rect 2091 15660 2136 15688
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 7558 15688 7564 15700
rect 7519 15660 7564 15688
rect 7558 15648 7564 15660
rect 7616 15648 7622 15700
rect 8389 15691 8447 15697
rect 8389 15657 8401 15691
rect 8435 15688 8447 15691
rect 8478 15688 8484 15700
rect 8435 15660 8484 15688
rect 8435 15657 8447 15660
rect 8389 15651 8447 15657
rect 8478 15648 8484 15660
rect 8536 15648 8542 15700
rect 10226 15688 10232 15700
rect 10187 15660 10232 15688
rect 10226 15648 10232 15660
rect 10284 15648 10290 15700
rect 12161 15691 12219 15697
rect 12161 15657 12173 15691
rect 12207 15688 12219 15691
rect 12526 15688 12532 15700
rect 12207 15660 12532 15688
rect 12207 15657 12219 15660
rect 12161 15651 12219 15657
rect 12526 15648 12532 15660
rect 12584 15648 12590 15700
rect 14274 15688 14280 15700
rect 14235 15660 14280 15688
rect 14274 15648 14280 15660
rect 14332 15648 14338 15700
rect 15120 15660 17172 15688
rect 15120 15620 15148 15660
rect 13740 15592 15148 15620
rect 2590 15552 2596 15564
rect 2332 15524 2596 15552
rect 2332 15493 2360 15524
rect 2590 15512 2596 15524
rect 2648 15512 2654 15564
rect 2774 15512 2780 15564
rect 2832 15552 2838 15564
rect 3789 15555 3847 15561
rect 3789 15552 3801 15555
rect 2832 15524 3801 15552
rect 2832 15512 2838 15524
rect 3789 15521 3801 15524
rect 3835 15521 3847 15555
rect 3789 15515 3847 15521
rect 6273 15555 6331 15561
rect 6273 15521 6285 15555
rect 6319 15552 6331 15555
rect 7101 15555 7159 15561
rect 7101 15552 7113 15555
rect 6319 15524 7113 15552
rect 6319 15521 6331 15524
rect 6273 15515 6331 15521
rect 7101 15521 7113 15524
rect 7147 15521 7159 15555
rect 7101 15515 7159 15521
rect 7193 15555 7251 15561
rect 7193 15521 7205 15555
rect 7239 15552 7251 15555
rect 7282 15552 7288 15564
rect 7239 15524 7288 15552
rect 7239 15521 7251 15524
rect 7193 15515 7251 15521
rect 7282 15512 7288 15524
rect 7340 15512 7346 15564
rect 2317 15487 2375 15493
rect 2317 15453 2329 15487
rect 2363 15453 2375 15487
rect 2317 15447 2375 15453
rect 2406 15444 2412 15496
rect 2464 15484 2470 15496
rect 3053 15487 3111 15493
rect 2464 15456 2509 15484
rect 2464 15444 2470 15456
rect 3053 15453 3065 15487
rect 3099 15484 3111 15487
rect 5997 15487 6055 15493
rect 5997 15484 6009 15487
rect 3099 15456 4200 15484
rect 3099 15453 3111 15456
rect 3053 15447 3111 15453
rect 4034 15419 4092 15425
rect 4034 15416 4046 15419
rect 3252 15388 4046 15416
rect 3252 15357 3280 15388
rect 4034 15385 4046 15388
rect 4080 15385 4092 15419
rect 4172 15416 4200 15456
rect 4356 15456 6009 15484
rect 4246 15416 4252 15428
rect 4172 15388 4252 15416
rect 4034 15379 4092 15385
rect 4246 15376 4252 15388
rect 4304 15376 4310 15428
rect 3237 15351 3295 15357
rect 3237 15317 3249 15351
rect 3283 15317 3295 15351
rect 3237 15311 3295 15317
rect 3786 15308 3792 15360
rect 3844 15348 3850 15360
rect 4356 15348 4384 15456
rect 5997 15453 6009 15456
rect 6043 15453 6055 15487
rect 5997 15447 6055 15453
rect 6086 15444 6092 15496
rect 6144 15484 6150 15496
rect 6638 15484 6644 15496
rect 6144 15456 6644 15484
rect 6144 15444 6150 15456
rect 6638 15444 6644 15456
rect 6696 15444 6702 15496
rect 6825 15487 6883 15493
rect 6825 15453 6837 15487
rect 6871 15453 6883 15487
rect 7006 15484 7012 15496
rect 6967 15456 7012 15484
rect 6825 15447 6883 15453
rect 6546 15376 6552 15428
rect 6604 15416 6610 15428
rect 6840 15416 6868 15447
rect 7006 15444 7012 15456
rect 7064 15444 7070 15496
rect 7374 15484 7380 15496
rect 7335 15456 7380 15484
rect 7374 15444 7380 15456
rect 7432 15444 7438 15496
rect 8294 15484 8300 15496
rect 8255 15456 8300 15484
rect 8294 15444 8300 15456
rect 8352 15444 8358 15496
rect 8389 15487 8447 15493
rect 8389 15453 8401 15487
rect 8435 15484 8447 15487
rect 9858 15484 9864 15496
rect 8435 15456 9864 15484
rect 8435 15453 8447 15456
rect 8389 15447 8447 15453
rect 9858 15444 9864 15456
rect 9916 15444 9922 15496
rect 10870 15444 10876 15496
rect 10928 15484 10934 15496
rect 12066 15484 12072 15496
rect 10928 15456 12072 15484
rect 10928 15444 10934 15456
rect 12066 15444 12072 15456
rect 12124 15484 12130 15496
rect 13541 15487 13599 15493
rect 13541 15484 13553 15487
rect 12124 15456 13553 15484
rect 12124 15444 12130 15456
rect 13541 15453 13553 15456
rect 13587 15484 13599 15487
rect 13630 15484 13636 15496
rect 13587 15456 13636 15484
rect 13587 15453 13599 15456
rect 13541 15447 13599 15453
rect 13630 15444 13636 15456
rect 13688 15444 13694 15496
rect 6604 15388 6868 15416
rect 6604 15376 6610 15388
rect 12802 15376 12808 15428
rect 12860 15416 12866 15428
rect 13274 15419 13332 15425
rect 13274 15416 13286 15419
rect 12860 15388 13286 15416
rect 12860 15376 12866 15388
rect 13274 15385 13286 15388
rect 13320 15385 13332 15419
rect 13274 15379 13332 15385
rect 3844 15320 4384 15348
rect 3844 15308 3850 15320
rect 5074 15308 5080 15360
rect 5132 15348 5138 15360
rect 5169 15351 5227 15357
rect 5169 15348 5181 15351
rect 5132 15320 5181 15348
rect 5132 15308 5138 15320
rect 5169 15317 5181 15320
rect 5215 15317 5227 15351
rect 5626 15348 5632 15360
rect 5587 15320 5632 15348
rect 5169 15311 5227 15317
rect 5626 15308 5632 15320
rect 5684 15308 5690 15360
rect 6822 15308 6828 15360
rect 6880 15348 6886 15360
rect 8021 15351 8079 15357
rect 8021 15348 8033 15351
rect 6880 15320 8033 15348
rect 6880 15308 6886 15320
rect 8021 15317 8033 15320
rect 8067 15317 8079 15351
rect 10962 15348 10968 15360
rect 10923 15320 10968 15348
rect 8021 15311 8079 15317
rect 10962 15308 10968 15320
rect 11020 15308 11026 15360
rect 12986 15308 12992 15360
rect 13044 15348 13050 15360
rect 13740 15348 13768 15592
rect 13814 15512 13820 15564
rect 13872 15552 13878 15564
rect 13872 15524 14320 15552
rect 13872 15512 13878 15524
rect 13998 15444 14004 15496
rect 14056 15484 14062 15496
rect 14292 15493 14320 15524
rect 14093 15487 14151 15493
rect 14093 15484 14105 15487
rect 14056 15456 14105 15484
rect 14056 15444 14062 15456
rect 14093 15453 14105 15456
rect 14139 15453 14151 15487
rect 14093 15447 14151 15453
rect 14277 15487 14335 15493
rect 14277 15453 14289 15487
rect 14323 15453 14335 15487
rect 15102 15484 15108 15496
rect 15063 15456 15108 15484
rect 14277 15447 14335 15453
rect 14292 15416 14320 15447
rect 15102 15444 15108 15456
rect 15160 15444 15166 15496
rect 15378 15493 15384 15496
rect 15372 15484 15384 15493
rect 15339 15456 15384 15484
rect 15372 15447 15384 15456
rect 15378 15444 15384 15447
rect 15436 15444 15442 15496
rect 17144 15484 17172 15660
rect 19334 15648 19340 15700
rect 19392 15688 19398 15700
rect 19429 15691 19487 15697
rect 19429 15688 19441 15691
rect 19392 15660 19441 15688
rect 19392 15648 19398 15660
rect 19429 15657 19441 15660
rect 19475 15657 19487 15691
rect 19886 15688 19892 15700
rect 19847 15660 19892 15688
rect 19429 15651 19487 15657
rect 19886 15648 19892 15660
rect 19944 15648 19950 15700
rect 22094 15648 22100 15700
rect 22152 15688 22158 15700
rect 22741 15691 22799 15697
rect 22152 15660 22197 15688
rect 22152 15648 22158 15660
rect 22741 15657 22753 15691
rect 22787 15688 22799 15691
rect 23658 15688 23664 15700
rect 22787 15660 23664 15688
rect 22787 15657 22799 15660
rect 22741 15651 22799 15657
rect 23658 15648 23664 15660
rect 23716 15648 23722 15700
rect 26694 15648 26700 15700
rect 26752 15688 26758 15700
rect 27433 15691 27491 15697
rect 27433 15688 27445 15691
rect 26752 15660 27445 15688
rect 26752 15648 26758 15660
rect 27433 15657 27445 15660
rect 27479 15688 27491 15691
rect 29914 15688 29920 15700
rect 27479 15660 29920 15688
rect 27479 15657 27491 15660
rect 27433 15651 27491 15657
rect 29914 15648 29920 15660
rect 29972 15648 29978 15700
rect 30929 15691 30987 15697
rect 30929 15657 30941 15691
rect 30975 15688 30987 15691
rect 31202 15688 31208 15700
rect 30975 15660 31208 15688
rect 30975 15657 30987 15660
rect 30929 15651 30987 15657
rect 31202 15648 31208 15660
rect 31260 15648 31266 15700
rect 38286 15688 38292 15700
rect 38247 15660 38292 15688
rect 38286 15648 38292 15660
rect 38344 15648 38350 15700
rect 39850 15688 39856 15700
rect 39811 15660 39856 15688
rect 39850 15648 39856 15660
rect 39908 15648 39914 15700
rect 18690 15552 18696 15564
rect 18651 15524 18696 15552
rect 18690 15512 18696 15524
rect 18748 15512 18754 15564
rect 19518 15552 19524 15564
rect 19260 15524 19524 15552
rect 19260 15493 19288 15524
rect 19518 15512 19524 15524
rect 19576 15512 19582 15564
rect 19245 15487 19303 15493
rect 19245 15484 19257 15487
rect 15488 15456 17080 15484
rect 17144 15456 19257 15484
rect 15488 15416 15516 15456
rect 14292 15388 15516 15416
rect 16022 15376 16028 15428
rect 16080 15416 16086 15428
rect 16945 15419 17003 15425
rect 16945 15416 16957 15419
rect 16080 15388 16957 15416
rect 16080 15376 16086 15388
rect 16945 15385 16957 15388
rect 16991 15385 17003 15419
rect 17052 15416 17080 15456
rect 19245 15453 19257 15456
rect 19291 15453 19303 15487
rect 19245 15447 19303 15453
rect 19334 15444 19340 15496
rect 19392 15484 19398 15496
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 19392 15456 19441 15484
rect 19392 15444 19398 15456
rect 19429 15453 19441 15456
rect 19475 15453 19487 15487
rect 19904 15484 19932 15648
rect 20625 15623 20683 15629
rect 20625 15589 20637 15623
rect 20671 15620 20683 15623
rect 27062 15620 27068 15632
rect 20671 15592 27068 15620
rect 20671 15589 20683 15592
rect 20625 15583 20683 15589
rect 27062 15580 27068 15592
rect 27120 15580 27126 15632
rect 20254 15512 20260 15564
rect 20312 15552 20318 15564
rect 20312 15524 20668 15552
rect 20312 15512 20318 15524
rect 20640 15493 20668 15524
rect 34698 15512 34704 15564
rect 34756 15552 34762 15564
rect 35437 15555 35495 15561
rect 35437 15552 35449 15555
rect 34756 15524 35449 15552
rect 34756 15512 34762 15524
rect 35437 15521 35449 15524
rect 35483 15521 35495 15555
rect 35437 15515 35495 15521
rect 35713 15555 35771 15561
rect 35713 15521 35725 15555
rect 35759 15552 35771 15555
rect 36998 15552 37004 15564
rect 35759 15524 37004 15552
rect 35759 15521 35771 15524
rect 35713 15515 35771 15521
rect 36998 15512 37004 15524
rect 37056 15512 37062 15564
rect 39206 15512 39212 15564
rect 39264 15552 39270 15564
rect 39264 15524 40264 15552
rect 39264 15512 39270 15524
rect 20441 15487 20499 15493
rect 20441 15484 20453 15487
rect 19904 15456 20453 15484
rect 19429 15447 19487 15453
rect 20441 15453 20453 15456
rect 20487 15453 20499 15487
rect 20441 15447 20499 15453
rect 20625 15487 20683 15493
rect 20625 15453 20637 15487
rect 20671 15453 20683 15487
rect 20625 15447 20683 15453
rect 20806 15444 20812 15496
rect 20864 15484 20870 15496
rect 21453 15487 21511 15493
rect 21453 15484 21465 15487
rect 20864 15456 21465 15484
rect 20864 15444 20870 15456
rect 21453 15453 21465 15456
rect 21499 15484 21511 15487
rect 21634 15484 21640 15496
rect 21499 15456 21640 15484
rect 21499 15453 21511 15456
rect 21453 15447 21511 15453
rect 21634 15444 21640 15456
rect 21692 15484 21698 15496
rect 22557 15487 22615 15493
rect 22557 15484 22569 15487
rect 21692 15456 22569 15484
rect 21692 15444 21698 15456
rect 22557 15453 22569 15456
rect 22603 15453 22615 15487
rect 22557 15447 22615 15453
rect 22741 15487 22799 15493
rect 22741 15453 22753 15487
rect 22787 15453 22799 15487
rect 22741 15447 22799 15453
rect 22094 15416 22100 15428
rect 17052 15388 22100 15416
rect 16945 15379 17003 15385
rect 22094 15376 22100 15388
rect 22152 15376 22158 15428
rect 22186 15376 22192 15428
rect 22244 15416 22250 15428
rect 22756 15416 22784 15447
rect 27062 15444 27068 15496
rect 27120 15484 27126 15496
rect 27341 15487 27399 15493
rect 27341 15484 27353 15487
rect 27120 15456 27353 15484
rect 27120 15444 27126 15456
rect 27341 15453 27353 15456
rect 27387 15453 27399 15487
rect 27522 15484 27528 15496
rect 27483 15456 27528 15484
rect 27341 15447 27399 15453
rect 23293 15419 23351 15425
rect 23293 15416 23305 15419
rect 22244 15388 23305 15416
rect 22244 15376 22250 15388
rect 23293 15385 23305 15388
rect 23339 15416 23351 15419
rect 23842 15416 23848 15428
rect 23339 15388 23848 15416
rect 23339 15385 23351 15388
rect 23293 15379 23351 15385
rect 23842 15376 23848 15388
rect 23900 15416 23906 15428
rect 24397 15419 24455 15425
rect 24397 15416 24409 15419
rect 23900 15388 24409 15416
rect 23900 15376 23906 15388
rect 24397 15385 24409 15388
rect 24443 15385 24455 15419
rect 27356 15416 27384 15447
rect 27522 15444 27528 15456
rect 27580 15444 27586 15496
rect 29546 15484 29552 15496
rect 29507 15456 29552 15484
rect 29546 15444 29552 15456
rect 29604 15444 29610 15496
rect 31202 15444 31208 15496
rect 31260 15484 31266 15496
rect 31573 15487 31631 15493
rect 31573 15484 31585 15487
rect 31260 15456 31585 15484
rect 31260 15444 31266 15456
rect 31573 15453 31585 15456
rect 31619 15453 31631 15487
rect 31573 15447 31631 15453
rect 33042 15444 33048 15496
rect 33100 15484 33106 15496
rect 33229 15487 33287 15493
rect 33229 15484 33241 15487
rect 33100 15456 33241 15484
rect 33100 15444 33106 15456
rect 33229 15453 33241 15456
rect 33275 15453 33287 15487
rect 33229 15447 33287 15453
rect 33505 15487 33563 15493
rect 33505 15453 33517 15487
rect 33551 15484 33563 15487
rect 33594 15484 33600 15496
rect 33551 15456 33600 15484
rect 33551 15453 33563 15456
rect 33505 15447 33563 15453
rect 27985 15419 28043 15425
rect 27985 15416 27997 15419
rect 27356 15388 27997 15416
rect 24397 15379 24455 15385
rect 27985 15385 27997 15388
rect 28031 15385 28043 15419
rect 27985 15379 28043 15385
rect 13044 15320 13768 15348
rect 16485 15351 16543 15357
rect 13044 15308 13050 15320
rect 16485 15317 16497 15351
rect 16531 15348 16543 15351
rect 16850 15348 16856 15360
rect 16531 15320 16856 15348
rect 16531 15317 16543 15320
rect 16485 15311 16543 15317
rect 16850 15308 16856 15320
rect 16908 15308 16914 15360
rect 19518 15308 19524 15360
rect 19576 15348 19582 15360
rect 21174 15348 21180 15360
rect 19576 15320 21180 15348
rect 19576 15308 19582 15320
rect 21174 15308 21180 15320
rect 21232 15308 21238 15360
rect 28000 15348 28028 15379
rect 29638 15376 29644 15428
rect 29696 15416 29702 15428
rect 29794 15419 29852 15425
rect 29794 15416 29806 15419
rect 29696 15388 29806 15416
rect 29696 15376 29702 15388
rect 29794 15385 29806 15388
rect 29840 15385 29852 15419
rect 31386 15416 31392 15428
rect 31347 15388 31392 15416
rect 29794 15379 29852 15385
rect 31386 15376 31392 15388
rect 31444 15376 31450 15428
rect 33244 15416 33272 15447
rect 33594 15444 33600 15456
rect 33652 15444 33658 15496
rect 37461 15487 37519 15493
rect 37461 15453 37473 15487
rect 37507 15484 37519 15487
rect 37734 15484 37740 15496
rect 37507 15456 37740 15484
rect 37507 15453 37519 15456
rect 37461 15447 37519 15453
rect 37734 15444 37740 15456
rect 37792 15484 37798 15496
rect 37918 15484 37924 15496
rect 37792 15456 37924 15484
rect 37792 15444 37798 15456
rect 37918 15444 37924 15456
rect 37976 15444 37982 15496
rect 38286 15444 38292 15496
rect 38344 15484 38350 15496
rect 40236 15493 40264 15524
rect 40129 15487 40187 15493
rect 40129 15484 40141 15487
rect 38344 15456 40141 15484
rect 38344 15444 38350 15456
rect 40129 15453 40141 15456
rect 40175 15453 40187 15487
rect 40129 15447 40187 15453
rect 40221 15487 40279 15493
rect 40221 15453 40233 15487
rect 40267 15453 40279 15487
rect 40221 15447 40279 15453
rect 34701 15419 34759 15425
rect 34701 15416 34713 15419
rect 33244 15388 34713 15416
rect 34701 15385 34713 15388
rect 34747 15385 34759 15419
rect 34701 15379 34759 15385
rect 37645 15419 37703 15425
rect 37645 15385 37657 15419
rect 37691 15416 37703 15419
rect 38654 15416 38660 15428
rect 37691 15388 38660 15416
rect 37691 15385 37703 15388
rect 37645 15379 37703 15385
rect 38654 15376 38660 15388
rect 38712 15376 38718 15428
rect 40144 15416 40172 15447
rect 40310 15444 40316 15496
rect 40368 15484 40374 15496
rect 40497 15487 40555 15493
rect 40368 15456 40413 15484
rect 40368 15444 40374 15456
rect 40497 15453 40509 15487
rect 40543 15484 40555 15487
rect 41138 15484 41144 15496
rect 40543 15456 41144 15484
rect 40543 15453 40555 15456
rect 40497 15447 40555 15453
rect 41138 15444 41144 15456
rect 41196 15444 41202 15496
rect 40957 15419 41015 15425
rect 40957 15416 40969 15419
rect 40144 15388 40969 15416
rect 40957 15385 40969 15388
rect 41003 15385 41015 15419
rect 40957 15379 41015 15385
rect 30006 15348 30012 15360
rect 28000 15320 30012 15348
rect 30006 15308 30012 15320
rect 30064 15308 30070 15360
rect 30190 15308 30196 15360
rect 30248 15348 30254 15360
rect 30466 15348 30472 15360
rect 30248 15320 30472 15348
rect 30248 15308 30254 15320
rect 30466 15308 30472 15320
rect 30524 15308 30530 15360
rect 31754 15348 31760 15360
rect 31715 15320 31760 15348
rect 31754 15308 31760 15320
rect 31812 15308 31818 15360
rect 32401 15351 32459 15357
rect 32401 15317 32413 15351
rect 32447 15348 32459 15351
rect 32490 15348 32496 15360
rect 32447 15320 32496 15348
rect 32447 15317 32459 15320
rect 32401 15311 32459 15317
rect 32490 15308 32496 15320
rect 32548 15308 32554 15360
rect 37829 15351 37887 15357
rect 37829 15317 37841 15351
rect 37875 15348 37887 15351
rect 37918 15348 37924 15360
rect 37875 15320 37924 15348
rect 37875 15317 37887 15320
rect 37829 15311 37887 15317
rect 37918 15308 37924 15320
rect 37976 15308 37982 15360
rect 38746 15308 38752 15360
rect 38804 15348 38810 15360
rect 38841 15351 38899 15357
rect 38841 15348 38853 15351
rect 38804 15320 38853 15348
rect 38804 15308 38810 15320
rect 38841 15317 38853 15320
rect 38887 15317 38899 15351
rect 38841 15311 38899 15317
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 3786 15144 3792 15156
rect 3747 15116 3792 15144
rect 3786 15104 3792 15116
rect 3844 15104 3850 15156
rect 4246 15144 4252 15156
rect 4207 15116 4252 15144
rect 4246 15104 4252 15116
rect 4304 15104 4310 15156
rect 7006 15144 7012 15156
rect 6967 15116 7012 15144
rect 7006 15104 7012 15116
rect 7064 15104 7070 15156
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 17218 15144 17224 15156
rect 8352 15116 17080 15144
rect 17179 15116 17224 15144
rect 8352 15104 8358 15116
rect 2774 15076 2780 15088
rect 2424 15048 2780 15076
rect 2424 15017 2452 15048
rect 2774 15036 2780 15048
rect 2832 15036 2838 15088
rect 3234 15036 3240 15088
rect 3292 15076 3298 15088
rect 6730 15076 6736 15088
rect 3292 15048 6736 15076
rect 3292 15036 3298 15048
rect 6730 15036 6736 15048
rect 6788 15036 6794 15088
rect 9490 15076 9496 15088
rect 9451 15048 9496 15076
rect 9490 15036 9496 15048
rect 9548 15036 9554 15088
rect 12526 15036 12532 15088
rect 12584 15076 12590 15088
rect 12584 15048 12756 15076
rect 12584 15036 12590 15048
rect 2409 15011 2467 15017
rect 2409 14977 2421 15011
rect 2455 14977 2467 15011
rect 2409 14971 2467 14977
rect 2498 14968 2504 15020
rect 2556 15008 2562 15020
rect 2665 15011 2723 15017
rect 2665 15008 2677 15011
rect 2556 14980 2677 15008
rect 2556 14968 2562 14980
rect 2665 14977 2677 14980
rect 2711 14977 2723 15011
rect 2665 14971 2723 14977
rect 4433 15011 4491 15017
rect 4433 14977 4445 15011
rect 4479 15008 4491 15011
rect 4706 15008 4712 15020
rect 4479 14980 4712 15008
rect 4479 14977 4491 14980
rect 4433 14971 4491 14977
rect 4706 14968 4712 14980
rect 4764 14968 4770 15020
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 14977 7435 15011
rect 7377 14971 7435 14977
rect 9401 15011 9459 15017
rect 9401 14977 9413 15011
rect 9447 14977 9459 15011
rect 9582 15008 9588 15020
rect 9543 14980 9588 15008
rect 9401 14971 9459 14977
rect 4617 14943 4675 14949
rect 4617 14909 4629 14943
rect 4663 14909 4675 14943
rect 4617 14903 4675 14909
rect 7285 14943 7343 14949
rect 7285 14909 7297 14943
rect 7331 14909 7343 14943
rect 7285 14903 7343 14909
rect 4632 14872 4660 14903
rect 3712 14844 4660 14872
rect 2406 14764 2412 14816
rect 2464 14804 2470 14816
rect 3712 14804 3740 14844
rect 2464 14776 3740 14804
rect 2464 14764 2470 14776
rect 5902 14764 5908 14816
rect 5960 14804 5966 14816
rect 7193 14807 7251 14813
rect 7193 14804 7205 14807
rect 5960 14776 7205 14804
rect 5960 14764 5966 14776
rect 7193 14773 7205 14776
rect 7239 14773 7251 14807
rect 7300 14804 7328 14903
rect 7392 14872 7420 14971
rect 9416 14940 9444 14971
rect 9582 14968 9588 14980
rect 9640 14968 9646 15020
rect 10413 15011 10471 15017
rect 10413 14977 10425 15011
rect 10459 15008 10471 15011
rect 12158 15008 12164 15020
rect 10459 14980 12164 15008
rect 10459 14977 10471 14980
rect 10413 14971 10471 14977
rect 12158 14968 12164 14980
rect 12216 14968 12222 15020
rect 12618 15008 12624 15020
rect 12579 14980 12624 15008
rect 12618 14968 12624 14980
rect 12676 14968 12682 15020
rect 12728 15017 12756 15048
rect 12802 15036 12808 15088
rect 12860 15076 12866 15088
rect 12897 15079 12955 15085
rect 12897 15076 12909 15079
rect 12860 15048 12909 15076
rect 12860 15036 12866 15048
rect 12897 15045 12909 15048
rect 12943 15045 12955 15079
rect 13998 15076 14004 15088
rect 12897 15039 12955 15045
rect 13004 15048 14004 15076
rect 13004 15017 13032 15048
rect 13998 15036 14004 15048
rect 14056 15036 14062 15088
rect 17052 15076 17080 15116
rect 17218 15104 17224 15116
rect 17276 15104 17282 15156
rect 17328 15116 19334 15144
rect 17328 15076 17356 15116
rect 18690 15076 18696 15088
rect 17052 15048 17356 15076
rect 18340 15048 18696 15076
rect 18340 15020 18368 15048
rect 18690 15036 18696 15048
rect 18748 15036 18754 15088
rect 12714 15011 12772 15017
rect 12714 14977 12726 15011
rect 12760 14977 12772 15011
rect 12714 14971 12772 14977
rect 12989 15011 13047 15017
rect 12989 14977 13001 15011
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 13127 15011 13185 15017
rect 13127 14977 13139 15011
rect 13173 14977 13185 15011
rect 13127 14971 13185 14977
rect 9766 14940 9772 14952
rect 9416 14912 9772 14940
rect 9766 14900 9772 14912
rect 9824 14900 9830 14952
rect 10321 14943 10379 14949
rect 10321 14909 10333 14943
rect 10367 14940 10379 14943
rect 11330 14940 11336 14952
rect 10367 14912 11336 14940
rect 10367 14909 10379 14912
rect 10321 14903 10379 14909
rect 11330 14900 11336 14912
rect 11388 14900 11394 14952
rect 11698 14900 11704 14952
rect 11756 14940 11762 14952
rect 13142 14940 13170 14971
rect 13906 14968 13912 15020
rect 13964 15008 13970 15020
rect 17129 15011 17187 15017
rect 17129 15008 17141 15011
rect 13964 14980 17141 15008
rect 13964 14968 13970 14980
rect 17129 14977 17141 14980
rect 17175 15008 17187 15011
rect 17175 14980 17264 15008
rect 17175 14977 17187 14980
rect 17129 14971 17187 14977
rect 14642 14940 14648 14952
rect 11756 14912 14648 14940
rect 11756 14900 11762 14912
rect 14642 14900 14648 14912
rect 14700 14900 14706 14952
rect 17236 14940 17264 14980
rect 17310 14968 17316 15020
rect 17368 15008 17374 15020
rect 18322 15008 18328 15020
rect 17368 14980 17413 15008
rect 18235 14980 18328 15008
rect 17368 14968 17374 14980
rect 18322 14968 18328 14980
rect 18380 14968 18386 15020
rect 18414 14968 18420 15020
rect 18472 15008 18478 15020
rect 18581 15011 18639 15017
rect 18581 15008 18593 15011
rect 18472 14980 18593 15008
rect 18472 14968 18478 14980
rect 18581 14977 18593 14980
rect 18627 14977 18639 15011
rect 19306 15008 19334 15116
rect 19426 15104 19432 15156
rect 19484 15144 19490 15156
rect 19705 15147 19763 15153
rect 19705 15144 19717 15147
rect 19484 15116 19717 15144
rect 19484 15104 19490 15116
rect 19705 15113 19717 15116
rect 19751 15113 19763 15147
rect 19705 15107 19763 15113
rect 20717 15147 20775 15153
rect 20717 15113 20729 15147
rect 20763 15144 20775 15147
rect 20898 15144 20904 15156
rect 20763 15116 20904 15144
rect 20763 15113 20775 15116
rect 20717 15107 20775 15113
rect 19720 15076 19748 15107
rect 20898 15104 20904 15116
rect 20956 15104 20962 15156
rect 21174 15144 21180 15156
rect 21135 15116 21180 15144
rect 21174 15104 21180 15116
rect 21232 15104 21238 15156
rect 29638 15144 29644 15156
rect 29599 15116 29644 15144
rect 29638 15104 29644 15116
rect 29696 15104 29702 15156
rect 29914 15104 29920 15156
rect 29972 15144 29978 15156
rect 36173 15147 36231 15153
rect 29972 15116 31892 15144
rect 29972 15104 29978 15116
rect 19720 15048 22692 15076
rect 20533 15011 20591 15017
rect 19306 14980 20484 15008
rect 18581 14971 18639 14977
rect 17865 14943 17923 14949
rect 17865 14940 17877 14943
rect 17236 14912 17877 14940
rect 17865 14909 17877 14912
rect 17911 14909 17923 14943
rect 17865 14903 17923 14909
rect 13265 14875 13323 14881
rect 13265 14872 13277 14875
rect 7392 14844 13277 14872
rect 13265 14841 13277 14844
rect 13311 14841 13323 14875
rect 13265 14835 13323 14841
rect 8754 14804 8760 14816
rect 7300 14776 8760 14804
rect 7193 14767 7251 14773
rect 8754 14764 8760 14776
rect 8812 14764 8818 14816
rect 8846 14764 8852 14816
rect 8904 14804 8910 14816
rect 9582 14804 9588 14816
rect 8904 14776 9588 14804
rect 8904 14764 8910 14776
rect 9582 14764 9588 14776
rect 9640 14764 9646 14816
rect 10042 14804 10048 14816
rect 10003 14776 10048 14804
rect 10042 14764 10048 14776
rect 10100 14764 10106 14816
rect 10413 14807 10471 14813
rect 10413 14773 10425 14807
rect 10459 14804 10471 14807
rect 10502 14804 10508 14816
rect 10459 14776 10508 14804
rect 10459 14773 10471 14776
rect 10413 14767 10471 14773
rect 10502 14764 10508 14776
rect 10560 14764 10566 14816
rect 13906 14804 13912 14816
rect 13867 14776 13912 14804
rect 13906 14764 13912 14776
rect 13964 14764 13970 14816
rect 15194 14764 15200 14816
rect 15252 14804 15258 14816
rect 16022 14804 16028 14816
rect 15252 14776 16028 14804
rect 15252 14764 15258 14776
rect 16022 14764 16028 14776
rect 16080 14764 16086 14816
rect 16298 14764 16304 14816
rect 16356 14804 16362 14816
rect 17310 14804 17316 14816
rect 16356 14776 17316 14804
rect 16356 14764 16362 14776
rect 17310 14764 17316 14776
rect 17368 14764 17374 14816
rect 17880 14804 17908 14903
rect 19886 14900 19892 14952
rect 19944 14940 19950 14952
rect 20349 14943 20407 14949
rect 20349 14940 20361 14943
rect 19944 14912 20361 14940
rect 19944 14900 19950 14912
rect 20349 14909 20361 14912
rect 20395 14909 20407 14943
rect 20349 14903 20407 14909
rect 20456 14872 20484 14980
rect 20533 14977 20545 15011
rect 20579 15008 20591 15011
rect 20622 15008 20628 15020
rect 20579 14980 20628 15008
rect 20579 14977 20591 14980
rect 20533 14971 20591 14977
rect 20622 14968 20628 14980
rect 20680 14968 20686 15020
rect 21174 14968 21180 15020
rect 21232 15008 21238 15020
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21232 14980 22017 15008
rect 21232 14968 21238 14980
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 22094 14968 22100 15020
rect 22152 15008 22158 15020
rect 22664 15017 22692 15048
rect 22738 15036 22744 15088
rect 22796 15076 22802 15088
rect 22833 15079 22891 15085
rect 22833 15076 22845 15079
rect 22796 15048 22845 15076
rect 22796 15036 22802 15048
rect 22833 15045 22845 15048
rect 22879 15045 22891 15079
rect 22833 15039 22891 15045
rect 22925 15079 22983 15085
rect 22925 15045 22937 15079
rect 22971 15076 22983 15079
rect 31754 15076 31760 15088
rect 22971 15048 25084 15076
rect 22971 15045 22983 15048
rect 22925 15039 22983 15045
rect 25056 15020 25084 15048
rect 30208 15048 31760 15076
rect 22189 15011 22247 15017
rect 22189 15008 22201 15011
rect 22152 14980 22201 15008
rect 22152 14968 22158 14980
rect 22189 14977 22201 14980
rect 22235 14977 22247 15011
rect 22189 14971 22247 14977
rect 22649 15011 22707 15017
rect 22649 14977 22661 15011
rect 22695 14977 22707 15011
rect 22649 14971 22707 14977
rect 23017 15011 23075 15017
rect 23017 14977 23029 15011
rect 23063 14977 23075 15011
rect 23017 14971 23075 14977
rect 23032 14940 23060 14971
rect 23474 14968 23480 15020
rect 23532 15008 23538 15020
rect 23661 15011 23719 15017
rect 23661 15008 23673 15011
rect 23532 14980 23673 15008
rect 23532 14968 23538 14980
rect 23661 14977 23673 14980
rect 23707 14977 23719 15011
rect 23842 15008 23848 15020
rect 23803 14980 23848 15008
rect 23661 14971 23719 14977
rect 23566 14940 23572 14952
rect 23032 14912 23572 14940
rect 23566 14900 23572 14912
rect 23624 14900 23630 14952
rect 23676 14940 23704 14971
rect 23842 14968 23848 14980
rect 23900 14968 23906 15020
rect 25038 14968 25044 15020
rect 25096 15008 25102 15020
rect 27157 15011 27215 15017
rect 27157 15008 27169 15011
rect 25096 14980 27169 15008
rect 25096 14968 25102 14980
rect 27157 14977 27169 14980
rect 27203 14977 27215 15011
rect 27157 14971 27215 14977
rect 27341 15011 27399 15017
rect 27341 14977 27353 15011
rect 27387 15008 27399 15011
rect 28626 15008 28632 15020
rect 27387 14980 28632 15008
rect 27387 14977 27399 14980
rect 27341 14971 27399 14977
rect 28626 14968 28632 14980
rect 28684 14968 28690 15020
rect 29086 14968 29092 15020
rect 29144 15008 29150 15020
rect 30122 15017 30180 15023
rect 29871 15011 29929 15017
rect 29871 15008 29883 15011
rect 29144 14980 29883 15008
rect 29144 14968 29150 14980
rect 29871 14977 29883 14980
rect 29917 14977 29929 15011
rect 29871 14971 29929 14977
rect 30009 15011 30067 15017
rect 30009 14977 30021 15011
rect 30055 14977 30067 15011
rect 30122 14983 30134 15017
rect 30168 15014 30180 15017
rect 30208 15014 30236 15048
rect 31754 15036 31760 15048
rect 31812 15036 31818 15088
rect 31864 15076 31892 15116
rect 36173 15113 36185 15147
rect 36219 15144 36231 15147
rect 37734 15144 37740 15156
rect 36219 15116 37740 15144
rect 36219 15113 36231 15116
rect 36173 15107 36231 15113
rect 37734 15104 37740 15116
rect 37792 15104 37798 15156
rect 38562 15144 38568 15156
rect 38120 15116 38568 15144
rect 38120 15076 38148 15116
rect 38562 15104 38568 15116
rect 38620 15104 38626 15156
rect 38654 15104 38660 15156
rect 38712 15144 38718 15156
rect 40221 15147 40279 15153
rect 40221 15144 40233 15147
rect 38712 15116 40233 15144
rect 38712 15104 38718 15116
rect 40221 15113 40233 15116
rect 40267 15113 40279 15147
rect 40221 15107 40279 15113
rect 31864 15048 36308 15076
rect 36280 15020 36308 15048
rect 37752 15048 38148 15076
rect 38381 15079 38439 15085
rect 30168 14986 30236 15014
rect 30297 15011 30355 15017
rect 30168 14983 30180 14986
rect 30122 14977 30180 14983
rect 30297 14977 30309 15011
rect 30343 15006 30355 15011
rect 30466 15008 30472 15020
rect 30392 15006 30472 15008
rect 30343 14980 30472 15006
rect 30343 14978 30420 14980
rect 30343 14977 30355 14978
rect 30009 14971 30067 14977
rect 30297 14971 30355 14977
rect 24305 14943 24363 14949
rect 24305 14940 24317 14943
rect 23676 14912 24317 14940
rect 24305 14909 24317 14912
rect 24351 14909 24363 14943
rect 24305 14903 24363 14909
rect 24394 14900 24400 14952
rect 24452 14940 24458 14952
rect 27062 14940 27068 14952
rect 24452 14912 27068 14940
rect 24452 14900 24458 14912
rect 27062 14900 27068 14912
rect 27120 14900 27126 14952
rect 22186 14872 22192 14884
rect 20456 14844 22094 14872
rect 22147 14844 22192 14872
rect 19426 14804 19432 14816
rect 17880 14776 19432 14804
rect 19426 14764 19432 14776
rect 19484 14804 19490 14816
rect 20254 14804 20260 14816
rect 19484 14776 20260 14804
rect 19484 14764 19490 14776
rect 20254 14764 20260 14776
rect 20312 14764 20318 14816
rect 22066 14804 22094 14844
rect 22186 14832 22192 14844
rect 22244 14832 22250 14884
rect 23106 14804 23112 14816
rect 22066 14776 23112 14804
rect 23106 14764 23112 14776
rect 23164 14764 23170 14816
rect 23201 14807 23259 14813
rect 23201 14773 23213 14807
rect 23247 14804 23259 14807
rect 23566 14804 23572 14816
rect 23247 14776 23572 14804
rect 23247 14773 23259 14776
rect 23201 14767 23259 14773
rect 23566 14764 23572 14776
rect 23624 14764 23630 14816
rect 23842 14804 23848 14816
rect 23803 14776 23848 14804
rect 23842 14764 23848 14776
rect 23900 14764 23906 14816
rect 26973 14807 27031 14813
rect 26973 14773 26985 14807
rect 27019 14804 27031 14807
rect 27338 14804 27344 14816
rect 27019 14776 27344 14804
rect 27019 14773 27031 14776
rect 26973 14767 27031 14773
rect 27338 14764 27344 14776
rect 27396 14764 27402 14816
rect 27706 14764 27712 14816
rect 27764 14804 27770 14816
rect 29086 14804 29092 14816
rect 27764 14776 29092 14804
rect 27764 14764 27770 14776
rect 29086 14764 29092 14776
rect 29144 14764 29150 14816
rect 30021 14804 30049 14971
rect 30466 14968 30472 14980
rect 30524 15008 30530 15020
rect 32398 15008 32404 15020
rect 30524 14980 32404 15008
rect 30524 14968 30530 14980
rect 32398 14968 32404 14980
rect 32456 15008 32462 15020
rect 33321 15011 33379 15017
rect 33321 15008 33333 15011
rect 32456 14980 33333 15008
rect 32456 14968 32462 14980
rect 33321 14977 33333 14980
rect 33367 14977 33379 15011
rect 33594 15008 33600 15020
rect 33555 14980 33600 15008
rect 33321 14971 33379 14977
rect 33594 14968 33600 14980
rect 33652 14968 33658 15020
rect 35069 15011 35127 15017
rect 35069 14977 35081 15011
rect 35115 15008 35127 15011
rect 35434 15008 35440 15020
rect 35115 14980 35440 15008
rect 35115 14977 35127 14980
rect 35069 14971 35127 14977
rect 35434 14968 35440 14980
rect 35492 15008 35498 15020
rect 35989 15011 36047 15017
rect 35989 15008 36001 15011
rect 35492 14980 36001 15008
rect 35492 14968 35498 14980
rect 35989 14977 36001 14980
rect 36035 14977 36047 15011
rect 35989 14971 36047 14977
rect 36262 14968 36268 15020
rect 36320 15008 36326 15020
rect 37752 15017 37780 15048
rect 38381 15045 38393 15079
rect 38427 15076 38439 15079
rect 39086 15079 39144 15085
rect 39086 15076 39098 15079
rect 38427 15048 39098 15076
rect 38427 15045 38439 15048
rect 38381 15039 38439 15045
rect 39086 15045 39098 15048
rect 39132 15045 39144 15079
rect 40957 15079 41015 15085
rect 40957 15076 40969 15079
rect 39086 15039 39144 15045
rect 39224 15048 40969 15076
rect 37918 15017 37924 15020
rect 37737 15011 37795 15017
rect 37737 15008 37749 15011
rect 36320 14980 37749 15008
rect 36320 14968 36326 14980
rect 37737 14977 37749 14980
rect 37783 14977 37795 15011
rect 37916 15008 37924 15017
rect 37879 14980 37924 15008
rect 37737 14971 37795 14977
rect 37916 14971 37924 14980
rect 37918 14968 37924 14971
rect 37976 14968 37982 15020
rect 38016 15011 38074 15017
rect 38016 14977 38028 15011
rect 38062 14977 38074 15011
rect 38016 14971 38074 14977
rect 38151 15011 38209 15017
rect 38151 14977 38163 15011
rect 38197 15008 38209 15011
rect 38286 15008 38292 15020
rect 38197 14980 38292 15008
rect 38197 14977 38209 14980
rect 38151 14971 38209 14977
rect 35342 14940 35348 14952
rect 35303 14912 35348 14940
rect 35342 14900 35348 14912
rect 35400 14900 35406 14952
rect 35802 14940 35808 14952
rect 35715 14912 35808 14940
rect 35802 14900 35808 14912
rect 35860 14940 35866 14952
rect 36633 14943 36691 14949
rect 36633 14940 36645 14943
rect 35860 14912 36645 14940
rect 35860 14900 35866 14912
rect 36633 14909 36645 14912
rect 36679 14909 36691 14943
rect 36633 14903 36691 14909
rect 37550 14900 37556 14952
rect 37608 14940 37614 14952
rect 38028 14940 38056 14971
rect 38286 14968 38292 14980
rect 38344 14968 38350 15020
rect 38562 14968 38568 15020
rect 38620 15008 38626 15020
rect 38746 15008 38752 15020
rect 38620 14980 38752 15008
rect 38620 14968 38626 14980
rect 38746 14968 38752 14980
rect 38804 15008 38810 15020
rect 39224 15008 39252 15048
rect 40957 15045 40969 15048
rect 41003 15076 41015 15079
rect 41322 15076 41328 15088
rect 41003 15048 41328 15076
rect 41003 15045 41015 15048
rect 40957 15039 41015 15045
rect 41322 15036 41328 15048
rect 41380 15036 41386 15088
rect 38804 14980 39252 15008
rect 38804 14968 38810 14980
rect 40310 14968 40316 15020
rect 40368 15008 40374 15020
rect 40678 15008 40684 15020
rect 40368 14980 40684 15008
rect 40368 14968 40374 14980
rect 40678 14968 40684 14980
rect 40736 15008 40742 15020
rect 40773 15011 40831 15017
rect 40773 15008 40785 15011
rect 40736 14980 40785 15008
rect 40736 14968 40742 14980
rect 40773 14977 40785 14980
rect 40819 14977 40831 15011
rect 40773 14971 40831 14977
rect 37608 14912 38056 14940
rect 37608 14900 37614 14912
rect 38654 14900 38660 14952
rect 38712 14940 38718 14952
rect 38841 14943 38899 14949
rect 38841 14940 38853 14943
rect 38712 14912 38853 14940
rect 38712 14900 38718 14912
rect 38841 14909 38853 14912
rect 38887 14909 38899 14943
rect 38841 14903 38899 14909
rect 30098 14804 30104 14816
rect 30021 14776 30104 14804
rect 30098 14764 30104 14776
rect 30156 14764 30162 14816
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 4617 14603 4675 14609
rect 4617 14569 4629 14603
rect 4663 14600 4675 14603
rect 4706 14600 4712 14612
rect 4663 14572 4712 14600
rect 4663 14569 4675 14572
rect 4617 14563 4675 14569
rect 4706 14560 4712 14572
rect 4764 14560 4770 14612
rect 7374 14560 7380 14612
rect 7432 14600 7438 14612
rect 10042 14600 10048 14612
rect 7432 14572 10048 14600
rect 7432 14560 7438 14572
rect 10042 14560 10048 14572
rect 10100 14560 10106 14612
rect 14918 14600 14924 14612
rect 12406 14572 14924 14600
rect 4982 14492 4988 14544
rect 5040 14532 5046 14544
rect 9033 14535 9091 14541
rect 5040 14504 5212 14532
rect 5040 14492 5046 14504
rect 5074 14464 5080 14476
rect 5035 14436 5080 14464
rect 5074 14424 5080 14436
rect 5132 14424 5138 14476
rect 5184 14473 5212 14504
rect 9033 14501 9045 14535
rect 9079 14532 9091 14535
rect 9398 14532 9404 14544
rect 9079 14504 9404 14532
rect 9079 14501 9091 14504
rect 9033 14495 9091 14501
rect 5169 14467 5227 14473
rect 5169 14433 5181 14467
rect 5215 14433 5227 14467
rect 5169 14427 5227 14433
rect 6457 14467 6515 14473
rect 6457 14433 6469 14467
rect 6503 14464 6515 14467
rect 7929 14467 7987 14473
rect 7929 14464 7941 14467
rect 6503 14436 7941 14464
rect 6503 14433 6515 14436
rect 6457 14427 6515 14433
rect 7929 14433 7941 14436
rect 7975 14433 7987 14467
rect 9048 14464 9076 14495
rect 9398 14492 9404 14504
rect 9456 14492 9462 14544
rect 9582 14492 9588 14544
rect 9640 14532 9646 14544
rect 12406 14532 12434 14572
rect 14918 14560 14924 14572
rect 14976 14560 14982 14612
rect 20346 14600 20352 14612
rect 15028 14572 20352 14600
rect 9640 14504 12434 14532
rect 9640 14492 9646 14504
rect 7929 14427 7987 14433
rect 8036 14436 9076 14464
rect 5092 14396 5120 14424
rect 6181 14399 6239 14405
rect 6181 14396 6193 14399
rect 5092 14368 6193 14396
rect 6181 14365 6193 14368
rect 6227 14365 6239 14399
rect 6181 14359 6239 14365
rect 6273 14399 6331 14405
rect 6273 14365 6285 14399
rect 6319 14396 6331 14399
rect 6638 14396 6644 14408
rect 6319 14368 6644 14396
rect 6319 14365 6331 14368
rect 6273 14359 6331 14365
rect 6638 14356 6644 14368
rect 6696 14356 6702 14408
rect 7650 14396 7656 14408
rect 7611 14368 7656 14396
rect 7650 14356 7656 14368
rect 7708 14356 7714 14408
rect 8036 14405 8064 14436
rect 7837 14399 7895 14405
rect 7837 14365 7849 14399
rect 7883 14365 7895 14399
rect 7837 14359 7895 14365
rect 8021 14399 8079 14405
rect 8021 14365 8033 14399
rect 8067 14365 8079 14399
rect 8202 14396 8208 14408
rect 8163 14368 8208 14396
rect 8021 14359 8079 14365
rect 7852 14328 7880 14359
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 11974 14356 11980 14408
rect 12032 14396 12038 14408
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 12032 14368 14105 14396
rect 12032 14356 12038 14368
rect 14093 14365 14105 14368
rect 14139 14365 14151 14399
rect 14093 14359 14151 14365
rect 9582 14328 9588 14340
rect 7852 14300 9588 14328
rect 9582 14288 9588 14300
rect 9640 14288 9646 14340
rect 9766 14288 9772 14340
rect 9824 14328 9830 14340
rect 10134 14328 10140 14340
rect 9824 14300 10140 14328
rect 9824 14288 9830 14300
rect 10134 14288 10140 14300
rect 10192 14328 10198 14340
rect 15028 14328 15056 14572
rect 20346 14560 20352 14572
rect 20404 14560 20410 14612
rect 21082 14560 21088 14612
rect 21140 14600 21146 14612
rect 21821 14603 21879 14609
rect 21821 14600 21833 14603
rect 21140 14572 21833 14600
rect 21140 14560 21146 14572
rect 21821 14569 21833 14572
rect 21867 14600 21879 14603
rect 22278 14600 22284 14612
rect 21867 14572 22284 14600
rect 21867 14569 21879 14572
rect 21821 14563 21879 14569
rect 22278 14560 22284 14572
rect 22336 14560 22342 14612
rect 22664 14572 22876 14600
rect 18230 14532 18236 14544
rect 18143 14504 18236 14532
rect 18230 14492 18236 14504
rect 18288 14532 18294 14544
rect 18288 14504 20852 14532
rect 18288 14492 18294 14504
rect 19889 14467 19947 14473
rect 19889 14433 19901 14467
rect 19935 14464 19947 14467
rect 20441 14467 20499 14473
rect 20441 14464 20453 14467
rect 19935 14436 20453 14464
rect 19935 14433 19947 14436
rect 19889 14427 19947 14433
rect 20441 14433 20453 14436
rect 20487 14464 20499 14467
rect 20530 14464 20536 14476
rect 20487 14436 20536 14464
rect 20487 14433 20499 14436
rect 20441 14427 20499 14433
rect 20530 14424 20536 14436
rect 20588 14424 20594 14476
rect 20622 14424 20628 14476
rect 20680 14464 20686 14476
rect 20717 14467 20775 14473
rect 20717 14464 20729 14467
rect 20680 14436 20729 14464
rect 20680 14424 20686 14436
rect 20717 14433 20729 14436
rect 20763 14433 20775 14467
rect 20717 14427 20775 14433
rect 15102 14356 15108 14408
rect 15160 14396 15166 14408
rect 16853 14399 16911 14405
rect 16853 14396 16865 14399
rect 15160 14368 16865 14396
rect 15160 14356 15166 14368
rect 16853 14365 16865 14368
rect 16899 14396 16911 14399
rect 18322 14396 18328 14408
rect 16899 14368 18328 14396
rect 16899 14365 16911 14368
rect 16853 14359 16911 14365
rect 18322 14356 18328 14368
rect 18380 14356 18386 14408
rect 19426 14356 19432 14408
rect 19484 14396 19490 14408
rect 19797 14399 19855 14405
rect 19797 14396 19809 14399
rect 19484 14368 19809 14396
rect 19484 14356 19490 14368
rect 19797 14365 19809 14368
rect 19843 14365 19855 14399
rect 19797 14359 19855 14365
rect 19981 14399 20039 14405
rect 19981 14365 19993 14399
rect 20027 14396 20039 14399
rect 20070 14396 20076 14408
rect 20027 14368 20076 14396
rect 20027 14365 20039 14368
rect 19981 14359 20039 14365
rect 20070 14356 20076 14368
rect 20128 14356 20134 14408
rect 10192 14300 15056 14328
rect 10192 14288 10198 14300
rect 15930 14288 15936 14340
rect 15988 14328 15994 14340
rect 17126 14337 17132 14340
rect 17120 14328 17132 14337
rect 15988 14300 16988 14328
rect 17087 14300 17132 14328
rect 15988 14288 15994 14300
rect 4985 14263 5043 14269
rect 4985 14229 4997 14263
rect 5031 14260 5043 14263
rect 5534 14260 5540 14272
rect 5031 14232 5540 14260
rect 5031 14229 5043 14232
rect 4985 14223 5043 14229
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 5626 14220 5632 14272
rect 5684 14260 5690 14272
rect 5813 14263 5871 14269
rect 5813 14260 5825 14263
rect 5684 14232 5825 14260
rect 5684 14220 5690 14232
rect 5813 14229 5825 14232
rect 5859 14229 5871 14263
rect 7466 14260 7472 14272
rect 7427 14232 7472 14260
rect 5813 14223 5871 14229
rect 7466 14220 7472 14232
rect 7524 14220 7530 14272
rect 14277 14263 14335 14269
rect 14277 14229 14289 14263
rect 14323 14260 14335 14263
rect 15286 14260 15292 14272
rect 14323 14232 15292 14260
rect 14323 14229 14335 14232
rect 14277 14223 14335 14229
rect 15286 14220 15292 14232
rect 15344 14220 15350 14272
rect 15838 14220 15844 14272
rect 15896 14260 15902 14272
rect 16298 14260 16304 14272
rect 15896 14232 16304 14260
rect 15896 14220 15902 14232
rect 16298 14220 16304 14232
rect 16356 14220 16362 14272
rect 16960 14260 16988 14300
rect 17120 14291 17132 14300
rect 17126 14288 17132 14291
rect 17184 14288 17190 14340
rect 19886 14328 19892 14340
rect 19260 14300 19892 14328
rect 19260 14269 19288 14300
rect 19886 14288 19892 14300
rect 19944 14288 19950 14340
rect 20824 14328 20852 14504
rect 21726 14396 21732 14408
rect 21687 14368 21732 14396
rect 21726 14356 21732 14368
rect 21784 14356 21790 14408
rect 21910 14396 21916 14408
rect 21871 14368 21916 14396
rect 21910 14356 21916 14368
rect 21968 14396 21974 14408
rect 22664 14396 22692 14572
rect 22738 14492 22744 14544
rect 22796 14492 22802 14544
rect 22848 14532 22876 14572
rect 23842 14560 23848 14612
rect 23900 14600 23906 14612
rect 36081 14603 36139 14609
rect 23900 14572 27844 14600
rect 23900 14560 23906 14572
rect 24394 14532 24400 14544
rect 22848 14504 24400 14532
rect 24394 14492 24400 14504
rect 24452 14492 24458 14544
rect 24489 14535 24547 14541
rect 24489 14501 24501 14535
rect 24535 14532 24547 14535
rect 24578 14532 24584 14544
rect 24535 14504 24584 14532
rect 24535 14501 24547 14504
rect 24489 14495 24547 14501
rect 24578 14492 24584 14504
rect 24636 14492 24642 14544
rect 25038 14532 25044 14544
rect 24999 14504 25044 14532
rect 25038 14492 25044 14504
rect 25096 14492 25102 14544
rect 27816 14532 27844 14572
rect 36081 14569 36093 14603
rect 36127 14600 36139 14603
rect 37550 14600 37556 14612
rect 36127 14572 37556 14600
rect 36127 14569 36139 14572
rect 36081 14563 36139 14569
rect 37550 14560 37556 14572
rect 37608 14600 37614 14612
rect 37608 14572 39252 14600
rect 37608 14560 37614 14572
rect 34698 14532 34704 14544
rect 27816 14504 34704 14532
rect 34698 14492 34704 14504
rect 34756 14492 34762 14544
rect 34790 14492 34796 14544
rect 34848 14532 34854 14544
rect 35342 14532 35348 14544
rect 34848 14504 35348 14532
rect 34848 14492 34854 14504
rect 35342 14492 35348 14504
rect 35400 14532 35406 14544
rect 35400 14504 36216 14532
rect 35400 14492 35406 14504
rect 22756 14464 22784 14492
rect 22756 14436 22968 14464
rect 22940 14405 22968 14436
rect 28258 14424 28264 14476
rect 28316 14464 28322 14476
rect 33321 14467 33379 14473
rect 33321 14464 33333 14467
rect 28316 14436 33333 14464
rect 28316 14424 28322 14436
rect 33321 14433 33333 14436
rect 33367 14464 33379 14467
rect 33781 14467 33839 14473
rect 33781 14464 33793 14467
rect 33367 14436 33793 14464
rect 33367 14433 33379 14436
rect 33321 14427 33379 14433
rect 33781 14433 33793 14436
rect 33827 14464 33839 14467
rect 35802 14464 35808 14476
rect 33827 14436 35808 14464
rect 33827 14433 33839 14436
rect 33781 14427 33839 14433
rect 35802 14424 35808 14436
rect 35860 14424 35866 14476
rect 21968 14368 22692 14396
rect 22741 14399 22799 14405
rect 21968 14356 21974 14368
rect 22741 14365 22753 14399
rect 22787 14365 22799 14399
rect 22741 14359 22799 14365
rect 22925 14399 22983 14405
rect 22925 14365 22937 14399
rect 22971 14365 22983 14399
rect 22925 14359 22983 14365
rect 23109 14399 23167 14405
rect 23109 14365 23121 14399
rect 23155 14396 23167 14399
rect 23474 14396 23480 14408
rect 23155 14368 23480 14396
rect 23155 14365 23167 14368
rect 23109 14359 23167 14365
rect 22756 14328 22784 14359
rect 23474 14356 23480 14368
rect 23532 14356 23538 14408
rect 25406 14356 25412 14408
rect 25464 14396 25470 14408
rect 26421 14399 26479 14405
rect 26421 14396 26433 14399
rect 25464 14368 26433 14396
rect 25464 14356 25470 14368
rect 26421 14365 26433 14368
rect 26467 14396 26479 14399
rect 26881 14399 26939 14405
rect 26881 14396 26893 14399
rect 26467 14368 26893 14396
rect 26467 14365 26479 14368
rect 26421 14359 26479 14365
rect 26881 14365 26893 14368
rect 26927 14365 26939 14399
rect 26881 14359 26939 14365
rect 28626 14356 28632 14408
rect 28684 14396 28690 14408
rect 29549 14399 29607 14405
rect 29549 14396 29561 14399
rect 28684 14368 29561 14396
rect 28684 14356 28690 14368
rect 29549 14365 29561 14368
rect 29595 14396 29607 14399
rect 31386 14396 31392 14408
rect 29595 14368 31392 14396
rect 29595 14365 29607 14368
rect 29549 14359 29607 14365
rect 31386 14356 31392 14368
rect 31444 14356 31450 14408
rect 33965 14399 34023 14405
rect 33965 14365 33977 14399
rect 34011 14365 34023 14399
rect 34698 14396 34704 14408
rect 34659 14368 34704 14396
rect 33965 14359 34023 14365
rect 20824 14300 22784 14328
rect 23017 14331 23075 14337
rect 23017 14297 23029 14331
rect 23063 14328 23075 14331
rect 26176 14331 26234 14337
rect 23063 14300 26096 14328
rect 23063 14297 23075 14300
rect 23017 14291 23075 14297
rect 19245 14263 19303 14269
rect 19245 14260 19257 14263
rect 16960 14232 19257 14260
rect 19245 14229 19257 14232
rect 19291 14229 19303 14263
rect 19245 14223 19303 14229
rect 19334 14220 19340 14272
rect 19392 14260 19398 14272
rect 20070 14260 20076 14272
rect 19392 14232 20076 14260
rect 19392 14220 19398 14232
rect 20070 14220 20076 14232
rect 20128 14260 20134 14272
rect 20622 14260 20628 14272
rect 20128 14232 20628 14260
rect 20128 14220 20134 14232
rect 20622 14220 20628 14232
rect 20680 14220 20686 14272
rect 23293 14263 23351 14269
rect 23293 14229 23305 14263
rect 23339 14260 23351 14263
rect 23658 14260 23664 14272
rect 23339 14232 23664 14260
rect 23339 14229 23351 14232
rect 23293 14223 23351 14229
rect 23658 14220 23664 14232
rect 23716 14220 23722 14272
rect 23842 14260 23848 14272
rect 23803 14232 23848 14260
rect 23842 14220 23848 14232
rect 23900 14220 23906 14272
rect 26068 14260 26096 14300
rect 26176 14297 26188 14331
rect 26222 14328 26234 14331
rect 26970 14328 26976 14340
rect 26222 14300 26976 14328
rect 26222 14297 26234 14300
rect 26176 14291 26234 14297
rect 26970 14288 26976 14300
rect 27028 14288 27034 14340
rect 27154 14337 27160 14340
rect 27148 14291 27160 14337
rect 27212 14328 27218 14340
rect 27212 14300 27248 14328
rect 27154 14288 27160 14291
rect 27212 14288 27218 14300
rect 29638 14288 29644 14340
rect 29696 14328 29702 14340
rect 29733 14331 29791 14337
rect 29733 14328 29745 14331
rect 29696 14300 29745 14328
rect 29696 14288 29702 14300
rect 29733 14297 29745 14300
rect 29779 14297 29791 14331
rect 33980 14328 34008 14359
rect 34698 14356 34704 14368
rect 34756 14356 34762 14408
rect 34977 14399 35035 14405
rect 34977 14365 34989 14399
rect 35023 14396 35035 14399
rect 35526 14396 35532 14408
rect 35023 14368 35532 14396
rect 35023 14365 35035 14368
rect 34977 14359 35035 14365
rect 34992 14328 35020 14359
rect 35526 14356 35532 14368
rect 35584 14356 35590 14408
rect 36188 14405 36216 14504
rect 37274 14492 37280 14544
rect 37332 14492 37338 14544
rect 37292 14464 37320 14492
rect 37292 14436 38424 14464
rect 38396 14408 38424 14436
rect 35989 14399 36047 14405
rect 35989 14365 36001 14399
rect 36035 14365 36047 14399
rect 35989 14359 36047 14365
rect 36173 14399 36231 14405
rect 36173 14365 36185 14399
rect 36219 14365 36231 14399
rect 36173 14359 36231 14365
rect 37277 14399 37335 14405
rect 37277 14365 37289 14399
rect 37323 14396 37335 14399
rect 37458 14396 37464 14408
rect 37323 14368 37464 14396
rect 37323 14365 37335 14368
rect 37277 14359 37335 14365
rect 33980 14300 35020 14328
rect 29733 14291 29791 14297
rect 35434 14288 35440 14340
rect 35492 14328 35498 14340
rect 36004 14328 36032 14359
rect 37458 14356 37464 14368
rect 37516 14356 37522 14408
rect 37553 14399 37611 14405
rect 37553 14365 37565 14399
rect 37599 14396 37611 14399
rect 37734 14396 37740 14408
rect 37599 14368 37740 14396
rect 37599 14365 37611 14368
rect 37553 14359 37611 14365
rect 37734 14356 37740 14368
rect 37792 14356 37798 14408
rect 38378 14396 38384 14408
rect 38291 14368 38384 14396
rect 38378 14356 38384 14368
rect 38436 14356 38442 14408
rect 39224 14405 39252 14572
rect 39209 14399 39267 14405
rect 39209 14365 39221 14399
rect 39255 14365 39267 14399
rect 58158 14396 58164 14408
rect 58119 14368 58164 14396
rect 39209 14359 39267 14365
rect 58158 14356 58164 14368
rect 58216 14356 58222 14408
rect 35492 14300 36032 14328
rect 37476 14328 37504 14356
rect 38197 14331 38255 14337
rect 38197 14328 38209 14331
rect 37476 14300 38209 14328
rect 35492 14288 35498 14300
rect 38197 14297 38209 14300
rect 38243 14297 38255 14331
rect 39022 14328 39028 14340
rect 38983 14300 39028 14328
rect 38197 14291 38255 14297
rect 39022 14288 39028 14300
rect 39080 14288 39086 14340
rect 40310 14328 40316 14340
rect 40271 14300 40316 14328
rect 40310 14288 40316 14300
rect 40368 14288 40374 14340
rect 28261 14263 28319 14269
rect 28261 14260 28273 14263
rect 26068 14232 28273 14260
rect 28261 14229 28273 14232
rect 28307 14260 28319 14263
rect 28442 14260 28448 14272
rect 28307 14232 28448 14260
rect 28307 14229 28319 14232
rect 28261 14223 28319 14229
rect 28442 14220 28448 14232
rect 28500 14220 28506 14272
rect 29822 14220 29828 14272
rect 29880 14260 29886 14272
rect 29917 14263 29975 14269
rect 29917 14260 29929 14263
rect 29880 14232 29929 14260
rect 29880 14220 29886 14232
rect 29917 14229 29929 14232
rect 29963 14229 29975 14263
rect 29917 14223 29975 14229
rect 34149 14263 34207 14269
rect 34149 14229 34161 14263
rect 34195 14260 34207 14263
rect 36722 14260 36728 14272
rect 34195 14232 36728 14260
rect 34195 14229 34207 14232
rect 34149 14223 34207 14229
rect 36722 14220 36728 14232
rect 36780 14220 36786 14272
rect 38562 14260 38568 14272
rect 38523 14232 38568 14260
rect 38562 14220 38568 14232
rect 38620 14220 38626 14272
rect 40402 14260 40408 14272
rect 40363 14232 40408 14260
rect 40402 14220 40408 14232
rect 40460 14220 40466 14272
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 7650 14016 7656 14068
rect 7708 14056 7714 14068
rect 8481 14059 8539 14065
rect 8481 14056 8493 14059
rect 7708 14028 8493 14056
rect 7708 14016 7714 14028
rect 8481 14025 8493 14028
rect 8527 14056 8539 14059
rect 9766 14056 9772 14068
rect 8527 14028 9772 14056
rect 8527 14025 8539 14028
rect 8481 14019 8539 14025
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 13173 14059 13231 14065
rect 13173 14025 13185 14059
rect 13219 14056 13231 14059
rect 13998 14056 14004 14068
rect 13219 14028 14004 14056
rect 13219 14025 13231 14028
rect 13173 14019 13231 14025
rect 13998 14016 14004 14028
rect 14056 14016 14062 14068
rect 16850 14016 16856 14068
rect 16908 14056 16914 14068
rect 21269 14059 21327 14065
rect 16908 14028 20668 14056
rect 16908 14016 16914 14028
rect 7368 13991 7426 13997
rect 7368 13957 7380 13991
rect 7414 13988 7426 13991
rect 7466 13988 7472 14000
rect 7414 13960 7472 13988
rect 7414 13957 7426 13960
rect 7368 13951 7426 13957
rect 7466 13948 7472 13960
rect 7524 13948 7530 14000
rect 7558 13948 7564 14000
rect 7616 13988 7622 14000
rect 7616 13960 12204 13988
rect 7616 13948 7622 13960
rect 12176 13932 12204 13960
rect 14918 13948 14924 14000
rect 14976 13988 14982 14000
rect 18325 13991 18383 13997
rect 18325 13988 18337 13991
rect 14976 13960 18337 13988
rect 14976 13948 14982 13960
rect 18325 13957 18337 13960
rect 18371 13988 18383 13991
rect 18877 13991 18935 13997
rect 18877 13988 18889 13991
rect 18371 13960 18889 13988
rect 18371 13957 18383 13960
rect 18325 13951 18383 13957
rect 18877 13957 18889 13960
rect 18923 13988 18935 13991
rect 19334 13988 19340 14000
rect 18923 13960 19340 13988
rect 18923 13957 18935 13960
rect 18877 13951 18935 13957
rect 19334 13948 19340 13960
rect 19392 13948 19398 14000
rect 19426 13948 19432 14000
rect 19484 13988 19490 14000
rect 19613 13991 19671 13997
rect 19613 13988 19625 13991
rect 19484 13960 19625 13988
rect 19484 13948 19490 13960
rect 19613 13957 19625 13960
rect 19659 13957 19671 13991
rect 20530 13988 20536 14000
rect 20491 13960 20536 13988
rect 19613 13951 19671 13957
rect 20530 13948 20536 13960
rect 20588 13948 20594 14000
rect 20640 13988 20668 14028
rect 21269 14025 21281 14059
rect 21315 14056 21327 14059
rect 21910 14056 21916 14068
rect 21315 14028 21916 14056
rect 21315 14025 21327 14028
rect 21269 14019 21327 14025
rect 21910 14016 21916 14028
rect 21968 14016 21974 14068
rect 22738 14056 22744 14068
rect 22572 14028 22744 14056
rect 22572 13997 22600 14028
rect 22738 14016 22744 14028
rect 22796 14016 22802 14068
rect 23106 14016 23112 14068
rect 23164 14056 23170 14068
rect 23385 14059 23443 14065
rect 23385 14056 23397 14059
rect 23164 14028 23397 14056
rect 23164 14016 23170 14028
rect 23385 14025 23397 14028
rect 23431 14025 23443 14059
rect 23385 14019 23443 14025
rect 25406 14016 25412 14068
rect 25464 14056 25470 14068
rect 25593 14059 25651 14065
rect 25593 14056 25605 14059
rect 25464 14028 25605 14056
rect 25464 14016 25470 14028
rect 25593 14025 25605 14028
rect 25639 14025 25651 14059
rect 27154 14056 27160 14068
rect 27115 14028 27160 14056
rect 25593 14019 25651 14025
rect 27154 14016 27160 14028
rect 27212 14016 27218 14068
rect 29638 14056 29644 14068
rect 27264 14028 29644 14056
rect 22557 13991 22615 13997
rect 20640 13960 22416 13988
rect 10042 13880 10048 13932
rect 10100 13920 10106 13932
rect 10606 13923 10664 13929
rect 10606 13920 10618 13923
rect 10100 13892 10618 13920
rect 10100 13880 10106 13892
rect 10606 13889 10618 13892
rect 10652 13889 10664 13923
rect 10870 13920 10876 13932
rect 10831 13892 10876 13920
rect 10606 13883 10664 13889
rect 10870 13880 10876 13892
rect 10928 13880 10934 13932
rect 11974 13920 11980 13932
rect 11935 13892 11980 13920
rect 11974 13880 11980 13892
rect 12032 13880 12038 13932
rect 12158 13920 12164 13932
rect 12119 13892 12164 13920
rect 12158 13880 12164 13892
rect 12216 13880 12222 13932
rect 14274 13920 14280 13932
rect 14332 13929 14338 13932
rect 14244 13892 14280 13920
rect 14274 13880 14280 13892
rect 14332 13883 14344 13929
rect 14553 13923 14611 13929
rect 14553 13889 14565 13923
rect 14599 13920 14611 13923
rect 15102 13920 15108 13932
rect 14599 13892 15108 13920
rect 14599 13889 14611 13892
rect 14553 13883 14611 13889
rect 14332 13880 14338 13883
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 16298 13880 16304 13932
rect 16356 13920 16362 13932
rect 21821 13923 21879 13929
rect 21821 13920 21833 13923
rect 16356 13892 21833 13920
rect 16356 13880 16362 13892
rect 21821 13889 21833 13892
rect 21867 13920 21879 13923
rect 22094 13920 22100 13932
rect 21867 13892 22100 13920
rect 21867 13889 21879 13892
rect 21821 13883 21879 13889
rect 22094 13880 22100 13892
rect 22152 13880 22158 13932
rect 22388 13929 22416 13960
rect 22557 13957 22569 13991
rect 22603 13957 22615 13991
rect 22557 13951 22615 13957
rect 22649 13991 22707 13997
rect 22649 13957 22661 13991
rect 22695 13988 22707 13991
rect 27264 13988 27292 14028
rect 29638 14016 29644 14028
rect 29696 14016 29702 14068
rect 30006 14016 30012 14068
rect 30064 14056 30070 14068
rect 34517 14059 34575 14065
rect 34517 14056 34529 14059
rect 30064 14028 34529 14056
rect 30064 14016 30070 14028
rect 34517 14025 34529 14028
rect 34563 14056 34575 14059
rect 34790 14056 34796 14068
rect 34563 14028 34796 14056
rect 34563 14025 34575 14028
rect 34517 14019 34575 14025
rect 34790 14016 34796 14028
rect 34848 14016 34854 14068
rect 28261 13991 28319 13997
rect 28261 13988 28273 13991
rect 22695 13960 27292 13988
rect 27724 13960 28273 13988
rect 22695 13957 22707 13960
rect 22649 13951 22707 13957
rect 22373 13923 22431 13929
rect 22373 13889 22385 13923
rect 22419 13889 22431 13923
rect 22373 13883 22431 13889
rect 22741 13923 22799 13929
rect 22741 13889 22753 13923
rect 22787 13920 22799 13923
rect 23474 13920 23480 13932
rect 22787 13892 23480 13920
rect 22787 13889 22799 13892
rect 22741 13883 22799 13889
rect 23474 13880 23480 13892
rect 23532 13880 23538 13932
rect 23569 13923 23627 13929
rect 23569 13889 23581 13923
rect 23615 13889 23627 13923
rect 23569 13883 23627 13889
rect 23845 13923 23903 13929
rect 23845 13889 23857 13923
rect 23891 13889 23903 13923
rect 23845 13883 23903 13889
rect 24305 13923 24363 13929
rect 24305 13889 24317 13923
rect 24351 13920 24363 13923
rect 25958 13920 25964 13932
rect 24351 13892 25964 13920
rect 24351 13889 24363 13892
rect 24305 13883 24363 13889
rect 5534 13852 5540 13864
rect 5495 13824 5540 13852
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 7098 13852 7104 13864
rect 7059 13824 7104 13852
rect 7098 13812 7104 13824
rect 7156 13812 7162 13864
rect 14642 13812 14648 13864
rect 14700 13852 14706 13864
rect 20717 13855 20775 13861
rect 20717 13852 20729 13855
rect 14700 13824 20729 13852
rect 14700 13812 14706 13824
rect 20717 13821 20729 13824
rect 20763 13852 20775 13855
rect 21726 13852 21732 13864
rect 20763 13824 21732 13852
rect 20763 13821 20775 13824
rect 20717 13815 20775 13821
rect 21726 13812 21732 13824
rect 21784 13812 21790 13864
rect 8754 13744 8760 13796
rect 8812 13784 8818 13796
rect 9858 13784 9864 13796
rect 8812 13756 9864 13784
rect 8812 13744 8818 13756
rect 9858 13744 9864 13756
rect 9916 13744 9922 13796
rect 17586 13744 17592 13796
rect 17644 13784 17650 13796
rect 17770 13784 17776 13796
rect 17644 13756 17776 13784
rect 17644 13744 17650 13756
rect 17770 13744 17776 13756
rect 17828 13744 17834 13796
rect 23584 13784 23612 13883
rect 23750 13852 23756 13864
rect 23711 13824 23756 13852
rect 23750 13812 23756 13824
rect 23808 13812 23814 13864
rect 23860 13852 23888 13883
rect 25958 13880 25964 13892
rect 26016 13880 26022 13932
rect 27062 13880 27068 13932
rect 27120 13920 27126 13932
rect 27522 13929 27528 13932
rect 27413 13923 27471 13929
rect 27413 13920 27425 13923
rect 27120 13892 27425 13920
rect 27120 13880 27126 13892
rect 27413 13889 27425 13892
rect 27459 13889 27471 13923
rect 27413 13883 27471 13889
rect 27506 13923 27528 13929
rect 27506 13889 27518 13923
rect 27506 13883 27528 13889
rect 27522 13880 27528 13883
rect 27580 13880 27586 13932
rect 27617 13923 27675 13929
rect 27617 13889 27629 13923
rect 27663 13920 27675 13923
rect 27724 13920 27752 13960
rect 28261 13957 28273 13960
rect 28307 13957 28319 13991
rect 28442 13988 28448 14000
rect 28403 13960 28448 13988
rect 28261 13951 28319 13957
rect 28442 13948 28448 13960
rect 28500 13948 28506 14000
rect 28626 13988 28632 14000
rect 28587 13960 28632 13988
rect 28626 13948 28632 13960
rect 28684 13948 28690 14000
rect 30190 13988 30196 14000
rect 29656 13960 30196 13988
rect 27663 13892 27752 13920
rect 27801 13926 27859 13929
rect 27801 13923 27936 13926
rect 27663 13889 27675 13892
rect 27617 13883 27675 13889
rect 27801 13889 27813 13923
rect 27847 13920 27936 13923
rect 28074 13920 28080 13932
rect 27847 13898 28080 13920
rect 27847 13889 27859 13898
rect 27908 13892 28080 13898
rect 27801 13883 27859 13889
rect 28074 13880 28080 13892
rect 28132 13880 28138 13932
rect 29086 13920 29092 13932
rect 29047 13892 29092 13920
rect 29086 13880 29092 13892
rect 29144 13880 29150 13932
rect 29656 13929 29684 13960
rect 30190 13948 30196 13960
rect 30248 13948 30254 14000
rect 36446 13948 36452 14000
rect 36504 13988 36510 14000
rect 36541 13991 36599 13997
rect 36541 13988 36553 13991
rect 36504 13960 36553 13988
rect 36504 13948 36510 13960
rect 36541 13957 36553 13960
rect 36587 13957 36599 13991
rect 37642 13988 37648 14000
rect 37603 13960 37648 13988
rect 36541 13951 36599 13957
rect 37642 13948 37648 13960
rect 37700 13948 37706 14000
rect 29641 13923 29699 13929
rect 29641 13889 29653 13923
rect 29687 13889 29699 13923
rect 29822 13920 29828 13932
rect 29783 13892 29828 13920
rect 29641 13883 29699 13889
rect 29822 13880 29828 13892
rect 29880 13880 29886 13932
rect 29917 13923 29975 13929
rect 29917 13889 29929 13923
rect 29963 13889 29975 13923
rect 29917 13883 29975 13889
rect 30009 13923 30067 13929
rect 30009 13889 30021 13923
rect 30055 13920 30067 13923
rect 35621 13923 35679 13929
rect 30055 13892 30236 13920
rect 30055 13889 30067 13892
rect 30009 13883 30067 13889
rect 24578 13852 24584 13864
rect 23860 13824 24584 13852
rect 24578 13812 24584 13824
rect 24636 13812 24642 13864
rect 27540 13852 27568 13880
rect 29932 13852 29960 13883
rect 30098 13852 30104 13864
rect 27540 13824 30104 13852
rect 30098 13812 30104 13824
rect 30156 13812 30162 13864
rect 23842 13784 23848 13796
rect 23584 13756 23848 13784
rect 23842 13744 23848 13756
rect 23900 13784 23906 13796
rect 24302 13784 24308 13796
rect 23900 13756 24308 13784
rect 23900 13744 23906 13756
rect 24302 13744 24308 13756
rect 24360 13744 24366 13796
rect 29086 13744 29092 13796
rect 29144 13784 29150 13796
rect 30208 13784 30236 13892
rect 35621 13889 35633 13923
rect 35667 13920 35679 13923
rect 36262 13920 36268 13932
rect 35667 13892 36268 13920
rect 35667 13889 35679 13892
rect 35621 13883 35679 13889
rect 36262 13880 36268 13892
rect 36320 13880 36326 13932
rect 36722 13920 36728 13932
rect 36635 13892 36728 13920
rect 36722 13880 36728 13892
rect 36780 13920 36786 13932
rect 37458 13920 37464 13932
rect 36780 13892 37464 13920
rect 36780 13880 36786 13892
rect 37458 13880 37464 13892
rect 37516 13920 37522 13932
rect 38194 13920 38200 13932
rect 37516 13892 38200 13920
rect 37516 13880 37522 13892
rect 38194 13880 38200 13892
rect 38252 13880 38258 13932
rect 30285 13855 30343 13861
rect 30285 13821 30297 13855
rect 30331 13852 30343 13855
rect 30742 13852 30748 13864
rect 30331 13824 30748 13852
rect 30331 13821 30343 13824
rect 30285 13815 30343 13821
rect 30742 13812 30748 13824
rect 30800 13812 30806 13864
rect 33594 13812 33600 13864
rect 33652 13852 33658 13864
rect 35897 13855 35955 13861
rect 35897 13852 35909 13855
rect 33652 13824 35909 13852
rect 33652 13812 33658 13824
rect 35897 13821 35909 13824
rect 35943 13852 35955 13855
rect 40310 13852 40316 13864
rect 35943 13824 40316 13852
rect 35943 13821 35955 13824
rect 35897 13815 35955 13821
rect 40310 13812 40316 13824
rect 40368 13812 40374 13864
rect 29144 13756 30236 13784
rect 29144 13744 29150 13756
rect 9490 13716 9496 13728
rect 9451 13688 9496 13716
rect 9490 13676 9496 13688
rect 9548 13676 9554 13728
rect 22925 13719 22983 13725
rect 22925 13685 22937 13719
rect 22971 13716 22983 13719
rect 23198 13716 23204 13728
rect 22971 13688 23204 13716
rect 22971 13685 22983 13688
rect 22925 13679 22983 13685
rect 23198 13676 23204 13688
rect 23256 13676 23262 13728
rect 23566 13716 23572 13728
rect 23527 13688 23572 13716
rect 23566 13676 23572 13688
rect 23624 13676 23630 13728
rect 23934 13676 23940 13728
rect 23992 13716 23998 13728
rect 27798 13716 27804 13728
rect 23992 13688 27804 13716
rect 23992 13676 23998 13688
rect 27798 13676 27804 13688
rect 27856 13676 27862 13728
rect 29270 13676 29276 13728
rect 29328 13716 29334 13728
rect 30834 13716 30840 13728
rect 29328 13688 30840 13716
rect 29328 13676 29334 13688
rect 30834 13676 30840 13688
rect 30892 13676 30898 13728
rect 36078 13676 36084 13728
rect 36136 13716 36142 13728
rect 36357 13719 36415 13725
rect 36357 13716 36369 13719
rect 36136 13688 36369 13716
rect 36136 13676 36142 13688
rect 36357 13685 36369 13688
rect 36403 13685 36415 13719
rect 36357 13679 36415 13685
rect 38654 13676 38660 13728
rect 38712 13716 38718 13728
rect 38933 13719 38991 13725
rect 38933 13716 38945 13719
rect 38712 13688 38945 13716
rect 38712 13676 38718 13688
rect 38933 13685 38945 13688
rect 38979 13685 38991 13719
rect 38933 13679 38991 13685
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 2317 13515 2375 13521
rect 2317 13481 2329 13515
rect 2363 13512 2375 13515
rect 2406 13512 2412 13524
rect 2363 13484 2412 13512
rect 2363 13481 2375 13484
rect 2317 13475 2375 13481
rect 2406 13472 2412 13484
rect 2464 13472 2470 13524
rect 4525 13515 4583 13521
rect 4525 13481 4537 13515
rect 4571 13512 4583 13515
rect 4614 13512 4620 13524
rect 4571 13484 4620 13512
rect 4571 13481 4583 13484
rect 4525 13475 4583 13481
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 9582 13472 9588 13524
rect 9640 13512 9646 13524
rect 9953 13515 10011 13521
rect 9640 13484 9720 13512
rect 9640 13472 9646 13484
rect 9398 13404 9404 13456
rect 9456 13404 9462 13456
rect 6638 13336 6644 13388
rect 6696 13376 6702 13388
rect 6825 13379 6883 13385
rect 6825 13376 6837 13379
rect 6696 13348 6837 13376
rect 6696 13336 6702 13348
rect 6825 13345 6837 13348
rect 6871 13345 6883 13379
rect 9416 13376 9444 13404
rect 9493 13379 9551 13385
rect 9493 13376 9505 13379
rect 9416 13348 9505 13376
rect 6825 13339 6883 13345
rect 9493 13345 9505 13348
rect 9539 13345 9551 13379
rect 9493 13339 9551 13345
rect 9585 13379 9643 13385
rect 9585 13345 9597 13379
rect 9631 13376 9643 13379
rect 9692 13376 9720 13484
rect 9953 13481 9965 13515
rect 9999 13512 10011 13515
rect 10042 13512 10048 13524
rect 9999 13484 10048 13512
rect 9999 13481 10011 13484
rect 9953 13475 10011 13481
rect 10042 13472 10048 13484
rect 10100 13472 10106 13524
rect 10505 13515 10563 13521
rect 10505 13481 10517 13515
rect 10551 13512 10563 13515
rect 10594 13512 10600 13524
rect 10551 13484 10600 13512
rect 10551 13481 10563 13484
rect 10505 13475 10563 13481
rect 10594 13472 10600 13484
rect 10652 13472 10658 13524
rect 17770 13472 17776 13524
rect 17828 13512 17834 13524
rect 18601 13515 18659 13521
rect 18601 13512 18613 13515
rect 17828 13484 18613 13512
rect 17828 13472 17834 13484
rect 18601 13481 18613 13484
rect 18647 13481 18659 13515
rect 20530 13512 20536 13524
rect 20491 13484 20536 13512
rect 18601 13475 18659 13481
rect 20530 13472 20536 13484
rect 20588 13472 20594 13524
rect 23198 13512 23204 13524
rect 23159 13484 23204 13512
rect 23198 13472 23204 13484
rect 23256 13472 23262 13524
rect 23658 13472 23664 13524
rect 23716 13512 23722 13524
rect 24857 13515 24915 13521
rect 24857 13512 24869 13515
rect 23716 13484 24869 13512
rect 23716 13472 23722 13484
rect 24857 13481 24869 13484
rect 24903 13481 24915 13515
rect 25958 13512 25964 13524
rect 25871 13484 25964 13512
rect 24857 13475 24915 13481
rect 25958 13472 25964 13484
rect 26016 13512 26022 13524
rect 32490 13512 32496 13524
rect 26016 13484 32496 13512
rect 26016 13472 26022 13484
rect 32490 13472 32496 13484
rect 32548 13512 32554 13524
rect 37642 13512 37648 13524
rect 32548 13484 37648 13512
rect 32548 13472 32554 13484
rect 37642 13472 37648 13484
rect 37700 13472 37706 13524
rect 9858 13404 9864 13456
rect 9916 13444 9922 13456
rect 23017 13447 23075 13453
rect 23017 13444 23029 13447
rect 9916 13416 23029 13444
rect 9916 13404 9922 13416
rect 23017 13413 23029 13416
rect 23063 13413 23075 13447
rect 23017 13407 23075 13413
rect 24489 13447 24547 13453
rect 24489 13413 24501 13447
rect 24535 13413 24547 13447
rect 26970 13444 26976 13456
rect 26931 13416 26976 13444
rect 24489 13407 24547 13413
rect 9631 13348 9720 13376
rect 9631 13345 9643 13348
rect 9585 13339 9643 13345
rect 11330 13336 11336 13388
rect 11388 13376 11394 13388
rect 24504 13376 24532 13407
rect 26970 13404 26976 13416
rect 27028 13404 27034 13456
rect 27522 13444 27528 13456
rect 27353 13416 27528 13444
rect 11388 13348 24532 13376
rect 11388 13336 11394 13348
rect 2501 13311 2559 13317
rect 2501 13277 2513 13311
rect 2547 13308 2559 13311
rect 3878 13308 3884 13320
rect 2547 13280 3884 13308
rect 2547 13277 2559 13280
rect 2501 13271 2559 13277
rect 3878 13268 3884 13280
rect 3936 13268 3942 13320
rect 5074 13268 5080 13320
rect 5132 13308 5138 13320
rect 6733 13311 6791 13317
rect 6733 13308 6745 13311
rect 5132 13280 6745 13308
rect 5132 13268 5138 13280
rect 6733 13277 6745 13280
rect 6779 13277 6791 13311
rect 6733 13271 6791 13277
rect 8202 13268 8208 13320
rect 8260 13308 8266 13320
rect 9217 13311 9275 13317
rect 9217 13308 9229 13311
rect 8260 13280 9229 13308
rect 8260 13268 8266 13280
rect 9217 13277 9229 13280
rect 9263 13277 9275 13311
rect 9217 13271 9275 13277
rect 9401 13311 9459 13317
rect 9401 13277 9413 13311
rect 9447 13308 9459 13311
rect 9769 13311 9827 13317
rect 9447 13306 9545 13308
rect 9447 13280 9674 13306
rect 9447 13277 9459 13280
rect 9517 13278 9674 13280
rect 9401 13271 9459 13277
rect 9646 13240 9674 13278
rect 9769 13277 9781 13311
rect 9815 13308 9827 13311
rect 9858 13308 9864 13320
rect 9815 13280 9864 13308
rect 9815 13277 9827 13280
rect 9769 13271 9827 13277
rect 9858 13268 9864 13280
rect 9916 13268 9922 13320
rect 13998 13268 14004 13320
rect 14056 13308 14062 13320
rect 14277 13311 14335 13317
rect 14277 13308 14289 13311
rect 14056 13280 14289 13308
rect 14056 13268 14062 13280
rect 14277 13277 14289 13280
rect 14323 13277 14335 13311
rect 19426 13308 19432 13320
rect 14277 13271 14335 13277
rect 17696 13280 19432 13308
rect 10594 13240 10600 13252
rect 9646 13212 10600 13240
rect 10594 13200 10600 13212
rect 10652 13200 10658 13252
rect 14090 13240 14096 13252
rect 14051 13212 14096 13240
rect 14090 13200 14096 13212
rect 14148 13240 14154 13252
rect 17696 13249 17724 13280
rect 19426 13268 19432 13280
rect 19484 13268 19490 13320
rect 23198 13308 23204 13320
rect 23159 13280 23204 13308
rect 23198 13268 23204 13280
rect 23256 13268 23262 13320
rect 23293 13311 23351 13317
rect 23293 13277 23305 13311
rect 23339 13308 23351 13311
rect 24210 13308 24216 13320
rect 23339 13280 24216 13308
rect 23339 13277 23351 13280
rect 23293 13271 23351 13277
rect 24210 13268 24216 13280
rect 24268 13268 24274 13320
rect 24578 13268 24584 13320
rect 24636 13308 24642 13320
rect 24673 13311 24731 13317
rect 24673 13308 24685 13311
rect 24636 13280 24685 13308
rect 24636 13268 24642 13280
rect 24673 13277 24685 13280
rect 24719 13277 24731 13311
rect 24673 13271 24731 13277
rect 24765 13311 24823 13317
rect 24765 13277 24777 13311
rect 24811 13277 24823 13311
rect 24765 13271 24823 13277
rect 24949 13311 25007 13317
rect 24949 13277 24961 13311
rect 24995 13308 25007 13311
rect 25222 13308 25228 13320
rect 24995 13280 25228 13308
rect 24995 13277 25007 13280
rect 24949 13271 25007 13277
rect 17681 13243 17739 13249
rect 17681 13240 17693 13243
rect 14148 13212 17693 13240
rect 14148 13200 14154 13212
rect 17681 13209 17693 13212
rect 17727 13209 17739 13243
rect 17862 13240 17868 13252
rect 17823 13212 17868 13240
rect 17681 13203 17739 13209
rect 17862 13200 17868 13212
rect 17920 13200 17926 13252
rect 19797 13243 19855 13249
rect 19797 13240 19809 13243
rect 17972 13212 19809 13240
rect 6362 13172 6368 13184
rect 6323 13144 6368 13172
rect 6362 13132 6368 13144
rect 6420 13132 6426 13184
rect 6914 13132 6920 13184
rect 6972 13172 6978 13184
rect 7009 13175 7067 13181
rect 7009 13172 7021 13175
rect 6972 13144 7021 13172
rect 6972 13132 6978 13144
rect 7009 13141 7021 13144
rect 7055 13141 7067 13175
rect 7466 13172 7472 13184
rect 7427 13144 7472 13172
rect 7009 13135 7067 13141
rect 7466 13132 7472 13144
rect 7524 13132 7530 13184
rect 9030 13132 9036 13184
rect 9088 13172 9094 13184
rect 9490 13172 9496 13184
rect 9088 13144 9496 13172
rect 9088 13132 9094 13144
rect 9490 13132 9496 13144
rect 9548 13172 9554 13184
rect 9858 13172 9864 13184
rect 9548 13144 9864 13172
rect 9548 13132 9554 13144
rect 9858 13132 9864 13144
rect 9916 13132 9922 13184
rect 14461 13175 14519 13181
rect 14461 13141 14473 13175
rect 14507 13172 14519 13175
rect 14642 13172 14648 13184
rect 14507 13144 14648 13172
rect 14507 13141 14519 13144
rect 14461 13135 14519 13141
rect 14642 13132 14648 13144
rect 14700 13132 14706 13184
rect 17770 13132 17776 13184
rect 17828 13172 17834 13184
rect 17972 13172 18000 13212
rect 19797 13209 19809 13212
rect 19843 13209 19855 13243
rect 19797 13203 19855 13209
rect 19981 13243 20039 13249
rect 19981 13209 19993 13243
rect 20027 13240 20039 13243
rect 21361 13243 21419 13249
rect 21361 13240 21373 13243
rect 20027 13212 21373 13240
rect 20027 13209 20039 13212
rect 19981 13203 20039 13209
rect 21361 13209 21373 13212
rect 21407 13240 21419 13243
rect 22094 13240 22100 13252
rect 21407 13212 22100 13240
rect 21407 13209 21419 13212
rect 21361 13203 21419 13209
rect 22094 13200 22100 13212
rect 22152 13240 22158 13252
rect 23382 13240 23388 13252
rect 22152 13212 23388 13240
rect 22152 13200 22158 13212
rect 23382 13200 23388 13212
rect 23440 13200 23446 13252
rect 23477 13243 23535 13249
rect 23477 13209 23489 13243
rect 23523 13240 23535 13243
rect 23934 13240 23940 13252
rect 23523 13212 23940 13240
rect 23523 13209 23535 13212
rect 23477 13203 23535 13209
rect 23934 13200 23940 13212
rect 23992 13200 23998 13252
rect 17828 13144 18000 13172
rect 18049 13175 18107 13181
rect 17828 13132 17834 13144
rect 18049 13141 18061 13175
rect 18095 13172 18107 13175
rect 18506 13172 18512 13184
rect 18095 13144 18512 13172
rect 18095 13141 18107 13144
rect 18049 13135 18107 13141
rect 18506 13132 18512 13144
rect 18564 13132 18570 13184
rect 23106 13132 23112 13184
rect 23164 13172 23170 13184
rect 24780 13172 24808 13271
rect 25222 13268 25228 13280
rect 25280 13268 25286 13320
rect 27353 13317 27381 13416
rect 27522 13404 27528 13416
rect 27580 13404 27586 13456
rect 29638 13444 29644 13456
rect 29599 13416 29644 13444
rect 29638 13404 29644 13416
rect 29696 13404 29702 13456
rect 40402 13444 40408 13456
rect 38396 13416 40408 13444
rect 28169 13379 28227 13385
rect 28169 13345 28181 13379
rect 28215 13376 28227 13379
rect 29914 13376 29920 13388
rect 28215 13348 29920 13376
rect 28215 13345 28227 13348
rect 28169 13339 28227 13345
rect 27229 13311 27287 13317
rect 27229 13305 27241 13311
rect 27172 13277 27241 13305
rect 27275 13277 27287 13311
rect 27172 13240 27200 13277
rect 27229 13271 27287 13277
rect 27338 13311 27396 13317
rect 27338 13277 27350 13311
rect 27384 13277 27396 13311
rect 27338 13271 27396 13277
rect 27430 13268 27436 13320
rect 27488 13305 27494 13320
rect 27617 13311 27675 13317
rect 27488 13277 27530 13305
rect 27617 13277 27629 13311
rect 27663 13308 27675 13311
rect 27798 13308 27804 13320
rect 27663 13280 27804 13308
rect 27663 13277 27675 13280
rect 27488 13268 27494 13277
rect 27617 13271 27675 13277
rect 27798 13268 27804 13280
rect 27856 13308 27862 13320
rect 28074 13308 28080 13320
rect 27856 13280 28080 13308
rect 27856 13268 27862 13280
rect 28074 13268 28080 13280
rect 28132 13308 28138 13320
rect 28184 13308 28212 13339
rect 29914 13336 29920 13348
rect 29972 13336 29978 13388
rect 34149 13379 34207 13385
rect 34149 13345 34161 13379
rect 34195 13376 34207 13379
rect 35713 13379 35771 13385
rect 35713 13376 35725 13379
rect 34195 13348 35725 13376
rect 34195 13345 34207 13348
rect 34149 13339 34207 13345
rect 35713 13345 35725 13348
rect 35759 13345 35771 13379
rect 35713 13339 35771 13345
rect 28132 13280 28212 13308
rect 28132 13268 28138 13280
rect 29546 13268 29552 13320
rect 29604 13308 29610 13320
rect 31021 13311 31079 13317
rect 31021 13308 31033 13311
rect 29604 13280 31033 13308
rect 29604 13268 29610 13280
rect 31021 13277 31033 13280
rect 31067 13277 31079 13311
rect 31021 13271 31079 13277
rect 35069 13311 35127 13317
rect 35069 13277 35081 13311
rect 35115 13277 35127 13311
rect 35069 13271 35127 13277
rect 35253 13311 35311 13317
rect 35253 13277 35265 13311
rect 35299 13308 35311 13311
rect 35342 13308 35348 13320
rect 35299 13280 35348 13308
rect 35299 13277 35311 13280
rect 35253 13271 35311 13277
rect 26436 13212 27200 13240
rect 23164 13144 24808 13172
rect 23164 13132 23170 13144
rect 24854 13132 24860 13184
rect 24912 13172 24918 13184
rect 26436 13181 26464 13212
rect 29362 13200 29368 13252
rect 29420 13240 29426 13252
rect 30098 13240 30104 13252
rect 29420 13212 30104 13240
rect 29420 13200 29426 13212
rect 30098 13200 30104 13212
rect 30156 13200 30162 13252
rect 30742 13200 30748 13252
rect 30800 13249 30806 13252
rect 30800 13240 30812 13249
rect 31938 13240 31944 13252
rect 30800 13212 30845 13240
rect 31899 13212 31944 13240
rect 30800 13203 30812 13212
rect 30800 13200 30806 13203
rect 31938 13200 31944 13212
rect 31996 13200 32002 13252
rect 32122 13200 32128 13252
rect 32180 13240 32186 13252
rect 32180 13212 32812 13240
rect 32180 13200 32186 13212
rect 26421 13175 26479 13181
rect 26421 13172 26433 13175
rect 24912 13144 26433 13172
rect 24912 13132 24918 13144
rect 26421 13141 26433 13144
rect 26467 13141 26479 13175
rect 26421 13135 26479 13141
rect 29178 13132 29184 13184
rect 29236 13172 29242 13184
rect 29546 13172 29552 13184
rect 29236 13144 29552 13172
rect 29236 13132 29242 13144
rect 29546 13132 29552 13144
rect 29604 13132 29610 13184
rect 32309 13175 32367 13181
rect 32309 13141 32321 13175
rect 32355 13172 32367 13175
rect 32398 13172 32404 13184
rect 32355 13144 32404 13172
rect 32355 13141 32367 13144
rect 32309 13135 32367 13141
rect 32398 13132 32404 13144
rect 32456 13132 32462 13184
rect 32784 13181 32812 13212
rect 32950 13200 32956 13252
rect 33008 13240 33014 13252
rect 33882 13243 33940 13249
rect 33882 13240 33894 13243
rect 33008 13212 33894 13240
rect 33008 13200 33014 13212
rect 33882 13209 33894 13212
rect 33928 13209 33940 13243
rect 35084 13240 35112 13271
rect 35342 13268 35348 13280
rect 35400 13268 35406 13320
rect 35728 13308 35756 13339
rect 38396 13317 38424 13416
rect 40402 13404 40408 13416
rect 40460 13404 40466 13456
rect 38838 13376 38844 13388
rect 38672 13348 38844 13376
rect 38381 13311 38439 13317
rect 35728 13280 38332 13308
rect 35526 13240 35532 13252
rect 35084 13212 35532 13240
rect 33882 13203 33940 13209
rect 35526 13200 35532 13212
rect 35584 13200 35590 13252
rect 35618 13200 35624 13252
rect 35676 13240 35682 13252
rect 35958 13243 36016 13249
rect 35958 13240 35970 13243
rect 35676 13212 35970 13240
rect 35676 13200 35682 13212
rect 35958 13209 35970 13212
rect 36004 13209 36016 13243
rect 35958 13203 36016 13209
rect 32769 13175 32827 13181
rect 32769 13141 32781 13175
rect 32815 13141 32827 13175
rect 35250 13172 35256 13184
rect 35211 13144 35256 13172
rect 32769 13135 32827 13141
rect 35250 13132 35256 13144
rect 35308 13132 35314 13184
rect 36446 13132 36452 13184
rect 36504 13172 36510 13184
rect 37093 13175 37151 13181
rect 37093 13172 37105 13175
rect 36504 13144 37105 13172
rect 36504 13132 36510 13144
rect 37093 13141 37105 13144
rect 37139 13141 37151 13175
rect 38304 13172 38332 13280
rect 38381 13277 38393 13311
rect 38427 13277 38439 13311
rect 38562 13308 38568 13320
rect 38523 13280 38568 13308
rect 38381 13271 38439 13277
rect 38562 13268 38568 13280
rect 38620 13268 38626 13320
rect 38672 13317 38700 13348
rect 38838 13336 38844 13348
rect 38896 13376 38902 13388
rect 39022 13376 39028 13388
rect 38896 13348 39028 13376
rect 38896 13336 38902 13348
rect 39022 13336 39028 13348
rect 39080 13336 39086 13388
rect 38657 13311 38715 13317
rect 38657 13277 38669 13311
rect 38703 13277 38715 13311
rect 38657 13271 38715 13277
rect 38746 13268 38752 13320
rect 38804 13308 38810 13320
rect 39853 13311 39911 13317
rect 39853 13308 39865 13311
rect 38804 13280 39865 13308
rect 38804 13268 38810 13280
rect 39853 13277 39865 13280
rect 39899 13277 39911 13311
rect 58158 13308 58164 13320
rect 58119 13280 58164 13308
rect 39853 13271 39911 13277
rect 58158 13268 58164 13280
rect 58216 13268 58222 13320
rect 38654 13172 38660 13184
rect 38304 13144 38660 13172
rect 37093 13135 37151 13141
rect 38654 13132 38660 13144
rect 38712 13132 38718 13184
rect 39022 13172 39028 13184
rect 38983 13144 39028 13172
rect 39022 13132 39028 13144
rect 39080 13132 39086 13184
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 4617 12971 4675 12977
rect 4617 12968 4629 12971
rect 2746 12940 4629 12968
rect 2746 12900 2774 12940
rect 4617 12937 4629 12940
rect 4663 12937 4675 12971
rect 5074 12968 5080 12980
rect 5035 12940 5080 12968
rect 4617 12931 4675 12937
rect 5074 12928 5080 12940
rect 5132 12928 5138 12980
rect 14185 12971 14243 12977
rect 14185 12937 14197 12971
rect 14231 12968 14243 12971
rect 14274 12968 14280 12980
rect 14231 12940 14280 12968
rect 14231 12937 14243 12940
rect 14185 12931 14243 12937
rect 14274 12928 14280 12940
rect 14332 12928 14338 12980
rect 15746 12928 15752 12980
rect 15804 12968 15810 12980
rect 17037 12971 17095 12977
rect 17037 12968 17049 12971
rect 15804 12940 17049 12968
rect 15804 12928 15810 12940
rect 17037 12937 17049 12940
rect 17083 12968 17095 12971
rect 17862 12968 17868 12980
rect 17083 12940 17868 12968
rect 17083 12937 17095 12940
rect 17037 12931 17095 12937
rect 17862 12928 17868 12940
rect 17920 12928 17926 12980
rect 17972 12940 21128 12968
rect 2148 12872 2774 12900
rect 2148 12841 2176 12872
rect 6546 12860 6552 12912
rect 6604 12900 6610 12912
rect 7466 12900 7472 12912
rect 6604 12872 7472 12900
rect 6604 12860 6610 12872
rect 2133 12835 2191 12841
rect 2133 12801 2145 12835
rect 2179 12801 2191 12835
rect 2133 12795 2191 12801
rect 3044 12835 3102 12841
rect 3044 12801 3056 12835
rect 3090 12832 3102 12835
rect 3786 12832 3792 12844
rect 3090 12804 3792 12832
rect 3090 12801 3102 12804
rect 3044 12795 3102 12801
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 4614 12792 4620 12844
rect 4672 12832 4678 12844
rect 4798 12832 4804 12844
rect 4672 12804 4804 12832
rect 4672 12792 4678 12804
rect 4798 12792 4804 12804
rect 4856 12832 4862 12844
rect 6656 12841 6684 12872
rect 7466 12860 7472 12872
rect 7524 12860 7530 12912
rect 11517 12903 11575 12909
rect 11517 12900 11529 12903
rect 10428 12872 11529 12900
rect 4985 12835 5043 12841
rect 4985 12832 4997 12835
rect 4856 12804 4997 12832
rect 4856 12792 4862 12804
rect 4985 12801 4997 12804
rect 5031 12801 5043 12835
rect 4985 12795 5043 12801
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12801 6699 12835
rect 6822 12832 6828 12844
rect 6783 12804 6828 12832
rect 6641 12795 6699 12801
rect 6822 12792 6828 12804
rect 6880 12792 6886 12844
rect 6914 12792 6920 12844
rect 6972 12832 6978 12844
rect 7190 12832 7196 12844
rect 6972 12804 7017 12832
rect 7151 12804 7196 12832
rect 6972 12792 6978 12804
rect 7190 12792 7196 12804
rect 7248 12792 7254 12844
rect 8202 12792 8208 12844
rect 8260 12832 8266 12844
rect 10428 12841 10456 12872
rect 11517 12869 11529 12872
rect 11563 12900 11575 12903
rect 15381 12903 15439 12909
rect 15381 12900 15393 12903
rect 11563 12872 12434 12900
rect 11563 12869 11575 12872
rect 11517 12863 11575 12869
rect 8389 12835 8447 12841
rect 8389 12832 8401 12835
rect 8260 12804 8401 12832
rect 8260 12792 8266 12804
rect 8389 12801 8401 12804
rect 8435 12832 8447 12835
rect 10229 12835 10287 12841
rect 10229 12832 10241 12835
rect 8435 12804 10241 12832
rect 8435 12801 8447 12804
rect 8389 12795 8447 12801
rect 10229 12801 10241 12804
rect 10275 12801 10287 12835
rect 10229 12795 10287 12801
rect 10413 12835 10471 12841
rect 10413 12801 10425 12835
rect 10459 12801 10471 12835
rect 10413 12795 10471 12801
rect 10781 12835 10839 12841
rect 10781 12801 10793 12835
rect 10827 12832 10839 12835
rect 12158 12832 12164 12844
rect 10827 12804 12164 12832
rect 10827 12801 10839 12804
rect 10781 12795 10839 12801
rect 12158 12792 12164 12804
rect 12216 12792 12222 12844
rect 1949 12767 2007 12773
rect 1949 12733 1961 12767
rect 1995 12764 2007 12767
rect 2406 12764 2412 12776
rect 1995 12736 2412 12764
rect 1995 12733 2007 12736
rect 1949 12727 2007 12733
rect 2406 12724 2412 12736
rect 2464 12724 2470 12776
rect 2774 12724 2780 12776
rect 2832 12764 2838 12776
rect 5261 12767 5319 12773
rect 2832 12736 2877 12764
rect 2832 12724 2838 12736
rect 5261 12733 5273 12767
rect 5307 12764 5319 12767
rect 5350 12764 5356 12776
rect 5307 12736 5356 12764
rect 5307 12733 5319 12736
rect 5261 12727 5319 12733
rect 5350 12724 5356 12736
rect 5408 12724 5414 12776
rect 7009 12767 7067 12773
rect 7009 12733 7021 12767
rect 7055 12764 7067 12767
rect 7282 12764 7288 12776
rect 7055 12736 7288 12764
rect 7055 12733 7067 12736
rect 7009 12727 7067 12733
rect 7282 12724 7288 12736
rect 7340 12724 7346 12776
rect 8665 12767 8723 12773
rect 8665 12733 8677 12767
rect 8711 12733 8723 12767
rect 10502 12764 10508 12776
rect 10463 12736 10508 12764
rect 8665 12727 8723 12733
rect 3878 12656 3884 12708
rect 3936 12696 3942 12708
rect 8680 12696 8708 12727
rect 10502 12724 10508 12736
rect 10560 12724 10566 12776
rect 10597 12767 10655 12773
rect 10597 12733 10609 12767
rect 10643 12733 10655 12767
rect 10597 12727 10655 12733
rect 3936 12668 9536 12696
rect 3936 12656 3942 12668
rect 2317 12631 2375 12637
rect 2317 12597 2329 12631
rect 2363 12628 2375 12631
rect 2498 12628 2504 12640
rect 2363 12600 2504 12628
rect 2363 12597 2375 12600
rect 2317 12591 2375 12597
rect 2498 12588 2504 12600
rect 2556 12588 2562 12640
rect 4157 12631 4215 12637
rect 4157 12597 4169 12631
rect 4203 12628 4215 12631
rect 5258 12628 5264 12640
rect 4203 12600 5264 12628
rect 4203 12597 4215 12600
rect 4157 12591 4215 12597
rect 5258 12588 5264 12600
rect 5316 12588 5322 12640
rect 7377 12631 7435 12637
rect 7377 12597 7389 12631
rect 7423 12628 7435 12631
rect 8754 12628 8760 12640
rect 7423 12600 8760 12628
rect 7423 12597 7435 12600
rect 7377 12591 7435 12597
rect 8754 12588 8760 12600
rect 8812 12588 8818 12640
rect 9508 12628 9536 12668
rect 9582 12656 9588 12708
rect 9640 12696 9646 12708
rect 10612 12696 10640 12727
rect 11974 12696 11980 12708
rect 9640 12668 10640 12696
rect 10888 12668 11980 12696
rect 9640 12656 9646 12668
rect 10888 12628 10916 12668
rect 11974 12656 11980 12668
rect 12032 12656 12038 12708
rect 9508 12600 10916 12628
rect 10965 12631 11023 12637
rect 10965 12597 10977 12631
rect 11011 12628 11023 12631
rect 11054 12628 11060 12640
rect 11011 12600 11060 12628
rect 11011 12597 11023 12600
rect 10965 12591 11023 12597
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 12406 12628 12434 12872
rect 14476 12872 15393 12900
rect 14476 12844 14504 12872
rect 15381 12869 15393 12872
rect 15427 12900 15439 12903
rect 17972 12900 18000 12940
rect 15427 12872 18000 12900
rect 15427 12869 15439 12872
rect 15381 12863 15439 12869
rect 20254 12860 20260 12912
rect 20312 12900 20318 12912
rect 20993 12903 21051 12909
rect 20993 12900 21005 12903
rect 20312 12872 21005 12900
rect 20312 12860 20318 12872
rect 20993 12869 21005 12872
rect 21039 12869 21051 12903
rect 21100 12900 21128 12940
rect 22066 12940 25176 12968
rect 22066 12900 22094 12940
rect 24857 12903 24915 12909
rect 24857 12900 24869 12903
rect 21100 12872 22094 12900
rect 24136 12872 24869 12900
rect 20993 12863 21051 12869
rect 24136 12844 24164 12872
rect 24857 12869 24869 12872
rect 24903 12900 24915 12903
rect 24946 12900 24952 12912
rect 24903 12872 24952 12900
rect 24903 12869 24915 12872
rect 24857 12863 24915 12869
rect 24946 12860 24952 12872
rect 25004 12860 25010 12912
rect 25148 12900 25176 12940
rect 25222 12928 25228 12980
rect 25280 12968 25286 12980
rect 25317 12971 25375 12977
rect 25317 12968 25329 12971
rect 25280 12940 25329 12968
rect 25280 12928 25286 12940
rect 25317 12937 25329 12940
rect 25363 12937 25375 12971
rect 27798 12968 27804 12980
rect 27759 12940 27804 12968
rect 25317 12931 25375 12937
rect 27798 12928 27804 12940
rect 27856 12928 27862 12980
rect 29546 12928 29552 12980
rect 29604 12968 29610 12980
rect 29641 12971 29699 12977
rect 29641 12968 29653 12971
rect 29604 12940 29653 12968
rect 29604 12928 29610 12940
rect 29641 12937 29653 12940
rect 29687 12937 29699 12971
rect 31570 12968 31576 12980
rect 31483 12940 31576 12968
rect 29641 12931 29699 12937
rect 29086 12900 29092 12912
rect 25148 12872 29092 12900
rect 29086 12860 29092 12872
rect 29144 12860 29150 12912
rect 29656 12900 29684 12931
rect 31496 12909 31524 12940
rect 31570 12928 31576 12940
rect 31628 12968 31634 12980
rect 32950 12968 32956 12980
rect 31628 12940 32720 12968
rect 32911 12940 32956 12968
rect 31628 12928 31634 12940
rect 30285 12903 30343 12909
rect 30285 12900 30297 12903
rect 29656 12872 30297 12900
rect 30285 12869 30297 12872
rect 30331 12869 30343 12903
rect 30285 12863 30343 12869
rect 30469 12903 30527 12909
rect 30469 12869 30481 12903
rect 30515 12900 30527 12903
rect 31481 12903 31539 12909
rect 31481 12900 31493 12903
rect 30515 12872 31493 12900
rect 30515 12869 30527 12872
rect 30469 12863 30527 12869
rect 31481 12869 31493 12872
rect 31527 12869 31539 12903
rect 31481 12863 31539 12869
rect 14458 12832 14464 12844
rect 14371 12804 14464 12832
rect 14458 12792 14464 12804
rect 14516 12792 14522 12844
rect 14553 12835 14611 12841
rect 14553 12801 14565 12835
rect 14599 12801 14611 12835
rect 14553 12795 14611 12801
rect 14568 12764 14596 12795
rect 14642 12792 14648 12844
rect 14700 12832 14706 12844
rect 14829 12835 14887 12841
rect 14700 12804 14745 12832
rect 14700 12792 14706 12804
rect 14829 12801 14841 12835
rect 14875 12832 14887 12835
rect 15102 12832 15108 12844
rect 14875 12804 15108 12832
rect 14875 12801 14887 12804
rect 14829 12795 14887 12801
rect 15102 12792 15108 12804
rect 15160 12792 15166 12844
rect 18138 12832 18144 12844
rect 18196 12841 18202 12844
rect 18108 12804 18144 12832
rect 18138 12792 18144 12804
rect 18196 12795 18208 12841
rect 18196 12792 18202 12795
rect 18322 12792 18328 12844
rect 18380 12832 18386 12844
rect 18417 12835 18475 12841
rect 18417 12832 18429 12835
rect 18380 12804 18429 12832
rect 18380 12792 18386 12804
rect 18417 12801 18429 12804
rect 18463 12801 18475 12835
rect 19150 12832 19156 12844
rect 19111 12804 19156 12832
rect 18417 12795 18475 12801
rect 19150 12792 19156 12804
rect 19208 12792 19214 12844
rect 19245 12835 19303 12841
rect 19245 12801 19257 12835
rect 19291 12801 19303 12835
rect 19245 12795 19303 12801
rect 19337 12835 19395 12841
rect 19337 12801 19349 12835
rect 19383 12801 19395 12835
rect 19337 12795 19395 12801
rect 19533 12835 19591 12841
rect 19533 12801 19545 12835
rect 19579 12832 19591 12835
rect 20349 12835 20407 12841
rect 19579 12804 20300 12832
rect 19579 12801 19591 12804
rect 19533 12795 19591 12801
rect 14918 12764 14924 12776
rect 14568 12736 14924 12764
rect 14918 12724 14924 12736
rect 14976 12724 14982 12776
rect 18414 12656 18420 12708
rect 18472 12696 18478 12708
rect 19260 12696 19288 12795
rect 19352 12708 19380 12795
rect 20272 12764 20300 12804
rect 20349 12801 20361 12835
rect 20395 12832 20407 12835
rect 20809 12835 20867 12841
rect 20809 12832 20821 12835
rect 20395 12804 20821 12832
rect 20395 12801 20407 12804
rect 20349 12795 20407 12801
rect 20809 12801 20821 12804
rect 20855 12832 20867 12835
rect 20898 12832 20904 12844
rect 20855 12804 20904 12832
rect 20855 12801 20867 12804
rect 20809 12795 20867 12801
rect 20898 12792 20904 12804
rect 20956 12792 20962 12844
rect 22094 12792 22100 12844
rect 22152 12832 22158 12844
rect 24118 12832 24124 12844
rect 22152 12804 22197 12832
rect 24079 12804 24124 12832
rect 22152 12792 22158 12804
rect 24118 12792 24124 12804
rect 24176 12792 24182 12844
rect 24670 12832 24676 12844
rect 24631 12804 24676 12832
rect 24670 12792 24676 12804
rect 24728 12792 24734 12844
rect 31294 12792 31300 12844
rect 31352 12832 31358 12844
rect 32297 12835 32355 12841
rect 32232 12832 32309 12835
rect 31352 12807 32309 12832
rect 31352 12804 32260 12807
rect 31352 12792 31358 12804
rect 32297 12801 32309 12807
rect 32343 12801 32355 12835
rect 32297 12795 32355 12801
rect 32398 12792 32404 12844
rect 32456 12832 32462 12844
rect 32692 12841 32720 12940
rect 32950 12928 32956 12940
rect 33008 12928 33014 12980
rect 34977 12971 35035 12977
rect 34977 12937 34989 12971
rect 35023 12968 35035 12971
rect 35342 12968 35348 12980
rect 35023 12940 35348 12968
rect 35023 12937 35035 12940
rect 34977 12931 35035 12937
rect 35342 12928 35348 12940
rect 35400 12928 35406 12980
rect 35618 12968 35624 12980
rect 35579 12940 35624 12968
rect 35618 12928 35624 12940
rect 35676 12928 35682 12980
rect 38378 12928 38384 12980
rect 38436 12968 38442 12980
rect 39945 12971 40003 12977
rect 39945 12968 39957 12971
rect 38436 12940 39957 12968
rect 38436 12928 38442 12940
rect 39945 12937 39957 12940
rect 39991 12937 40003 12971
rect 39945 12931 40003 12937
rect 35250 12860 35256 12912
rect 35308 12900 35314 12912
rect 38832 12903 38890 12909
rect 35308 12872 38792 12900
rect 35308 12860 35314 12872
rect 32493 12835 32551 12841
rect 32493 12832 32505 12835
rect 32456 12804 32505 12832
rect 32456 12792 32462 12804
rect 32493 12801 32505 12804
rect 32539 12801 32551 12835
rect 32493 12795 32551 12801
rect 32588 12835 32646 12841
rect 32588 12801 32600 12835
rect 32634 12801 32646 12835
rect 32588 12795 32646 12801
rect 32677 12835 32735 12841
rect 32677 12801 32689 12835
rect 32723 12801 32735 12835
rect 35894 12832 35900 12844
rect 35855 12804 35900 12832
rect 32677 12795 32735 12801
rect 20530 12764 20536 12776
rect 20272 12736 20536 12764
rect 20530 12724 20536 12736
rect 20588 12724 20594 12776
rect 23845 12767 23903 12773
rect 23845 12733 23857 12767
rect 23891 12764 23903 12767
rect 24026 12764 24032 12776
rect 23891 12736 24032 12764
rect 23891 12733 23903 12736
rect 23845 12727 23903 12733
rect 24026 12724 24032 12736
rect 24084 12724 24090 12776
rect 24302 12724 24308 12776
rect 24360 12764 24366 12776
rect 24360 12736 31754 12764
rect 24360 12724 24366 12736
rect 18472 12668 19288 12696
rect 18472 12656 18478 12668
rect 17678 12628 17684 12640
rect 12406 12600 17684 12628
rect 17678 12588 17684 12600
rect 17736 12588 17742 12640
rect 18874 12628 18880 12640
rect 18835 12600 18880 12628
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 19260 12628 19288 12668
rect 19334 12656 19340 12708
rect 19392 12656 19398 12708
rect 19426 12656 19432 12708
rect 19484 12696 19490 12708
rect 20165 12699 20223 12705
rect 20165 12696 20177 12699
rect 19484 12668 20177 12696
rect 19484 12656 19490 12668
rect 20165 12665 20177 12668
rect 20211 12665 20223 12699
rect 20165 12659 20223 12665
rect 24578 12656 24584 12708
rect 24636 12696 24642 12708
rect 31726 12696 31754 12736
rect 31846 12724 31852 12776
rect 31904 12764 31910 12776
rect 32603 12764 32631 12795
rect 35894 12792 35900 12804
rect 35952 12792 35958 12844
rect 36004 12841 36032 12872
rect 35989 12835 36047 12841
rect 35989 12801 36001 12835
rect 36035 12801 36047 12835
rect 35989 12795 36047 12801
rect 36078 12792 36084 12844
rect 36136 12832 36142 12844
rect 36136 12804 36181 12832
rect 36136 12792 36142 12804
rect 36262 12792 36268 12844
rect 36320 12832 36326 12844
rect 38565 12835 38623 12841
rect 36320 12804 36365 12832
rect 36320 12792 36326 12804
rect 38565 12801 38577 12835
rect 38611 12832 38623 12835
rect 38654 12832 38660 12844
rect 38611 12804 38660 12832
rect 38611 12801 38623 12804
rect 38565 12795 38623 12801
rect 38654 12792 38660 12804
rect 38712 12792 38718 12844
rect 38764 12832 38792 12872
rect 38832 12869 38844 12903
rect 38878 12900 38890 12903
rect 39022 12900 39028 12912
rect 38878 12872 39028 12900
rect 38878 12869 38890 12872
rect 38832 12863 38890 12869
rect 39022 12860 39028 12872
rect 39080 12860 39086 12912
rect 39206 12832 39212 12844
rect 38764 12804 39212 12832
rect 39206 12792 39212 12804
rect 39264 12792 39270 12844
rect 31904 12736 32631 12764
rect 31904 12724 31910 12736
rect 34606 12696 34612 12708
rect 24636 12668 31616 12696
rect 31726 12668 34612 12696
rect 24636 12656 24642 12668
rect 20806 12628 20812 12640
rect 19260 12600 20812 12628
rect 20806 12588 20812 12600
rect 20864 12588 20870 12640
rect 21177 12631 21235 12637
rect 21177 12597 21189 12631
rect 21223 12628 21235 12631
rect 22002 12628 22008 12640
rect 21223 12600 22008 12628
rect 21223 12597 21235 12600
rect 21177 12591 21235 12597
rect 22002 12588 22008 12600
rect 22060 12588 22066 12640
rect 27062 12628 27068 12640
rect 27023 12600 27068 12628
rect 27062 12588 27068 12600
rect 27120 12588 27126 12640
rect 31588 12628 31616 12668
rect 34606 12656 34612 12668
rect 34664 12656 34670 12708
rect 34698 12628 34704 12640
rect 31588 12600 34704 12628
rect 34698 12588 34704 12600
rect 34756 12588 34762 12640
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 7098 12424 7104 12436
rect 2832 12396 7104 12424
rect 2832 12384 2838 12396
rect 7098 12384 7104 12396
rect 7156 12424 7162 12436
rect 7926 12424 7932 12436
rect 7156 12396 7932 12424
rect 7156 12384 7162 12396
rect 7926 12384 7932 12396
rect 7984 12384 7990 12436
rect 14826 12424 14832 12436
rect 9508 12396 14832 12424
rect 9508 12368 9536 12396
rect 14826 12384 14832 12396
rect 14884 12384 14890 12436
rect 19245 12427 19303 12433
rect 19245 12393 19257 12427
rect 19291 12424 19303 12427
rect 19334 12424 19340 12436
rect 19291 12396 19340 12424
rect 19291 12393 19303 12396
rect 19245 12387 19303 12393
rect 19334 12384 19340 12396
rect 19392 12384 19398 12436
rect 22554 12384 22560 12436
rect 22612 12424 22618 12436
rect 22649 12427 22707 12433
rect 22649 12424 22661 12427
rect 22612 12396 22661 12424
rect 22612 12384 22618 12396
rect 22649 12393 22661 12396
rect 22695 12393 22707 12427
rect 22649 12387 22707 12393
rect 23661 12427 23719 12433
rect 23661 12393 23673 12427
rect 23707 12424 23719 12427
rect 23934 12424 23940 12436
rect 23707 12396 23940 12424
rect 23707 12393 23719 12396
rect 23661 12387 23719 12393
rect 23934 12384 23940 12396
rect 23992 12384 23998 12436
rect 24946 12424 24952 12436
rect 24907 12396 24952 12424
rect 24946 12384 24952 12396
rect 25004 12384 25010 12436
rect 29730 12384 29736 12436
rect 29788 12424 29794 12436
rect 30745 12427 30803 12433
rect 30745 12424 30757 12427
rect 29788 12396 30757 12424
rect 29788 12384 29794 12396
rect 30745 12393 30757 12396
rect 30791 12424 30803 12427
rect 30791 12396 31708 12424
rect 30791 12393 30803 12396
rect 30745 12387 30803 12393
rect 9490 12316 9496 12368
rect 9548 12316 9554 12368
rect 12158 12356 12164 12368
rect 12071 12328 12164 12356
rect 12158 12316 12164 12328
rect 12216 12356 12222 12368
rect 13722 12356 13728 12368
rect 12216 12328 13728 12356
rect 12216 12316 12222 12328
rect 13722 12316 13728 12328
rect 13780 12316 13786 12368
rect 28166 12356 28172 12368
rect 28127 12328 28172 12356
rect 28166 12316 28172 12328
rect 28224 12316 28230 12368
rect 31680 12356 31708 12396
rect 37642 12384 37648 12436
rect 37700 12424 37706 12436
rect 37918 12424 37924 12436
rect 37700 12396 37924 12424
rect 37700 12384 37706 12396
rect 37918 12384 37924 12396
rect 37976 12384 37982 12436
rect 31680 12328 31728 12356
rect 5350 12288 5356 12300
rect 5311 12260 5356 12288
rect 5350 12248 5356 12260
rect 5408 12248 5414 12300
rect 12434 12248 12440 12300
rect 12492 12288 12498 12300
rect 13262 12288 13268 12300
rect 12492 12260 13268 12288
rect 12492 12248 12498 12260
rect 13262 12248 13268 12260
rect 13320 12288 13326 12300
rect 16666 12288 16672 12300
rect 13320 12260 16672 12288
rect 13320 12248 13326 12260
rect 16666 12248 16672 12260
rect 16724 12248 16730 12300
rect 19426 12248 19432 12300
rect 19484 12248 19490 12300
rect 20806 12288 20812 12300
rect 20767 12260 20812 12288
rect 20806 12248 20812 12260
rect 20864 12248 20870 12300
rect 21082 12288 21088 12300
rect 21043 12260 21088 12288
rect 21082 12248 21088 12260
rect 21140 12288 21146 12300
rect 21140 12260 21947 12288
rect 21140 12248 21146 12260
rect 2498 12220 2504 12232
rect 2459 12192 2504 12220
rect 2498 12180 2504 12192
rect 2556 12180 2562 12232
rect 7926 12180 7932 12232
rect 7984 12220 7990 12232
rect 11054 12229 11060 12232
rect 10781 12223 10839 12229
rect 10781 12220 10793 12223
rect 7984 12192 10793 12220
rect 7984 12180 7990 12192
rect 10781 12189 10793 12192
rect 10827 12189 10839 12223
rect 10781 12183 10839 12189
rect 11048 12183 11060 12229
rect 11112 12220 11118 12232
rect 13541 12223 13599 12229
rect 11112 12192 11148 12220
rect 11054 12180 11060 12183
rect 11112 12180 11118 12192
rect 13541 12189 13553 12223
rect 13587 12220 13599 12223
rect 14090 12220 14096 12232
rect 13587 12192 14096 12220
rect 13587 12189 13599 12192
rect 13541 12183 13599 12189
rect 14090 12180 14096 12192
rect 14148 12180 14154 12232
rect 14645 12223 14703 12229
rect 14645 12189 14657 12223
rect 14691 12189 14703 12223
rect 14645 12183 14703 12189
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12189 14795 12223
rect 14737 12183 14795 12189
rect 5166 12152 5172 12164
rect 4632 12124 5172 12152
rect 4632 12096 4660 12124
rect 5166 12112 5172 12124
rect 5224 12112 5230 12164
rect 5810 12112 5816 12164
rect 5868 12152 5874 12164
rect 6641 12155 6699 12161
rect 6641 12152 6653 12155
rect 5868 12124 6653 12152
rect 5868 12112 5874 12124
rect 6641 12121 6653 12124
rect 6687 12152 6699 12155
rect 8941 12155 8999 12161
rect 8941 12152 8953 12155
rect 6687 12124 8953 12152
rect 6687 12121 6699 12124
rect 6641 12115 6699 12121
rect 8941 12121 8953 12124
rect 8987 12152 8999 12155
rect 9674 12152 9680 12164
rect 8987 12124 9680 12152
rect 8987 12121 8999 12124
rect 8941 12115 8999 12121
rect 9674 12112 9680 12124
rect 9732 12112 9738 12164
rect 13354 12152 13360 12164
rect 13315 12124 13360 12152
rect 13354 12112 13360 12124
rect 13412 12112 13418 12164
rect 2682 12084 2688 12096
rect 2643 12056 2688 12084
rect 2682 12044 2688 12056
rect 2740 12044 2746 12096
rect 4341 12087 4399 12093
rect 4341 12053 4353 12087
rect 4387 12084 4399 12087
rect 4614 12084 4620 12096
rect 4387 12056 4620 12084
rect 4387 12053 4399 12056
rect 4341 12047 4399 12053
rect 4614 12044 4620 12056
rect 4672 12044 4678 12096
rect 4801 12087 4859 12093
rect 4801 12053 4813 12087
rect 4847 12084 4859 12087
rect 4890 12084 4896 12096
rect 4847 12056 4896 12084
rect 4847 12053 4859 12056
rect 4801 12047 4859 12053
rect 4890 12044 4896 12056
rect 4948 12044 4954 12096
rect 5258 12044 5264 12096
rect 5316 12084 5322 12096
rect 13173 12087 13231 12093
rect 5316 12056 5361 12084
rect 5316 12044 5322 12056
rect 13173 12053 13185 12087
rect 13219 12084 13231 12087
rect 14274 12084 14280 12096
rect 13219 12056 14280 12084
rect 13219 12053 13231 12056
rect 13173 12047 13231 12053
rect 14274 12044 14280 12056
rect 14332 12044 14338 12096
rect 14366 12044 14372 12096
rect 14424 12084 14430 12096
rect 14660 12084 14688 12183
rect 14752 12152 14780 12183
rect 14826 12180 14832 12232
rect 14884 12220 14890 12232
rect 15013 12223 15071 12229
rect 14884 12192 14929 12220
rect 14884 12180 14890 12192
rect 15013 12189 15025 12223
rect 15059 12220 15071 12223
rect 15102 12220 15108 12232
rect 15059 12192 15108 12220
rect 15059 12189 15071 12192
rect 15013 12183 15071 12189
rect 15102 12180 15108 12192
rect 15160 12180 15166 12232
rect 15470 12180 15476 12232
rect 15528 12220 15534 12232
rect 18417 12223 18475 12229
rect 18417 12220 18429 12223
rect 15528 12192 18429 12220
rect 15528 12180 15534 12192
rect 18417 12189 18429 12192
rect 18463 12189 18475 12223
rect 19444 12220 19472 12248
rect 19613 12223 19671 12229
rect 19613 12220 19625 12223
rect 19444 12192 19625 12220
rect 18417 12183 18475 12189
rect 19613 12189 19625 12192
rect 19659 12189 19671 12223
rect 21818 12220 21824 12232
rect 21779 12192 21824 12220
rect 19613 12183 19671 12189
rect 21818 12180 21824 12192
rect 21876 12180 21882 12232
rect 21919 12229 21947 12260
rect 21910 12223 21968 12229
rect 21910 12189 21922 12223
rect 21956 12189 21968 12223
rect 21910 12183 21968 12189
rect 22002 12180 22008 12232
rect 22060 12220 22066 12232
rect 22189 12223 22247 12229
rect 22060 12192 22105 12220
rect 22060 12180 22066 12192
rect 22189 12189 22201 12223
rect 22235 12220 22247 12223
rect 22554 12220 22560 12232
rect 22235 12192 22560 12220
rect 22235 12189 22247 12192
rect 22189 12183 22247 12189
rect 22554 12180 22560 12192
rect 22612 12220 22618 12232
rect 24946 12220 24952 12232
rect 22612 12192 24952 12220
rect 22612 12180 22618 12192
rect 24946 12180 24952 12192
rect 25004 12180 25010 12232
rect 25038 12180 25044 12232
rect 25096 12220 25102 12232
rect 25406 12220 25412 12232
rect 25096 12192 25412 12220
rect 25096 12180 25102 12192
rect 25406 12180 25412 12192
rect 25464 12220 25470 12232
rect 25501 12223 25559 12229
rect 25501 12220 25513 12223
rect 25464 12192 25513 12220
rect 25464 12180 25470 12192
rect 25501 12189 25513 12192
rect 25547 12189 25559 12223
rect 31294 12220 31300 12232
rect 31255 12192 31300 12220
rect 25501 12183 25559 12189
rect 31294 12180 31300 12192
rect 31352 12180 31358 12232
rect 31478 12220 31484 12232
rect 31439 12192 31484 12220
rect 31478 12180 31484 12192
rect 31536 12180 31542 12232
rect 31700 12229 31728 12328
rect 37274 12288 37280 12300
rect 33704 12260 37280 12288
rect 31592 12223 31650 12229
rect 31592 12220 31604 12223
rect 31591 12189 31604 12220
rect 31638 12189 31650 12223
rect 31591 12183 31650 12189
rect 31685 12223 31743 12229
rect 31685 12189 31697 12223
rect 31731 12189 31743 12223
rect 31685 12183 31743 12189
rect 14918 12152 14924 12164
rect 14752 12124 14924 12152
rect 14918 12112 14924 12124
rect 14976 12112 14982 12164
rect 18172 12155 18230 12161
rect 18172 12121 18184 12155
rect 18218 12152 18230 12155
rect 18874 12152 18880 12164
rect 18218 12124 18880 12152
rect 18218 12121 18230 12124
rect 18172 12115 18230 12121
rect 18874 12112 18880 12124
rect 18932 12112 18938 12164
rect 19429 12155 19487 12161
rect 19429 12121 19441 12155
rect 19475 12121 19487 12155
rect 19429 12115 19487 12121
rect 14826 12084 14832 12096
rect 14424 12056 14469 12084
rect 14660 12056 14832 12084
rect 14424 12044 14430 12056
rect 14826 12044 14832 12056
rect 14884 12084 14890 12096
rect 15473 12087 15531 12093
rect 15473 12084 15485 12087
rect 14884 12056 15485 12084
rect 14884 12044 14890 12056
rect 15473 12053 15485 12056
rect 15519 12053 15531 12087
rect 15473 12047 15531 12053
rect 16942 12044 16948 12096
rect 17000 12084 17006 12096
rect 17037 12087 17095 12093
rect 17037 12084 17049 12087
rect 17000 12056 17049 12084
rect 17000 12044 17006 12056
rect 17037 12053 17049 12056
rect 17083 12084 17095 12087
rect 19444 12084 19472 12115
rect 20162 12112 20168 12164
rect 20220 12152 20226 12164
rect 20220 12124 22094 12152
rect 20220 12112 20226 12124
rect 21542 12084 21548 12096
rect 17083 12056 19472 12084
rect 21503 12056 21548 12084
rect 17083 12053 17095 12056
rect 17037 12047 17095 12053
rect 21542 12044 21548 12056
rect 21600 12044 21606 12096
rect 22066 12084 22094 12124
rect 25590 12112 25596 12164
rect 25648 12152 25654 12164
rect 25746 12155 25804 12161
rect 25746 12152 25758 12155
rect 25648 12124 25758 12152
rect 25648 12112 25654 12124
rect 25746 12121 25758 12124
rect 25792 12121 25804 12155
rect 25746 12115 25804 12121
rect 27617 12155 27675 12161
rect 27617 12121 27629 12155
rect 27663 12152 27675 12155
rect 28350 12152 28356 12164
rect 27663 12124 28356 12152
rect 27663 12121 27675 12124
rect 27617 12115 27675 12121
rect 28350 12112 28356 12124
rect 28408 12112 28414 12164
rect 31591 12152 31619 12183
rect 32030 12180 32036 12232
rect 32088 12220 32094 12232
rect 33704 12220 33732 12260
rect 37274 12248 37280 12260
rect 37332 12248 37338 12300
rect 37458 12248 37464 12300
rect 37516 12288 37522 12300
rect 38197 12291 38255 12297
rect 38197 12288 38209 12291
rect 37516 12260 38209 12288
rect 37516 12248 37522 12260
rect 38197 12257 38209 12260
rect 38243 12257 38255 12291
rect 38197 12251 38255 12257
rect 32088 12192 33732 12220
rect 33781 12223 33839 12229
rect 32088 12180 32094 12192
rect 33781 12189 33793 12223
rect 33827 12220 33839 12223
rect 34790 12220 34796 12232
rect 33827 12192 34796 12220
rect 33827 12189 33839 12192
rect 33781 12183 33839 12189
rect 34790 12180 34796 12192
rect 34848 12180 34854 12232
rect 37550 12180 37556 12232
rect 37608 12220 37614 12232
rect 37921 12223 37979 12229
rect 37921 12220 37933 12223
rect 37608 12192 37933 12220
rect 37608 12180 37614 12192
rect 37921 12189 37933 12192
rect 37967 12189 37979 12223
rect 37921 12183 37979 12189
rect 31846 12152 31852 12164
rect 31591 12124 31852 12152
rect 31846 12112 31852 12124
rect 31904 12112 31910 12164
rect 31941 12155 31999 12161
rect 31941 12121 31953 12155
rect 31987 12152 31999 12155
rect 33514 12155 33572 12161
rect 33514 12152 33526 12155
rect 31987 12124 33526 12152
rect 31987 12121 31999 12124
rect 31941 12115 31999 12121
rect 33514 12121 33526 12124
rect 33560 12121 33572 12155
rect 33514 12115 33572 12121
rect 35342 12112 35348 12164
rect 35400 12152 35406 12164
rect 35526 12152 35532 12164
rect 35400 12124 35532 12152
rect 35400 12112 35406 12124
rect 35526 12112 35532 12124
rect 35584 12112 35590 12164
rect 24486 12084 24492 12096
rect 22066 12056 24492 12084
rect 24486 12044 24492 12056
rect 24544 12044 24550 12096
rect 25958 12044 25964 12096
rect 26016 12084 26022 12096
rect 26881 12087 26939 12093
rect 26881 12084 26893 12087
rect 26016 12056 26893 12084
rect 26016 12044 26022 12056
rect 26881 12053 26893 12056
rect 26927 12053 26939 12087
rect 27522 12084 27528 12096
rect 27483 12056 27528 12084
rect 26881 12047 26939 12053
rect 27522 12044 27528 12056
rect 27580 12044 27586 12096
rect 27706 12044 27712 12096
rect 27764 12084 27770 12096
rect 32030 12084 32036 12096
rect 27764 12056 32036 12084
rect 27764 12044 27770 12056
rect 32030 12044 32036 12056
rect 32088 12044 32094 12096
rect 32398 12084 32404 12096
rect 32359 12056 32404 12084
rect 32398 12044 32404 12056
rect 32456 12044 32462 12096
rect 35250 12044 35256 12096
rect 35308 12084 35314 12096
rect 35437 12087 35495 12093
rect 35437 12084 35449 12087
rect 35308 12056 35449 12084
rect 35308 12044 35314 12056
rect 35437 12053 35449 12056
rect 35483 12084 35495 12087
rect 35894 12084 35900 12096
rect 35483 12056 35900 12084
rect 35483 12053 35495 12056
rect 35437 12047 35495 12053
rect 35894 12044 35900 12056
rect 35952 12044 35958 12096
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 4249 11883 4307 11889
rect 4249 11849 4261 11883
rect 4295 11880 4307 11883
rect 5074 11880 5080 11892
rect 4295 11852 5080 11880
rect 4295 11849 4307 11852
rect 4249 11843 4307 11849
rect 5074 11840 5080 11852
rect 5132 11840 5138 11892
rect 14001 11883 14059 11889
rect 14001 11849 14013 11883
rect 14047 11880 14059 11883
rect 14734 11880 14740 11892
rect 14047 11852 14740 11880
rect 14047 11849 14059 11852
rect 14001 11843 14059 11849
rect 14734 11840 14740 11852
rect 14792 11840 14798 11892
rect 14918 11880 14924 11892
rect 14844 11852 14924 11880
rect 2682 11772 2688 11824
rect 2740 11812 2746 11824
rect 3114 11815 3172 11821
rect 3114 11812 3126 11815
rect 2740 11784 3126 11812
rect 2740 11772 2746 11784
rect 3114 11781 3126 11784
rect 3160 11781 3172 11815
rect 3114 11775 3172 11781
rect 7926 11772 7932 11824
rect 7984 11812 7990 11824
rect 13633 11815 13691 11821
rect 7984 11784 9076 11812
rect 7984 11772 7990 11784
rect 2774 11704 2780 11756
rect 2832 11744 2838 11756
rect 2869 11747 2927 11753
rect 2869 11744 2881 11747
rect 2832 11716 2881 11744
rect 2832 11704 2838 11716
rect 2869 11713 2881 11716
rect 2915 11713 2927 11747
rect 4890 11744 4896 11756
rect 4851 11716 4896 11744
rect 2869 11707 2927 11713
rect 4890 11704 4896 11716
rect 4948 11704 4954 11756
rect 6638 11744 6644 11756
rect 6599 11716 6644 11744
rect 6638 11704 6644 11716
rect 6696 11704 6702 11756
rect 8754 11704 8760 11756
rect 8812 11753 8818 11756
rect 9048 11753 9076 11784
rect 13633 11781 13645 11815
rect 13679 11812 13691 11815
rect 14090 11812 14096 11824
rect 13679 11784 14096 11812
rect 13679 11781 13691 11784
rect 13633 11775 13691 11781
rect 14090 11772 14096 11784
rect 14148 11772 14154 11824
rect 14274 11772 14280 11824
rect 14332 11812 14338 11824
rect 14844 11812 14872 11852
rect 14918 11840 14924 11852
rect 14976 11840 14982 11892
rect 18049 11883 18107 11889
rect 18049 11849 18061 11883
rect 18095 11880 18107 11883
rect 18138 11880 18144 11892
rect 18095 11852 18144 11880
rect 18095 11849 18107 11852
rect 18049 11843 18107 11849
rect 18138 11840 18144 11852
rect 18196 11840 18202 11892
rect 18230 11840 18236 11892
rect 18288 11880 18294 11892
rect 19889 11883 19947 11889
rect 18288 11852 19564 11880
rect 18288 11840 18294 11852
rect 14332 11784 14872 11812
rect 17497 11815 17555 11821
rect 14332 11772 14338 11784
rect 17497 11781 17509 11815
rect 17543 11812 17555 11815
rect 19536 11812 19564 11852
rect 19889 11849 19901 11883
rect 19935 11880 19947 11883
rect 20254 11880 20260 11892
rect 19935 11852 20260 11880
rect 19935 11849 19947 11852
rect 19889 11843 19947 11849
rect 20254 11840 20260 11852
rect 20312 11840 20318 11892
rect 21174 11840 21180 11892
rect 21232 11880 21238 11892
rect 22462 11880 22468 11892
rect 21232 11852 22468 11880
rect 21232 11840 21238 11852
rect 22462 11840 22468 11852
rect 22520 11840 22526 11892
rect 23566 11880 23572 11892
rect 22572 11852 23572 11880
rect 20162 11812 20168 11824
rect 17543 11784 19334 11812
rect 19536 11784 20168 11812
rect 17543 11781 17555 11784
rect 17497 11775 17555 11781
rect 8812 11744 8824 11753
rect 9033 11747 9091 11753
rect 8812 11716 8857 11744
rect 8812 11707 8824 11716
rect 9033 11713 9045 11747
rect 9079 11713 9091 11747
rect 9033 11707 9091 11713
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11744 11851 11747
rect 11974 11744 11980 11756
rect 11839 11716 11980 11744
rect 11839 11713 11851 11716
rect 11793 11707 11851 11713
rect 8812 11704 8818 11707
rect 11974 11704 11980 11716
rect 12032 11704 12038 11756
rect 13814 11704 13820 11756
rect 13872 11744 13878 11756
rect 13998 11744 14004 11756
rect 13872 11716 14004 11744
rect 13872 11704 13878 11716
rect 13998 11704 14004 11716
rect 14056 11704 14062 11756
rect 14737 11747 14795 11753
rect 14737 11713 14749 11747
rect 14783 11713 14795 11747
rect 14737 11707 14795 11713
rect 14829 11747 14887 11753
rect 14829 11713 14841 11747
rect 14875 11713 14887 11747
rect 14829 11707 14887 11713
rect 4706 11636 4712 11688
rect 4764 11676 4770 11688
rect 5074 11676 5080 11688
rect 4764 11648 4844 11676
rect 5035 11648 5080 11676
rect 4764 11636 4770 11648
rect 4816 11552 4844 11648
rect 5074 11636 5080 11648
rect 5132 11636 5138 11688
rect 6365 11679 6423 11685
rect 6365 11645 6377 11679
rect 6411 11676 6423 11679
rect 6914 11676 6920 11688
rect 6411 11648 6920 11676
rect 6411 11645 6423 11648
rect 6365 11639 6423 11645
rect 6914 11636 6920 11648
rect 6972 11636 6978 11688
rect 11514 11676 11520 11688
rect 11475 11648 11520 11676
rect 11514 11636 11520 11648
rect 11572 11636 11578 11688
rect 14752 11608 14780 11707
rect 14844 11676 14872 11707
rect 14918 11704 14924 11756
rect 14976 11747 14982 11756
rect 14976 11719 15018 11747
rect 14976 11704 14982 11719
rect 15102 11704 15108 11756
rect 15160 11744 15166 11756
rect 15654 11744 15660 11756
rect 15160 11716 15660 11744
rect 15160 11704 15166 11716
rect 15654 11704 15660 11716
rect 15712 11704 15718 11756
rect 18138 11704 18144 11756
rect 18196 11744 18202 11756
rect 18279 11747 18337 11753
rect 18279 11744 18291 11747
rect 18196 11716 18291 11744
rect 18196 11704 18202 11716
rect 18279 11713 18291 11716
rect 18325 11713 18337 11747
rect 18414 11744 18420 11756
rect 18375 11716 18420 11744
rect 18279 11707 18337 11713
rect 18414 11704 18420 11716
rect 18472 11704 18478 11756
rect 18506 11704 18512 11756
rect 18564 11744 18570 11756
rect 18708 11753 18736 11784
rect 18693 11747 18751 11753
rect 18564 11716 18609 11744
rect 18564 11704 18570 11716
rect 18693 11713 18705 11747
rect 18739 11713 18751 11747
rect 18693 11707 18751 11713
rect 19058 11704 19064 11756
rect 19116 11744 19122 11756
rect 19153 11747 19211 11753
rect 19153 11744 19165 11747
rect 19116 11716 19165 11744
rect 19116 11704 19122 11716
rect 19153 11713 19165 11716
rect 19199 11713 19211 11747
rect 19306 11744 19334 11784
rect 20162 11772 20168 11784
rect 20220 11772 20226 11824
rect 21024 11815 21082 11821
rect 21024 11781 21036 11815
rect 21070 11812 21082 11815
rect 21542 11812 21548 11824
rect 21070 11784 21548 11812
rect 21070 11781 21082 11784
rect 21024 11775 21082 11781
rect 21542 11772 21548 11784
rect 21600 11772 21606 11824
rect 20530 11744 20536 11756
rect 19306 11716 20536 11744
rect 19153 11707 19211 11713
rect 20530 11704 20536 11716
rect 20588 11704 20594 11756
rect 22094 11704 22100 11756
rect 22152 11744 22158 11756
rect 22572 11753 22600 11852
rect 23566 11840 23572 11852
rect 23624 11840 23630 11892
rect 25590 11880 25596 11892
rect 25551 11852 25596 11880
rect 25590 11840 25596 11852
rect 25648 11840 25654 11892
rect 25700 11852 26280 11880
rect 25700 11812 25728 11852
rect 22848 11784 25728 11812
rect 22465 11747 22523 11753
rect 22465 11744 22477 11747
rect 22152 11716 22477 11744
rect 22152 11704 22158 11716
rect 22465 11713 22477 11716
rect 22511 11713 22523 11747
rect 22465 11707 22523 11713
rect 22557 11747 22615 11753
rect 22557 11713 22569 11747
rect 22603 11713 22615 11747
rect 22557 11707 22615 11713
rect 22646 11704 22652 11756
rect 22704 11744 22710 11756
rect 22848 11753 22876 11784
rect 22833 11747 22891 11753
rect 22704 11716 22749 11744
rect 22704 11704 22710 11716
rect 22833 11713 22845 11747
rect 22879 11713 22891 11747
rect 22833 11707 22891 11713
rect 23385 11747 23443 11753
rect 23385 11713 23397 11747
rect 23431 11744 23443 11747
rect 23658 11744 23664 11756
rect 23431 11716 23664 11744
rect 23431 11713 23443 11716
rect 23385 11707 23443 11713
rect 15010 11676 15016 11688
rect 14844 11648 15016 11676
rect 15010 11636 15016 11648
rect 15068 11676 15074 11688
rect 18432 11676 18460 11704
rect 15068 11648 18460 11676
rect 21269 11679 21327 11685
rect 15068 11636 15074 11648
rect 21269 11645 21281 11679
rect 21315 11676 21327 11679
rect 21634 11676 21640 11688
rect 21315 11648 21640 11676
rect 21315 11645 21327 11648
rect 21269 11639 21327 11645
rect 21634 11636 21640 11648
rect 21692 11636 21698 11688
rect 22738 11636 22744 11688
rect 22796 11676 22802 11688
rect 22848 11676 22876 11707
rect 23658 11704 23664 11716
rect 23716 11744 23722 11756
rect 24394 11744 24400 11756
rect 23716 11716 24400 11744
rect 23716 11704 23722 11716
rect 24394 11704 24400 11716
rect 24452 11704 24458 11756
rect 25869 11747 25927 11753
rect 25869 11744 25881 11747
rect 25056 11716 25881 11744
rect 22796 11648 22876 11676
rect 22796 11636 22802 11648
rect 25056 11617 25084 11716
rect 25869 11713 25881 11716
rect 25915 11713 25927 11747
rect 25869 11707 25927 11713
rect 25961 11747 26019 11753
rect 25961 11713 25973 11747
rect 26007 11713 26019 11747
rect 25961 11707 26019 11713
rect 26053 11747 26111 11753
rect 26053 11713 26065 11747
rect 26099 11744 26111 11747
rect 26142 11744 26148 11756
rect 26099 11716 26148 11744
rect 26099 11713 26111 11716
rect 26053 11707 26111 11713
rect 15565 11611 15623 11617
rect 15565 11608 15577 11611
rect 14752 11580 15577 11608
rect 15028 11552 15056 11580
rect 15565 11577 15577 11580
rect 15611 11577 15623 11611
rect 25041 11611 25099 11617
rect 25041 11608 25053 11611
rect 15565 11571 15623 11577
rect 22112 11580 25053 11608
rect 4706 11540 4712 11552
rect 4667 11512 4712 11540
rect 4706 11500 4712 11512
rect 4764 11500 4770 11552
rect 4798 11500 4804 11552
rect 4856 11500 4862 11552
rect 5442 11500 5448 11552
rect 5500 11540 5506 11552
rect 7190 11540 7196 11552
rect 5500 11512 7196 11540
rect 5500 11500 5506 11512
rect 7190 11500 7196 11512
rect 7248 11540 7254 11552
rect 7653 11543 7711 11549
rect 7653 11540 7665 11543
rect 7248 11512 7665 11540
rect 7248 11500 7254 11512
rect 7653 11509 7665 11512
rect 7699 11509 7711 11543
rect 14458 11540 14464 11552
rect 14419 11512 14464 11540
rect 7653 11503 7711 11509
rect 14458 11500 14464 11512
rect 14516 11500 14522 11552
rect 15010 11500 15016 11552
rect 15068 11500 15074 11552
rect 19337 11543 19395 11549
rect 19337 11509 19349 11543
rect 19383 11540 19395 11543
rect 21266 11540 21272 11552
rect 19383 11512 21272 11540
rect 19383 11509 19395 11512
rect 19337 11503 19395 11509
rect 21266 11500 21272 11512
rect 21324 11540 21330 11552
rect 22112 11540 22140 11580
rect 25041 11577 25053 11580
rect 25087 11577 25099 11611
rect 25884 11608 25912 11707
rect 25976 11676 26004 11707
rect 26142 11704 26148 11716
rect 26200 11704 26206 11756
rect 26252 11753 26280 11852
rect 31478 11840 31484 11892
rect 31536 11880 31542 11892
rect 32493 11883 32551 11889
rect 32493 11880 32505 11883
rect 31536 11852 32505 11880
rect 31536 11840 31542 11852
rect 32493 11849 32505 11852
rect 32539 11849 32551 11883
rect 32493 11843 32551 11849
rect 34698 11840 34704 11892
rect 34756 11880 34762 11892
rect 35161 11883 35219 11889
rect 35161 11880 35173 11883
rect 34756 11852 35173 11880
rect 34756 11840 34762 11852
rect 35161 11849 35173 11852
rect 35207 11849 35219 11883
rect 36538 11880 36544 11892
rect 35161 11843 35219 11849
rect 35452 11852 36544 11880
rect 35250 11812 35256 11824
rect 27632 11784 35256 11812
rect 26237 11747 26295 11753
rect 26237 11713 26249 11747
rect 26283 11744 26295 11747
rect 27522 11744 27528 11756
rect 26283 11716 27528 11744
rect 26283 11713 26295 11716
rect 26237 11707 26295 11713
rect 27522 11704 27528 11716
rect 27580 11704 27586 11756
rect 26326 11676 26332 11688
rect 25976 11648 26332 11676
rect 26326 11636 26332 11648
rect 26384 11636 26390 11688
rect 27632 11608 27660 11784
rect 35250 11772 35256 11784
rect 35308 11772 35314 11824
rect 35452 11821 35480 11852
rect 36538 11840 36544 11852
rect 36596 11840 36602 11892
rect 37274 11840 37280 11892
rect 37332 11880 37338 11892
rect 38197 11883 38255 11889
rect 38197 11880 38209 11883
rect 37332 11852 38209 11880
rect 37332 11840 37338 11852
rect 38197 11849 38209 11852
rect 38243 11880 38255 11883
rect 38746 11880 38752 11892
rect 38243 11852 38752 11880
rect 38243 11849 38255 11852
rect 38197 11843 38255 11849
rect 38746 11840 38752 11852
rect 38804 11840 38810 11892
rect 35437 11815 35495 11821
rect 35437 11781 35449 11815
rect 35483 11781 35495 11815
rect 35437 11775 35495 11781
rect 36265 11815 36323 11821
rect 36265 11781 36277 11815
rect 36311 11781 36323 11815
rect 36265 11775 36323 11781
rect 36449 11815 36507 11821
rect 36449 11781 36461 11815
rect 36495 11812 36507 11815
rect 36630 11812 36636 11824
rect 36495 11784 36636 11812
rect 36495 11781 36507 11784
rect 36449 11775 36507 11781
rect 28169 11747 28227 11753
rect 28169 11713 28181 11747
rect 28215 11713 28227 11747
rect 28169 11707 28227 11713
rect 28184 11676 28212 11707
rect 30742 11704 30748 11756
rect 30800 11744 30806 11756
rect 31938 11744 31944 11756
rect 30800 11716 31944 11744
rect 30800 11704 30806 11716
rect 31938 11704 31944 11716
rect 31996 11744 32002 11756
rect 32125 11747 32183 11753
rect 32125 11744 32137 11747
rect 31996 11716 32137 11744
rect 31996 11704 32002 11716
rect 32125 11713 32137 11716
rect 32171 11713 32183 11747
rect 32125 11707 32183 11713
rect 32309 11747 32367 11753
rect 32309 11713 32321 11747
rect 32355 11744 32367 11747
rect 32398 11744 32404 11756
rect 32355 11716 32404 11744
rect 32355 11713 32367 11716
rect 32309 11707 32367 11713
rect 32398 11704 32404 11716
rect 32456 11744 32462 11756
rect 32950 11744 32956 11756
rect 32456 11716 32956 11744
rect 32456 11704 32462 11716
rect 32950 11704 32956 11716
rect 33008 11704 33014 11756
rect 33042 11704 33048 11756
rect 33100 11744 33106 11756
rect 33321 11747 33379 11753
rect 33100 11716 33145 11744
rect 33100 11704 33106 11716
rect 33321 11713 33333 11747
rect 33367 11713 33379 11747
rect 35342 11744 35348 11756
rect 35303 11716 35348 11744
rect 33321 11707 33379 11713
rect 28350 11676 28356 11688
rect 28184 11648 28356 11676
rect 28350 11636 28356 11648
rect 28408 11676 28414 11688
rect 33336 11676 33364 11707
rect 35342 11704 35348 11716
rect 35400 11704 35406 11756
rect 35526 11744 35532 11756
rect 35487 11716 35532 11744
rect 35526 11704 35532 11716
rect 35584 11704 35590 11756
rect 35618 11704 35624 11756
rect 35676 11744 35682 11756
rect 35713 11747 35771 11753
rect 35713 11744 35725 11747
rect 35676 11716 35725 11744
rect 35676 11704 35682 11716
rect 35713 11713 35725 11716
rect 35759 11713 35771 11747
rect 35713 11707 35771 11713
rect 36280 11676 36308 11775
rect 36630 11772 36636 11784
rect 36688 11772 36694 11824
rect 38749 11747 38807 11753
rect 38749 11713 38761 11747
rect 38795 11744 38807 11747
rect 39206 11744 39212 11756
rect 38795 11716 39212 11744
rect 38795 11713 38807 11716
rect 38749 11707 38807 11713
rect 39206 11704 39212 11716
rect 39264 11704 39270 11756
rect 39022 11676 39028 11688
rect 28408 11648 31754 11676
rect 28408 11636 28414 11648
rect 25884 11580 27660 11608
rect 31726 11608 31754 11648
rect 33336 11648 36308 11676
rect 38983 11648 39028 11676
rect 32306 11608 32312 11620
rect 31726 11580 32312 11608
rect 25041 11571 25099 11577
rect 32306 11568 32312 11580
rect 32364 11608 32370 11620
rect 33336 11608 33364 11648
rect 39022 11636 39028 11648
rect 39080 11636 39086 11688
rect 58158 11608 58164 11620
rect 32364 11580 33364 11608
rect 58119 11580 58164 11608
rect 32364 11568 32370 11580
rect 58158 11568 58164 11580
rect 58216 11568 58222 11620
rect 21324 11512 22140 11540
rect 21324 11500 21330 11512
rect 22186 11500 22192 11552
rect 22244 11540 22250 11552
rect 22244 11512 22289 11540
rect 22244 11500 22250 11512
rect 22462 11500 22468 11552
rect 22520 11540 22526 11552
rect 23658 11540 23664 11552
rect 22520 11512 23664 11540
rect 22520 11500 22526 11512
rect 23658 11500 23664 11512
rect 23716 11500 23722 11552
rect 24946 11500 24952 11552
rect 25004 11540 25010 11552
rect 28353 11543 28411 11549
rect 28353 11540 28365 11543
rect 25004 11512 28365 11540
rect 25004 11500 25010 11512
rect 28353 11509 28365 11512
rect 28399 11540 28411 11543
rect 34514 11540 34520 11552
rect 28399 11512 34520 11540
rect 28399 11509 28411 11512
rect 28353 11503 28411 11509
rect 34514 11500 34520 11512
rect 34572 11500 34578 11552
rect 34701 11543 34759 11549
rect 34701 11509 34713 11543
rect 34747 11540 34759 11543
rect 35434 11540 35440 11552
rect 34747 11512 35440 11540
rect 34747 11509 34759 11512
rect 34701 11503 34759 11509
rect 35434 11500 35440 11512
rect 35492 11500 35498 11552
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 3786 11336 3792 11348
rect 3747 11308 3792 11336
rect 3786 11296 3792 11308
rect 3844 11296 3850 11348
rect 6914 11336 6920 11348
rect 6564 11308 6920 11336
rect 3237 11203 3295 11209
rect 3237 11169 3249 11203
rect 3283 11200 3295 11203
rect 3878 11200 3884 11212
rect 3283 11172 3884 11200
rect 3283 11169 3295 11172
rect 3237 11163 3295 11169
rect 3878 11160 3884 11172
rect 3936 11160 3942 11212
rect 5258 11160 5264 11212
rect 5316 11200 5322 11212
rect 5629 11203 5687 11209
rect 5629 11200 5641 11203
rect 5316 11172 5641 11200
rect 5316 11160 5322 11172
rect 5629 11169 5641 11172
rect 5675 11169 5687 11203
rect 5629 11163 5687 11169
rect 5721 11203 5779 11209
rect 5721 11169 5733 11203
rect 5767 11200 5779 11203
rect 6564 11200 6592 11308
rect 6914 11296 6920 11308
rect 6972 11296 6978 11348
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 12492 11308 12537 11336
rect 12492 11296 12498 11308
rect 13354 11296 13360 11348
rect 13412 11336 13418 11348
rect 14185 11339 14243 11345
rect 14185 11336 14197 11339
rect 13412 11308 14197 11336
rect 13412 11296 13418 11308
rect 14185 11305 14197 11308
rect 14231 11305 14243 11339
rect 14185 11299 14243 11305
rect 18138 11296 18144 11348
rect 18196 11336 18202 11348
rect 18506 11336 18512 11348
rect 18196 11308 18512 11336
rect 18196 11296 18202 11308
rect 18506 11296 18512 11308
rect 18564 11296 18570 11348
rect 21085 11339 21143 11345
rect 21085 11305 21097 11339
rect 21131 11336 21143 11339
rect 21174 11336 21180 11348
rect 21131 11308 21180 11336
rect 21131 11305 21143 11308
rect 21085 11299 21143 11305
rect 21174 11296 21180 11308
rect 21232 11296 21238 11348
rect 22738 11336 22744 11348
rect 21376 11308 22744 11336
rect 6638 11228 6644 11280
rect 6696 11268 6702 11280
rect 6696 11240 7972 11268
rect 6696 11228 6702 11240
rect 6730 11200 6736 11212
rect 5767 11172 6592 11200
rect 6691 11172 6736 11200
rect 5767 11169 5779 11172
rect 5721 11163 5779 11169
rect 6730 11160 6736 11172
rect 6788 11160 6794 11212
rect 6831 11203 6889 11209
rect 6831 11169 6843 11203
rect 6877 11200 6889 11203
rect 7190 11200 7196 11212
rect 6877 11172 7196 11200
rect 6877 11169 6889 11172
rect 6831 11163 6889 11169
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 7282 11160 7288 11212
rect 7340 11200 7346 11212
rect 7837 11203 7895 11209
rect 7837 11200 7849 11203
rect 7340 11172 7849 11200
rect 7340 11160 7346 11172
rect 7837 11169 7849 11172
rect 7883 11169 7895 11203
rect 7837 11163 7895 11169
rect 2682 11092 2688 11144
rect 2740 11132 2746 11144
rect 2961 11135 3019 11141
rect 2961 11132 2973 11135
rect 2740 11104 2973 11132
rect 2740 11092 2746 11104
rect 2961 11101 2973 11104
rect 3007 11101 3019 11135
rect 2961 11095 3019 11101
rect 3973 11135 4031 11141
rect 3973 11101 3985 11135
rect 4019 11132 4031 11135
rect 4706 11132 4712 11144
rect 4019 11104 4712 11132
rect 4019 11101 4031 11104
rect 3973 11095 4031 11101
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 4890 11092 4896 11144
rect 4948 11132 4954 11144
rect 6549 11135 6607 11141
rect 6549 11132 6561 11135
rect 4948 11104 6561 11132
rect 4948 11092 4954 11104
rect 6549 11101 6561 11104
rect 6595 11101 6607 11135
rect 6549 11095 6607 11101
rect 6913 11133 6971 11139
rect 6913 11099 6925 11133
rect 6959 11132 6971 11133
rect 7101 11135 7159 11141
rect 6959 11104 7052 11132
rect 6959 11099 6971 11104
rect 6913 11093 6971 11099
rect 5261 11067 5319 11073
rect 5261 11033 5273 11067
rect 5307 11064 5319 11067
rect 5626 11064 5632 11076
rect 5307 11036 5632 11064
rect 5307 11033 5319 11036
rect 5261 11027 5319 11033
rect 5626 11024 5632 11036
rect 5684 11024 5690 11076
rect 5905 11067 5963 11073
rect 5905 11033 5917 11067
rect 5951 11064 5963 11067
rect 5951 11036 6776 11064
rect 5951 11033 5963 11036
rect 5905 11027 5963 11033
rect 4706 10956 4712 11008
rect 4764 10996 4770 11008
rect 4982 10996 4988 11008
rect 4764 10968 4988 10996
rect 4764 10956 4770 10968
rect 4982 10956 4988 10968
rect 5040 10956 5046 11008
rect 6362 10996 6368 11008
rect 6323 10968 6368 10996
rect 6362 10956 6368 10968
rect 6420 10956 6426 11008
rect 6748 10996 6776 11036
rect 7024 10996 7052 11104
rect 7101 11101 7113 11135
rect 7147 11132 7159 11135
rect 7466 11132 7472 11144
rect 7147 11104 7472 11132
rect 7147 11101 7159 11104
rect 7101 11095 7159 11101
rect 7466 11092 7472 11104
rect 7524 11092 7530 11144
rect 7561 11135 7619 11141
rect 7561 11101 7573 11135
rect 7607 11132 7619 11135
rect 7944 11132 7972 11240
rect 15930 11228 15936 11280
rect 15988 11268 15994 11280
rect 16025 11271 16083 11277
rect 16025 11268 16037 11271
rect 15988 11240 16037 11268
rect 15988 11228 15994 11240
rect 16025 11237 16037 11240
rect 16071 11237 16083 11271
rect 16025 11231 16083 11237
rect 17037 11271 17095 11277
rect 17037 11237 17049 11271
rect 17083 11268 17095 11271
rect 17218 11268 17224 11280
rect 17083 11240 17224 11268
rect 17083 11237 17095 11240
rect 17037 11231 17095 11237
rect 17218 11228 17224 11240
rect 17276 11268 17282 11280
rect 21266 11268 21272 11280
rect 17276 11240 21272 11268
rect 17276 11228 17282 11240
rect 21266 11228 21272 11240
rect 21324 11228 21330 11280
rect 15654 11160 15660 11212
rect 15712 11200 15718 11212
rect 21376 11200 21404 11308
rect 22738 11296 22744 11308
rect 22796 11296 22802 11348
rect 26142 11336 26148 11348
rect 26103 11308 26148 11336
rect 26142 11296 26148 11308
rect 26200 11296 26206 11348
rect 29917 11339 29975 11345
rect 29917 11305 29929 11339
rect 29963 11336 29975 11339
rect 30190 11336 30196 11348
rect 29963 11308 30196 11336
rect 29963 11305 29975 11308
rect 29917 11299 29975 11305
rect 30190 11296 30196 11308
rect 30248 11336 30254 11348
rect 30374 11336 30380 11348
rect 30248 11308 30380 11336
rect 30248 11296 30254 11308
rect 30374 11296 30380 11308
rect 30432 11296 30438 11348
rect 32953 11339 33011 11345
rect 32953 11336 32965 11339
rect 31726 11308 32965 11336
rect 24486 11228 24492 11280
rect 24544 11268 24550 11280
rect 31726 11268 31754 11308
rect 32953 11305 32965 11308
rect 32999 11336 33011 11339
rect 33042 11336 33048 11348
rect 32999 11308 33048 11336
rect 32999 11305 33011 11308
rect 32953 11299 33011 11305
rect 33042 11296 33048 11308
rect 33100 11296 33106 11348
rect 34514 11296 34520 11348
rect 34572 11336 34578 11348
rect 34701 11339 34759 11345
rect 34701 11336 34713 11339
rect 34572 11308 34713 11336
rect 34572 11296 34578 11308
rect 34701 11305 34713 11308
rect 34747 11305 34759 11339
rect 34701 11299 34759 11305
rect 24544 11240 31754 11268
rect 24544 11228 24550 11240
rect 21634 11200 21640 11212
rect 15712 11172 21404 11200
rect 21595 11172 21640 11200
rect 15712 11160 15718 11172
rect 21634 11160 21640 11172
rect 21692 11160 21698 11212
rect 23566 11200 23572 11212
rect 23479 11172 23572 11200
rect 23566 11160 23572 11172
rect 23624 11200 23630 11212
rect 24578 11200 24584 11212
rect 23624 11172 24584 11200
rect 23624 11160 23630 11172
rect 24578 11160 24584 11172
rect 24636 11200 24642 11212
rect 26326 11200 26332 11212
rect 24636 11172 26332 11200
rect 24636 11160 24642 11172
rect 26326 11160 26332 11172
rect 26384 11200 26390 11212
rect 28169 11203 28227 11209
rect 28169 11200 28181 11203
rect 26384 11172 28181 11200
rect 26384 11160 26390 11172
rect 28169 11169 28181 11172
rect 28215 11169 28227 11203
rect 28169 11163 28227 11169
rect 28445 11203 28503 11209
rect 28445 11169 28457 11203
rect 28491 11200 28503 11203
rect 29086 11200 29092 11212
rect 28491 11172 29092 11200
rect 28491 11169 28503 11172
rect 28445 11163 28503 11169
rect 29086 11160 29092 11172
rect 29144 11200 29150 11212
rect 31846 11200 31852 11212
rect 29144 11172 31852 11200
rect 29144 11160 29150 11172
rect 9122 11132 9128 11144
rect 7607 11104 7972 11132
rect 9083 11104 9128 11132
rect 7607 11101 7619 11104
rect 7561 11095 7619 11101
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 11514 11132 11520 11144
rect 11475 11104 11520 11132
rect 11514 11092 11520 11104
rect 11572 11132 11578 11144
rect 12253 11135 12311 11141
rect 12253 11132 12265 11135
rect 11572 11104 12265 11132
rect 11572 11092 11578 11104
rect 12253 11101 12265 11104
rect 12299 11101 12311 11135
rect 12253 11095 12311 11101
rect 14458 11092 14464 11144
rect 14516 11132 14522 11144
rect 15298 11135 15356 11141
rect 15298 11132 15310 11135
rect 14516 11104 15310 11132
rect 14516 11092 14522 11104
rect 15298 11101 15310 11104
rect 15344 11101 15356 11135
rect 15298 11095 15356 11101
rect 15470 11092 15476 11144
rect 15528 11132 15534 11144
rect 15565 11135 15623 11141
rect 15565 11132 15577 11135
rect 15528 11104 15577 11132
rect 15528 11092 15534 11104
rect 15565 11101 15577 11104
rect 15611 11101 15623 11135
rect 21652 11132 21680 11160
rect 21652 11104 23428 11132
rect 15565 11095 15623 11101
rect 14826 11024 14832 11076
rect 14884 11064 14890 11076
rect 16209 11067 16267 11073
rect 16209 11064 16221 11067
rect 14884 11036 16221 11064
rect 14884 11024 14890 11036
rect 16209 11033 16221 11036
rect 16255 11064 16267 11067
rect 16853 11067 16911 11073
rect 16853 11064 16865 11067
rect 16255 11036 16865 11064
rect 16255 11033 16267 11036
rect 16209 11027 16267 11033
rect 16853 11033 16865 11036
rect 16899 11033 16911 11067
rect 17770 11064 17776 11076
rect 17731 11036 17776 11064
rect 16853 11027 16911 11033
rect 17770 11024 17776 11036
rect 17828 11064 17834 11076
rect 18417 11067 18475 11073
rect 18417 11064 18429 11067
rect 17828 11036 18429 11064
rect 17828 11024 17834 11036
rect 18417 11033 18429 11036
rect 18463 11033 18475 11067
rect 18417 11027 18475 11033
rect 18506 11024 18512 11076
rect 18564 11064 18570 11076
rect 19334 11064 19340 11076
rect 18564 11036 19340 11064
rect 18564 11024 18570 11036
rect 19334 11024 19340 11036
rect 19392 11024 19398 11076
rect 20441 11067 20499 11073
rect 20441 11033 20453 11067
rect 20487 11064 20499 11067
rect 20806 11064 20812 11076
rect 20487 11036 20812 11064
rect 20487 11033 20499 11036
rect 20441 11027 20499 11033
rect 20806 11024 20812 11036
rect 20864 11064 20870 11076
rect 20993 11067 21051 11073
rect 20993 11064 21005 11067
rect 20864 11036 21005 11064
rect 20864 11024 20870 11036
rect 20993 11033 21005 11036
rect 21039 11064 21051 11067
rect 21450 11064 21456 11076
rect 21039 11036 21456 11064
rect 21039 11033 21051 11036
rect 20993 11027 21051 11033
rect 21450 11024 21456 11036
rect 21508 11024 21514 11076
rect 21904 11067 21962 11073
rect 21904 11033 21916 11067
rect 21950 11064 21962 11067
rect 22186 11064 22192 11076
rect 21950 11036 22192 11064
rect 21950 11033 21962 11036
rect 21904 11027 21962 11033
rect 22186 11024 22192 11036
rect 22244 11024 22250 11076
rect 23400 11064 23428 11104
rect 23474 11092 23480 11144
rect 23532 11132 23538 11144
rect 23658 11132 23664 11144
rect 23532 11104 23577 11132
rect 23619 11104 23664 11132
rect 23532 11092 23538 11104
rect 23658 11092 23664 11104
rect 23716 11092 23722 11144
rect 25958 11132 25964 11144
rect 25919 11104 25964 11132
rect 25958 11092 25964 11104
rect 26016 11092 26022 11144
rect 30190 11092 30196 11144
rect 30248 11132 30254 11144
rect 30760 11141 30788 11172
rect 31846 11160 31852 11172
rect 31904 11160 31910 11212
rect 30653 11135 30711 11141
rect 30653 11132 30665 11135
rect 30248 11104 30665 11132
rect 30248 11092 30254 11104
rect 30653 11101 30665 11104
rect 30699 11101 30711 11135
rect 30653 11095 30711 11101
rect 30745 11135 30803 11141
rect 30745 11101 30757 11135
rect 30791 11101 30803 11135
rect 30745 11095 30803 11101
rect 30834 11092 30840 11144
rect 30892 11132 30898 11144
rect 31021 11135 31079 11141
rect 30892 11104 30937 11132
rect 30892 11092 30898 11104
rect 31021 11101 31033 11135
rect 31067 11132 31079 11135
rect 31294 11132 31300 11144
rect 31067 11104 31300 11132
rect 31067 11101 31079 11104
rect 31021 11095 31079 11101
rect 25038 11064 25044 11076
rect 23400 11036 25044 11064
rect 25038 11024 25044 11036
rect 25096 11024 25102 11076
rect 25774 11064 25780 11076
rect 25735 11036 25780 11064
rect 25774 11024 25780 11036
rect 25832 11024 25838 11076
rect 30377 11067 30435 11073
rect 30377 11033 30389 11067
rect 30423 11064 30435 11067
rect 30466 11064 30472 11076
rect 30423 11036 30472 11064
rect 30423 11033 30435 11036
rect 30377 11027 30435 11033
rect 30466 11024 30472 11036
rect 30524 11024 30530 11076
rect 30558 11024 30564 11076
rect 30616 11064 30622 11076
rect 31036 11064 31064 11095
rect 31294 11092 31300 11104
rect 31352 11132 31358 11144
rect 32030 11132 32036 11144
rect 31352 11104 32036 11132
rect 31352 11092 31358 11104
rect 32030 11092 32036 11104
rect 32088 11092 32094 11144
rect 32306 11132 32312 11144
rect 32267 11104 32312 11132
rect 32306 11092 32312 11104
rect 32364 11092 32370 11144
rect 30616 11036 31064 11064
rect 34716 11064 34744 11299
rect 39022 11268 39028 11280
rect 35636 11240 39028 11268
rect 35434 11160 35440 11212
rect 35492 11160 35498 11212
rect 35250 11092 35256 11144
rect 35308 11132 35314 11144
rect 35452 11132 35480 11160
rect 35636 11141 35664 11240
rect 36357 11203 36415 11209
rect 36357 11200 36369 11203
rect 35728 11172 36369 11200
rect 35728 11141 35756 11172
rect 36357 11169 36369 11172
rect 36403 11169 36415 11203
rect 36357 11163 36415 11169
rect 38197 11203 38255 11209
rect 38197 11169 38209 11203
rect 38243 11200 38255 11203
rect 38243 11172 38884 11200
rect 38243 11169 38255 11172
rect 38197 11163 38255 11169
rect 35529 11135 35587 11141
rect 35529 11132 35541 11135
rect 35308 11104 35541 11132
rect 35308 11092 35314 11104
rect 35529 11101 35541 11104
rect 35575 11101 35587 11135
rect 35529 11095 35587 11101
rect 35621 11135 35679 11141
rect 35621 11101 35633 11135
rect 35667 11101 35679 11135
rect 35621 11095 35679 11101
rect 35713 11135 35771 11141
rect 35713 11101 35725 11135
rect 35759 11101 35771 11135
rect 35713 11095 35771 11101
rect 35897 11135 35955 11141
rect 35897 11101 35909 11135
rect 35943 11101 35955 11135
rect 36538 11132 36544 11144
rect 36499 11104 36544 11132
rect 35897 11095 35955 11101
rect 35912 11064 35940 11095
rect 36538 11092 36544 11104
rect 36596 11092 36602 11144
rect 36630 11092 36636 11144
rect 36688 11132 36694 11144
rect 38856 11141 38884 11172
rect 38948 11141 38976 11240
rect 39022 11228 39028 11240
rect 39080 11228 39086 11280
rect 38657 11135 38715 11141
rect 38657 11132 38669 11135
rect 36688 11104 38669 11132
rect 36688 11092 36694 11104
rect 38657 11101 38669 11104
rect 38703 11101 38715 11135
rect 38657 11095 38715 11101
rect 38841 11135 38899 11141
rect 38841 11101 38853 11135
rect 38887 11101 38899 11135
rect 38841 11095 38899 11101
rect 38933 11135 38991 11141
rect 38933 11101 38945 11135
rect 38979 11101 38991 11135
rect 38933 11095 38991 11101
rect 39025 11135 39083 11141
rect 39025 11101 39037 11135
rect 39071 11101 39083 11135
rect 39853 11135 39911 11141
rect 39853 11132 39865 11135
rect 39025 11095 39083 11101
rect 39132 11104 39865 11132
rect 34716 11036 35940 11064
rect 36725 11067 36783 11073
rect 30616 11024 30622 11036
rect 36725 11033 36737 11067
rect 36771 11064 36783 11067
rect 37550 11064 37556 11076
rect 36771 11036 37556 11064
rect 36771 11033 36783 11036
rect 36725 11027 36783 11033
rect 37550 11024 37556 11036
rect 37608 11064 37614 11076
rect 37829 11067 37887 11073
rect 37829 11064 37841 11067
rect 37608 11036 37841 11064
rect 37608 11024 37614 11036
rect 37829 11033 37841 11036
rect 37875 11033 37887 11067
rect 38010 11064 38016 11076
rect 37971 11036 38016 11064
rect 37829 11027 37887 11033
rect 38010 11024 38016 11036
rect 38068 11024 38074 11076
rect 8938 10996 8944 11008
rect 6748 10968 7052 10996
rect 8899 10968 8944 10996
rect 8938 10956 8944 10968
rect 8996 10956 9002 11008
rect 11701 10999 11759 11005
rect 11701 10965 11713 10999
rect 11747 10996 11759 10999
rect 14182 10996 14188 11008
rect 11747 10968 14188 10996
rect 11747 10965 11759 10968
rect 11701 10959 11759 10965
rect 14182 10956 14188 10968
rect 14240 10996 14246 11008
rect 18230 10996 18236 11008
rect 14240 10968 18236 10996
rect 14240 10956 14246 10968
rect 18230 10956 18236 10968
rect 18288 10956 18294 11008
rect 19242 10956 19248 11008
rect 19300 10996 19306 11008
rect 19705 10999 19763 11005
rect 19705 10996 19717 10999
rect 19300 10968 19717 10996
rect 19300 10956 19306 10968
rect 19705 10965 19717 10968
rect 19751 10996 19763 10999
rect 20070 10996 20076 11008
rect 19751 10968 20076 10996
rect 19751 10965 19763 10968
rect 19705 10959 19763 10965
rect 20070 10956 20076 10968
rect 20128 10956 20134 11008
rect 23014 10996 23020 11008
rect 22975 10968 23020 10996
rect 23014 10956 23020 10968
rect 23072 10956 23078 11008
rect 35253 10999 35311 11005
rect 35253 10965 35265 10999
rect 35299 10996 35311 10999
rect 35342 10996 35348 11008
rect 35299 10968 35348 10996
rect 35299 10965 35311 10968
rect 35253 10959 35311 10965
rect 35342 10956 35348 10968
rect 35400 10956 35406 11008
rect 38672 10996 38700 11095
rect 38746 11024 38752 11076
rect 38804 11064 38810 11076
rect 39040 11064 39068 11095
rect 38804 11036 39068 11064
rect 38804 11024 38810 11036
rect 39132 10996 39160 11104
rect 39853 11101 39865 11104
rect 39899 11101 39911 11135
rect 39853 11095 39911 11101
rect 39301 11067 39359 11073
rect 39301 11033 39313 11067
rect 39347 11064 39359 11067
rect 40126 11064 40132 11076
rect 39347 11036 40132 11064
rect 39347 11033 39359 11036
rect 39301 11027 39359 11033
rect 40126 11024 40132 11036
rect 40184 11024 40190 11076
rect 38672 10968 39160 10996
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 4341 10795 4399 10801
rect 4341 10761 4353 10795
rect 4387 10792 4399 10795
rect 5350 10792 5356 10804
rect 4387 10764 5356 10792
rect 4387 10761 4399 10764
rect 4341 10755 4399 10761
rect 5350 10752 5356 10764
rect 5408 10752 5414 10804
rect 7009 10795 7067 10801
rect 7009 10761 7021 10795
rect 7055 10792 7067 10795
rect 7466 10792 7472 10804
rect 7055 10764 7472 10792
rect 7055 10761 7067 10764
rect 7009 10755 7067 10761
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 7837 10795 7895 10801
rect 7837 10761 7849 10795
rect 7883 10792 7895 10795
rect 9122 10792 9128 10804
rect 7883 10764 9128 10792
rect 7883 10761 7895 10764
rect 7837 10755 7895 10761
rect 9122 10752 9128 10764
rect 9180 10752 9186 10804
rect 13998 10792 14004 10804
rect 13959 10764 14004 10792
rect 13998 10752 14004 10764
rect 14056 10752 14062 10804
rect 22646 10752 22652 10804
rect 22704 10792 22710 10804
rect 22741 10795 22799 10801
rect 22741 10792 22753 10795
rect 22704 10764 22753 10792
rect 22704 10752 22710 10764
rect 22741 10761 22753 10764
rect 22787 10761 22799 10795
rect 22741 10755 22799 10761
rect 23198 10752 23204 10804
rect 23256 10792 23262 10804
rect 27154 10792 27160 10804
rect 23256 10764 27160 10792
rect 23256 10752 23262 10764
rect 27154 10752 27160 10764
rect 27212 10752 27218 10804
rect 28261 10795 28319 10801
rect 28261 10761 28273 10795
rect 28307 10792 28319 10795
rect 28307 10764 30696 10792
rect 28307 10761 28319 10764
rect 28261 10755 28319 10761
rect 4614 10684 4620 10736
rect 4672 10724 4678 10736
rect 5258 10724 5264 10736
rect 4672 10696 5264 10724
rect 4672 10684 4678 10696
rect 5258 10684 5264 10696
rect 5316 10684 5322 10736
rect 8564 10727 8622 10733
rect 8564 10693 8576 10727
rect 8610 10724 8622 10727
rect 8938 10724 8944 10736
rect 8610 10696 8944 10724
rect 8610 10693 8622 10696
rect 8564 10687 8622 10693
rect 8938 10684 8944 10696
rect 8996 10684 9002 10736
rect 14366 10684 14372 10736
rect 14424 10724 14430 10736
rect 15114 10727 15172 10733
rect 15114 10724 15126 10727
rect 14424 10696 15126 10724
rect 14424 10684 14430 10696
rect 15114 10693 15126 10696
rect 15160 10693 15172 10727
rect 15114 10687 15172 10693
rect 22557 10727 22615 10733
rect 22557 10693 22569 10727
rect 22603 10724 22615 10727
rect 23014 10724 23020 10736
rect 22603 10696 23020 10724
rect 22603 10693 22615 10696
rect 22557 10687 22615 10693
rect 23014 10684 23020 10696
rect 23072 10684 23078 10736
rect 24412 10696 25820 10724
rect 2038 10616 2044 10668
rect 2096 10656 2102 10668
rect 2225 10659 2283 10665
rect 2225 10656 2237 10659
rect 2096 10628 2237 10656
rect 2096 10616 2102 10628
rect 2225 10625 2237 10628
rect 2271 10625 2283 10659
rect 2225 10619 2283 10625
rect 4433 10659 4491 10665
rect 4433 10625 4445 10659
rect 4479 10656 4491 10659
rect 4982 10656 4988 10668
rect 4479 10628 4988 10656
rect 4479 10625 4491 10628
rect 4433 10619 4491 10625
rect 4982 10616 4988 10628
rect 5040 10616 5046 10668
rect 7650 10656 7656 10668
rect 7611 10628 7656 10656
rect 7650 10616 7656 10628
rect 7708 10616 7714 10668
rect 7926 10616 7932 10668
rect 7984 10656 7990 10668
rect 8297 10659 8355 10665
rect 8297 10656 8309 10659
rect 7984 10628 8309 10656
rect 7984 10616 7990 10628
rect 8297 10625 8309 10628
rect 8343 10625 8355 10659
rect 12618 10656 12624 10668
rect 8297 10619 8355 10625
rect 8404 10628 12624 10656
rect 2682 10548 2688 10600
rect 2740 10588 2746 10600
rect 7469 10591 7527 10597
rect 7469 10588 7481 10591
rect 2740 10560 7481 10588
rect 2740 10548 2746 10560
rect 7469 10557 7481 10560
rect 7515 10588 7527 10591
rect 8404 10588 8432 10628
rect 12618 10616 12624 10628
rect 12676 10616 12682 10668
rect 22186 10616 22192 10668
rect 22244 10656 22250 10668
rect 22373 10659 22431 10665
rect 22373 10656 22385 10659
rect 22244 10628 22385 10656
rect 22244 10616 22250 10628
rect 22373 10625 22385 10628
rect 22419 10656 22431 10659
rect 24412 10656 24440 10696
rect 25792 10668 25820 10696
rect 28810 10684 28816 10736
rect 28868 10724 28874 10736
rect 30668 10733 30696 10764
rect 30834 10752 30840 10804
rect 30892 10792 30898 10804
rect 31021 10795 31079 10801
rect 31021 10792 31033 10795
rect 30892 10764 31033 10792
rect 30892 10752 30898 10764
rect 31021 10761 31033 10764
rect 31067 10761 31079 10795
rect 31021 10755 31079 10761
rect 36449 10795 36507 10801
rect 36449 10761 36461 10795
rect 36495 10792 36507 10795
rect 36538 10792 36544 10804
rect 36495 10764 36544 10792
rect 36495 10761 36507 10764
rect 36449 10755 36507 10761
rect 36538 10752 36544 10764
rect 36596 10752 36602 10804
rect 38010 10752 38016 10804
rect 38068 10792 38074 10804
rect 41233 10795 41291 10801
rect 41233 10792 41245 10795
rect 38068 10764 41245 10792
rect 38068 10752 38074 10764
rect 41233 10761 41245 10764
rect 41279 10761 41291 10795
rect 41233 10755 41291 10761
rect 29825 10727 29883 10733
rect 29825 10724 29837 10727
rect 28868 10696 29837 10724
rect 28868 10684 28874 10696
rect 24578 10656 24584 10668
rect 22419 10628 24440 10656
rect 24539 10628 24584 10656
rect 22419 10625 22431 10628
rect 22373 10619 22431 10625
rect 24578 10616 24584 10628
rect 24636 10616 24642 10668
rect 25038 10656 25044 10668
rect 24999 10628 25044 10656
rect 25038 10616 25044 10628
rect 25096 10616 25102 10668
rect 25314 10665 25320 10668
rect 25308 10619 25320 10665
rect 25372 10656 25378 10668
rect 25372 10628 25408 10656
rect 25314 10616 25320 10619
rect 25372 10616 25378 10628
rect 25774 10616 25780 10668
rect 25832 10656 25838 10668
rect 29012 10665 29040 10696
rect 29825 10693 29837 10696
rect 29871 10693 29883 10727
rect 29825 10687 29883 10693
rect 30653 10727 30711 10733
rect 30653 10693 30665 10727
rect 30699 10724 30711 10727
rect 30742 10724 30748 10736
rect 30699 10696 30748 10724
rect 30699 10693 30711 10696
rect 30653 10687 30711 10693
rect 30742 10684 30748 10696
rect 30800 10684 30806 10736
rect 37645 10727 37703 10733
rect 37645 10693 37657 10727
rect 37691 10724 37703 10727
rect 37918 10724 37924 10736
rect 37691 10696 37924 10724
rect 37691 10693 37703 10696
rect 37645 10687 37703 10693
rect 37918 10684 37924 10696
rect 37976 10684 37982 10736
rect 40126 10733 40132 10736
rect 40120 10724 40132 10733
rect 40087 10696 40132 10724
rect 40120 10687 40132 10696
rect 40126 10684 40132 10687
rect 40184 10684 40190 10736
rect 28077 10659 28135 10665
rect 28077 10656 28089 10659
rect 25832 10628 28089 10656
rect 25832 10616 25838 10628
rect 28077 10625 28089 10628
rect 28123 10625 28135 10659
rect 28077 10619 28135 10625
rect 28997 10659 29055 10665
rect 28997 10625 29009 10659
rect 29043 10625 29055 10659
rect 28997 10619 29055 10625
rect 29102 10662 29160 10668
rect 29102 10628 29114 10662
rect 29148 10628 29160 10662
rect 29102 10622 29160 10628
rect 29202 10659 29260 10665
rect 29202 10625 29214 10659
rect 29248 10656 29260 10659
rect 29365 10659 29423 10665
rect 29248 10628 29316 10656
rect 29248 10625 29260 10628
rect 15378 10588 15384 10600
rect 7515 10560 8432 10588
rect 15339 10560 15384 10588
rect 7515 10557 7527 10560
rect 7469 10551 7527 10557
rect 15378 10548 15384 10560
rect 15436 10548 15442 10600
rect 24302 10588 24308 10600
rect 24263 10560 24308 10588
rect 24302 10548 24308 10560
rect 24360 10548 24366 10600
rect 29104 10532 29132 10622
rect 29202 10619 29260 10625
rect 15470 10480 15476 10532
rect 15528 10520 15534 10532
rect 22830 10520 22836 10532
rect 15528 10492 22836 10520
rect 15528 10480 15534 10492
rect 22830 10480 22836 10492
rect 22888 10480 22894 10532
rect 29086 10480 29092 10532
rect 29144 10480 29150 10532
rect 29288 10520 29316 10628
rect 29365 10625 29377 10659
rect 29411 10656 29423 10659
rect 30558 10656 30564 10668
rect 29411 10628 30564 10656
rect 29411 10625 29423 10628
rect 29365 10619 29423 10625
rect 30558 10616 30564 10628
rect 30616 10616 30622 10668
rect 30834 10656 30840 10668
rect 30795 10628 30840 10656
rect 30834 10616 30840 10628
rect 30892 10616 30898 10668
rect 34790 10616 34796 10668
rect 34848 10656 34854 10668
rect 35342 10665 35348 10668
rect 35069 10659 35127 10665
rect 35069 10656 35081 10659
rect 34848 10628 35081 10656
rect 34848 10616 34854 10628
rect 35069 10625 35081 10628
rect 35115 10625 35127 10659
rect 35336 10656 35348 10665
rect 35303 10628 35348 10656
rect 35069 10619 35127 10625
rect 35336 10619 35348 10628
rect 35342 10616 35348 10619
rect 35400 10616 35406 10668
rect 39853 10591 39911 10597
rect 39853 10588 39865 10591
rect 38948 10560 39865 10588
rect 29362 10520 29368 10532
rect 29288 10492 29368 10520
rect 29362 10480 29368 10492
rect 29420 10480 29426 10532
rect 38948 10464 38976 10560
rect 39853 10557 39865 10560
rect 39899 10557 39911 10591
rect 39853 10551 39911 10557
rect 2406 10452 2412 10464
rect 2367 10424 2412 10452
rect 2406 10412 2412 10424
rect 2464 10412 2470 10464
rect 9677 10455 9735 10461
rect 9677 10421 9689 10455
rect 9723 10452 9735 10455
rect 9766 10452 9772 10464
rect 9723 10424 9772 10452
rect 9723 10421 9735 10424
rect 9677 10415 9735 10421
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 10226 10452 10232 10464
rect 10187 10424 10232 10452
rect 10226 10412 10232 10424
rect 10284 10412 10290 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12492 10424 12537 10452
rect 12492 10412 12498 10424
rect 12802 10412 12808 10464
rect 12860 10452 12866 10464
rect 12989 10455 13047 10461
rect 12989 10452 13001 10455
rect 12860 10424 13001 10452
rect 12860 10412 12866 10424
rect 12989 10421 13001 10424
rect 13035 10452 13047 10455
rect 16574 10452 16580 10464
rect 13035 10424 16580 10452
rect 13035 10421 13047 10424
rect 12989 10415 13047 10421
rect 16574 10412 16580 10424
rect 16632 10412 16638 10464
rect 18414 10412 18420 10464
rect 18472 10452 18478 10464
rect 18969 10455 19027 10461
rect 18969 10452 18981 10455
rect 18472 10424 18981 10452
rect 18472 10412 18478 10424
rect 18969 10421 18981 10424
rect 19015 10452 19027 10455
rect 19058 10452 19064 10464
rect 19015 10424 19064 10452
rect 19015 10421 19027 10424
rect 18969 10415 19027 10421
rect 19058 10412 19064 10424
rect 19116 10412 19122 10464
rect 19334 10412 19340 10464
rect 19392 10452 19398 10464
rect 19610 10452 19616 10464
rect 19392 10424 19616 10452
rect 19392 10412 19398 10424
rect 19610 10412 19616 10424
rect 19668 10412 19674 10464
rect 26326 10412 26332 10464
rect 26384 10452 26390 10464
rect 26421 10455 26479 10461
rect 26421 10452 26433 10455
rect 26384 10424 26433 10452
rect 26384 10412 26390 10424
rect 26421 10421 26433 10424
rect 26467 10421 26479 10455
rect 26421 10415 26479 10421
rect 28534 10412 28540 10464
rect 28592 10452 28598 10464
rect 28721 10455 28779 10461
rect 28721 10452 28733 10455
rect 28592 10424 28733 10452
rect 28592 10412 28598 10424
rect 28721 10421 28733 10424
rect 28767 10421 28779 10455
rect 38930 10452 38936 10464
rect 38891 10424 38936 10452
rect 28721 10415 28779 10421
rect 38930 10412 38936 10424
rect 38988 10412 38994 10464
rect 58158 10452 58164 10464
rect 58119 10424 58164 10452
rect 58158 10412 58164 10424
rect 58216 10412 58222 10464
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 2038 10248 2044 10260
rect 1999 10220 2044 10248
rect 2038 10208 2044 10220
rect 2096 10208 2102 10260
rect 5074 10208 5080 10260
rect 5132 10248 5138 10260
rect 5442 10248 5448 10260
rect 5132 10220 5448 10248
rect 5132 10208 5138 10220
rect 5442 10208 5448 10220
rect 5500 10248 5506 10260
rect 7006 10248 7012 10260
rect 5500 10220 7012 10248
rect 5500 10208 5506 10220
rect 7006 10208 7012 10220
rect 7064 10208 7070 10260
rect 7650 10208 7656 10260
rect 7708 10248 7714 10260
rect 8941 10251 8999 10257
rect 8941 10248 8953 10251
rect 7708 10220 8953 10248
rect 7708 10208 7714 10220
rect 8941 10217 8953 10220
rect 8987 10217 8999 10251
rect 21266 10248 21272 10260
rect 21227 10220 21272 10248
rect 8941 10211 8999 10217
rect 21266 10208 21272 10220
rect 21324 10208 21330 10260
rect 22186 10248 22192 10260
rect 22147 10220 22192 10248
rect 22186 10208 22192 10220
rect 22244 10208 22250 10260
rect 25314 10208 25320 10260
rect 25372 10248 25378 10260
rect 25409 10251 25467 10257
rect 25409 10248 25421 10251
rect 25372 10220 25421 10248
rect 25372 10208 25378 10220
rect 25409 10217 25421 10220
rect 25455 10217 25467 10251
rect 26418 10248 26424 10260
rect 26379 10220 26424 10248
rect 25409 10211 25467 10217
rect 26418 10208 26424 10220
rect 26476 10208 26482 10260
rect 27982 10248 27988 10260
rect 27943 10220 27988 10248
rect 27982 10208 27988 10220
rect 28040 10208 28046 10260
rect 29362 10208 29368 10260
rect 29420 10248 29426 10260
rect 29549 10251 29607 10257
rect 29549 10248 29561 10251
rect 29420 10220 29561 10248
rect 29420 10208 29426 10220
rect 29549 10217 29561 10220
rect 29595 10217 29607 10251
rect 30650 10248 30656 10260
rect 30611 10220 30656 10248
rect 29549 10211 29607 10217
rect 30650 10208 30656 10220
rect 30708 10208 30714 10260
rect 32490 10248 32496 10260
rect 32451 10220 32496 10248
rect 32490 10208 32496 10220
rect 32548 10208 32554 10260
rect 36630 10208 36636 10260
rect 36688 10248 36694 10260
rect 36817 10251 36875 10257
rect 36817 10248 36829 10251
rect 36688 10220 36829 10248
rect 36688 10208 36694 10220
rect 36817 10217 36829 10220
rect 36863 10217 36875 10251
rect 36817 10211 36875 10217
rect 37461 10251 37519 10257
rect 37461 10217 37473 10251
rect 37507 10248 37519 10251
rect 37918 10248 37924 10260
rect 37507 10220 37924 10248
rect 37507 10217 37519 10220
rect 37461 10211 37519 10217
rect 2501 10183 2559 10189
rect 2501 10149 2513 10183
rect 2547 10149 2559 10183
rect 2501 10143 2559 10149
rect 9600 10152 10548 10180
rect 1765 10047 1823 10053
rect 1765 10013 1777 10047
rect 1811 10013 1823 10047
rect 1765 10007 1823 10013
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10044 1915 10047
rect 2516 10044 2544 10143
rect 3145 10115 3203 10121
rect 3145 10081 3157 10115
rect 3191 10112 3203 10115
rect 3694 10112 3700 10124
rect 3191 10084 3700 10112
rect 3191 10081 3203 10084
rect 3145 10075 3203 10081
rect 3694 10072 3700 10084
rect 3752 10112 3758 10124
rect 5166 10112 5172 10124
rect 3752 10084 5172 10112
rect 3752 10072 3758 10084
rect 5166 10072 5172 10084
rect 5224 10112 5230 10124
rect 9600 10121 9628 10152
rect 9585 10115 9643 10121
rect 9585 10112 9597 10115
rect 5224 10084 9597 10112
rect 5224 10072 5230 10084
rect 9585 10081 9597 10084
rect 9631 10081 9643 10115
rect 9585 10075 9643 10081
rect 9674 10072 9680 10124
rect 9732 10112 9738 10124
rect 10413 10115 10471 10121
rect 10413 10112 10425 10115
rect 9732 10084 10425 10112
rect 9732 10072 9738 10084
rect 10413 10081 10425 10084
rect 10459 10081 10471 10115
rect 10520 10112 10548 10152
rect 10594 10140 10600 10192
rect 10652 10180 10658 10192
rect 15194 10180 15200 10192
rect 10652 10152 15200 10180
rect 10652 10140 10658 10152
rect 15194 10140 15200 10152
rect 15252 10140 15258 10192
rect 19610 10140 19616 10192
rect 19668 10180 19674 10192
rect 23845 10183 23903 10189
rect 23845 10180 23857 10183
rect 19668 10152 23857 10180
rect 19668 10140 19674 10152
rect 23845 10149 23857 10152
rect 23891 10180 23903 10183
rect 27706 10180 27712 10192
rect 23891 10152 27712 10180
rect 23891 10149 23903 10152
rect 23845 10143 23903 10149
rect 13173 10115 13231 10121
rect 13173 10112 13185 10115
rect 10520 10084 13185 10112
rect 10413 10075 10471 10081
rect 13173 10081 13185 10084
rect 13219 10081 13231 10115
rect 13173 10075 13231 10081
rect 1903 10016 2544 10044
rect 1903 10013 1915 10016
rect 1857 10007 1915 10013
rect 1780 9976 1808 10007
rect 3602 10004 3608 10056
rect 3660 10044 3666 10056
rect 6917 10047 6975 10053
rect 6917 10044 6929 10047
rect 3660 10016 6929 10044
rect 3660 10004 3666 10016
rect 6917 10013 6929 10016
rect 6963 10013 6975 10047
rect 6917 10007 6975 10013
rect 9309 10047 9367 10053
rect 9309 10013 9321 10047
rect 9355 10044 9367 10047
rect 10226 10044 10232 10056
rect 9355 10016 10232 10044
rect 9355 10013 9367 10016
rect 9309 10007 9367 10013
rect 2222 9976 2228 9988
rect 1780 9948 2228 9976
rect 2222 9936 2228 9948
rect 2280 9976 2286 9988
rect 2682 9976 2688 9988
rect 2280 9948 2688 9976
rect 2280 9936 2286 9948
rect 2682 9936 2688 9948
rect 2740 9936 2746 9988
rect 2869 9979 2927 9985
rect 2869 9945 2881 9979
rect 2915 9976 2927 9979
rect 4982 9976 4988 9988
rect 2915 9948 3924 9976
rect 4943 9948 4988 9976
rect 2915 9945 2927 9948
rect 2869 9939 2927 9945
rect 3896 9920 3924 9948
rect 4982 9936 4988 9948
rect 5040 9936 5046 9988
rect 6932 9976 6960 10007
rect 10226 10004 10232 10016
rect 10284 10004 10290 10056
rect 10428 10044 10456 10075
rect 16574 10072 16580 10124
rect 16632 10112 16638 10124
rect 20438 10112 20444 10124
rect 16632 10084 20444 10112
rect 16632 10072 16638 10084
rect 20438 10072 20444 10084
rect 20496 10072 20502 10124
rect 21266 10072 21272 10124
rect 21324 10112 21330 10124
rect 21821 10115 21879 10121
rect 21821 10112 21833 10115
rect 21324 10084 21833 10112
rect 21324 10072 21330 10084
rect 21821 10081 21833 10084
rect 21867 10081 21879 10115
rect 21821 10075 21879 10081
rect 24302 10072 24308 10124
rect 24360 10112 24366 10124
rect 24360 10084 25084 10112
rect 24360 10072 24366 10084
rect 10594 10044 10600 10056
rect 10428 10016 10600 10044
rect 10594 10004 10600 10016
rect 10652 10004 10658 10056
rect 12161 10047 12219 10053
rect 12161 10013 12173 10047
rect 12207 10044 12219 10047
rect 12802 10044 12808 10056
rect 12207 10016 12808 10044
rect 12207 10013 12219 10016
rect 12161 10007 12219 10013
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 15562 10004 15568 10056
rect 15620 10044 15626 10056
rect 16758 10044 16764 10056
rect 15620 10016 16764 10044
rect 15620 10004 15626 10016
rect 16758 10004 16764 10016
rect 16816 10004 16822 10056
rect 22005 10047 22063 10053
rect 22005 10013 22017 10047
rect 22051 10044 22063 10047
rect 22094 10044 22100 10056
rect 22051 10016 22100 10044
rect 22051 10013 22063 10016
rect 22005 10007 22063 10013
rect 22094 10004 22100 10016
rect 22152 10044 22158 10056
rect 23382 10044 23388 10056
rect 22152 10016 23388 10044
rect 22152 10004 22158 10016
rect 23382 10004 23388 10016
rect 23440 10004 23446 10056
rect 24026 10004 24032 10056
rect 24084 10044 24090 10056
rect 24765 10047 24823 10053
rect 24765 10044 24777 10047
rect 24084 10016 24777 10044
rect 24084 10004 24090 10016
rect 24765 10013 24777 10016
rect 24811 10013 24823 10047
rect 24946 10044 24952 10056
rect 24907 10016 24952 10044
rect 24765 10007 24823 10013
rect 24946 10004 24952 10016
rect 25004 10004 25010 10056
rect 25056 10053 25084 10084
rect 25148 10053 25176 10152
rect 27706 10140 27712 10152
rect 27764 10140 27770 10192
rect 28626 10140 28632 10192
rect 28684 10140 28690 10192
rect 28997 10183 29055 10189
rect 28997 10149 29009 10183
rect 29043 10180 29055 10183
rect 29270 10180 29276 10192
rect 29043 10152 29276 10180
rect 29043 10149 29055 10152
rect 28997 10143 29055 10149
rect 29270 10140 29276 10152
rect 29328 10140 29334 10192
rect 28258 10112 28264 10124
rect 27632 10084 28264 10112
rect 25041 10047 25099 10053
rect 25041 10013 25053 10047
rect 25087 10013 25099 10047
rect 25041 10007 25099 10013
rect 25133 10047 25191 10053
rect 25133 10013 25145 10047
rect 25179 10013 25191 10047
rect 25133 10007 25191 10013
rect 25869 10047 25927 10053
rect 25869 10013 25881 10047
rect 25915 10013 25927 10047
rect 25869 10007 25927 10013
rect 11514 9976 11520 9988
rect 6932 9948 11520 9976
rect 11514 9936 11520 9948
rect 11572 9936 11578 9988
rect 12434 9936 12440 9988
rect 12492 9976 12498 9988
rect 12989 9979 13047 9985
rect 12989 9976 13001 9979
rect 12492 9948 13001 9976
rect 12492 9936 12498 9948
rect 12989 9945 13001 9948
rect 13035 9945 13047 9979
rect 12989 9939 13047 9945
rect 20714 9936 20720 9988
rect 20772 9976 20778 9988
rect 25884 9976 25912 10007
rect 25958 10004 25964 10056
rect 26016 10044 26022 10056
rect 26145 10047 26203 10053
rect 26145 10044 26157 10047
rect 26016 10016 26157 10044
rect 26016 10004 26022 10016
rect 26145 10013 26157 10016
rect 26191 10013 26203 10047
rect 26145 10007 26203 10013
rect 26234 10004 26240 10056
rect 26292 10044 26298 10056
rect 27430 10044 27436 10056
rect 26292 10016 26337 10044
rect 27391 10016 27436 10044
rect 26292 10004 26298 10016
rect 27430 10004 27436 10016
rect 27488 10004 27494 10056
rect 27632 10053 27660 10084
rect 28258 10072 28264 10084
rect 28316 10072 28322 10124
rect 27617 10047 27675 10053
rect 27617 10013 27629 10047
rect 27663 10013 27675 10047
rect 27798 10044 27804 10056
rect 27759 10016 27804 10044
rect 27617 10007 27675 10013
rect 27798 10004 27804 10016
rect 27856 10004 27862 10056
rect 28442 10044 28448 10056
rect 28403 10016 28448 10044
rect 28442 10004 28448 10016
rect 28500 10004 28506 10056
rect 28644 10053 28672 10140
rect 28629 10047 28687 10053
rect 28629 10013 28641 10047
rect 28675 10013 28687 10047
rect 28810 10044 28816 10056
rect 28771 10016 28816 10044
rect 28629 10007 28687 10013
rect 28810 10004 28816 10016
rect 28868 10004 28874 10056
rect 30650 10004 30656 10056
rect 30708 10044 30714 10056
rect 31205 10047 31263 10053
rect 31205 10044 31217 10047
rect 30708 10016 31217 10044
rect 30708 10004 30714 10016
rect 31205 10013 31217 10016
rect 31251 10013 31263 10047
rect 36832 10044 36860 10211
rect 37918 10208 37924 10220
rect 37976 10208 37982 10260
rect 39022 10112 39028 10124
rect 38212 10084 39028 10112
rect 37090 10044 37096 10056
rect 36832 10016 37096 10044
rect 31205 10007 31263 10013
rect 37090 10004 37096 10016
rect 37148 10044 37154 10056
rect 37921 10047 37979 10053
rect 37921 10044 37933 10047
rect 37148 10016 37933 10044
rect 37148 10004 37154 10016
rect 37921 10013 37933 10016
rect 37967 10013 37979 10047
rect 38102 10044 38108 10056
rect 38063 10016 38108 10044
rect 37921 10007 37979 10013
rect 38102 10004 38108 10016
rect 38160 10004 38166 10056
rect 38212 10053 38240 10084
rect 39022 10072 39028 10084
rect 39080 10072 39086 10124
rect 38197 10047 38255 10053
rect 38197 10013 38209 10047
rect 38243 10013 38255 10047
rect 38197 10007 38255 10013
rect 38289 10047 38347 10053
rect 38289 10013 38301 10047
rect 38335 10013 38347 10047
rect 38289 10007 38347 10013
rect 20772 9948 25912 9976
rect 26053 9979 26111 9985
rect 20772 9936 20778 9948
rect 26053 9945 26065 9979
rect 26099 9976 26111 9979
rect 27522 9976 27528 9988
rect 26099 9948 27528 9976
rect 26099 9945 26111 9948
rect 26053 9939 26111 9945
rect 2961 9911 3019 9917
rect 2961 9877 2973 9911
rect 3007 9908 3019 9911
rect 3418 9908 3424 9920
rect 3007 9880 3424 9908
rect 3007 9877 3019 9880
rect 2961 9871 3019 9877
rect 3418 9868 3424 9880
rect 3476 9868 3482 9920
rect 3878 9908 3884 9920
rect 3839 9880 3884 9908
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 9401 9911 9459 9917
rect 9401 9877 9413 9911
rect 9447 9908 9459 9911
rect 9674 9908 9680 9920
rect 9447 9880 9680 9908
rect 9447 9877 9459 9880
rect 9401 9871 9459 9877
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 12621 9911 12679 9917
rect 12621 9877 12633 9911
rect 12667 9908 12679 9911
rect 12802 9908 12808 9920
rect 12667 9880 12808 9908
rect 12667 9877 12679 9880
rect 12621 9871 12679 9877
rect 12802 9868 12808 9880
rect 12860 9868 12866 9920
rect 13081 9911 13139 9917
rect 13081 9877 13093 9911
rect 13127 9908 13139 9911
rect 13262 9908 13268 9920
rect 13127 9880 13268 9908
rect 13127 9877 13139 9880
rect 13081 9871 13139 9877
rect 13262 9868 13268 9880
rect 13320 9868 13326 9920
rect 22462 9868 22468 9920
rect 22520 9908 22526 9920
rect 26068 9908 26096 9939
rect 27522 9936 27528 9948
rect 27580 9936 27586 9988
rect 27709 9979 27767 9985
rect 27709 9945 27721 9979
rect 27755 9945 27767 9979
rect 27709 9939 27767 9945
rect 28721 9979 28779 9985
rect 28721 9945 28733 9979
rect 28767 9976 28779 9979
rect 29638 9976 29644 9988
rect 28767 9948 29644 9976
rect 28767 9945 28779 9948
rect 28721 9939 28779 9945
rect 22520 9880 26096 9908
rect 22520 9868 22526 9880
rect 26326 9868 26332 9920
rect 26384 9908 26390 9920
rect 27724 9908 27752 9939
rect 29638 9936 29644 9948
rect 29696 9976 29702 9988
rect 29733 9979 29791 9985
rect 29733 9976 29745 9979
rect 29696 9948 29745 9976
rect 29696 9936 29702 9948
rect 29733 9945 29745 9948
rect 29779 9945 29791 9979
rect 29733 9939 29791 9945
rect 29917 9979 29975 9985
rect 29917 9945 29929 9979
rect 29963 9976 29975 9979
rect 30742 9976 30748 9988
rect 29963 9948 30748 9976
rect 29963 9945 29975 9948
rect 29917 9939 29975 9945
rect 30742 9936 30748 9948
rect 30800 9936 30806 9988
rect 37274 9936 37280 9988
rect 37332 9976 37338 9988
rect 38304 9976 38332 10007
rect 39025 9979 39083 9985
rect 39025 9976 39037 9979
rect 37332 9948 39037 9976
rect 37332 9936 37338 9948
rect 39025 9945 39037 9948
rect 39071 9945 39083 9979
rect 39025 9939 39083 9945
rect 26384 9880 27752 9908
rect 38565 9911 38623 9917
rect 26384 9868 26390 9880
rect 38565 9877 38577 9911
rect 38611 9908 38623 9911
rect 38838 9908 38844 9920
rect 38611 9880 38844 9908
rect 38611 9877 38623 9880
rect 38565 9871 38623 9877
rect 38838 9868 38844 9880
rect 38896 9868 38902 9920
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 15010 9664 15016 9716
rect 15068 9704 15074 9716
rect 15105 9707 15163 9713
rect 15105 9704 15117 9707
rect 15068 9676 15117 9704
rect 15068 9664 15074 9676
rect 15105 9673 15117 9676
rect 15151 9704 15163 9707
rect 15151 9676 15253 9704
rect 20548 9676 20852 9704
rect 15151 9673 15163 9676
rect 15105 9667 15163 9673
rect 2308 9639 2366 9645
rect 2308 9605 2320 9639
rect 2354 9636 2366 9639
rect 2406 9636 2412 9648
rect 2354 9608 2412 9636
rect 2354 9605 2366 9608
rect 2308 9599 2366 9605
rect 2406 9596 2412 9608
rect 2464 9596 2470 9648
rect 10229 9639 10287 9645
rect 10229 9605 10241 9639
rect 10275 9636 10287 9639
rect 10502 9636 10508 9648
rect 10275 9608 10508 9636
rect 10275 9605 10287 9608
rect 10229 9599 10287 9605
rect 10502 9596 10508 9608
rect 10560 9596 10566 9648
rect 15120 9636 15148 9667
rect 20548 9636 20576 9676
rect 15120 9608 20576 9636
rect 20622 9596 20628 9648
rect 20680 9636 20686 9648
rect 20717 9639 20775 9645
rect 20717 9636 20729 9639
rect 20680 9608 20729 9636
rect 20680 9596 20686 9608
rect 20717 9605 20729 9608
rect 20763 9605 20775 9639
rect 20824 9636 20852 9676
rect 24946 9664 24952 9716
rect 25004 9704 25010 9716
rect 25133 9707 25191 9713
rect 25133 9704 25145 9707
rect 25004 9676 25145 9704
rect 25004 9664 25010 9676
rect 25133 9673 25145 9676
rect 25179 9673 25191 9707
rect 25774 9704 25780 9716
rect 25133 9667 25191 9673
rect 25240 9676 25780 9704
rect 22278 9636 22284 9648
rect 20824 9608 22284 9636
rect 20717 9599 20775 9605
rect 22278 9596 22284 9608
rect 22336 9596 22342 9648
rect 22649 9639 22707 9645
rect 22649 9605 22661 9639
rect 22695 9636 22707 9639
rect 23014 9636 23020 9648
rect 22695 9608 23020 9636
rect 22695 9605 22707 9608
rect 22649 9599 22707 9605
rect 23014 9596 23020 9608
rect 23072 9596 23078 9648
rect 5534 9568 5540 9580
rect 5495 9540 5540 9568
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 9674 9528 9680 9580
rect 9732 9568 9738 9580
rect 11977 9571 12035 9577
rect 11977 9568 11989 9571
rect 9732 9540 10548 9568
rect 9732 9528 9738 9540
rect 2041 9503 2099 9509
rect 2041 9469 2053 9503
rect 2087 9469 2099 9503
rect 2041 9463 2099 9469
rect 2056 9364 2084 9463
rect 5626 9460 5632 9512
rect 5684 9500 5690 9512
rect 5813 9503 5871 9509
rect 5813 9500 5825 9503
rect 5684 9472 5825 9500
rect 5684 9460 5690 9472
rect 5813 9469 5825 9472
rect 5859 9500 5871 9503
rect 5902 9500 5908 9512
rect 5859 9472 5908 9500
rect 5859 9469 5871 9472
rect 5813 9463 5871 9469
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 10520 9509 10548 9540
rect 10612 9540 11989 9568
rect 10413 9503 10471 9509
rect 10413 9469 10425 9503
rect 10459 9469 10471 9503
rect 10413 9463 10471 9469
rect 10505 9503 10563 9509
rect 10505 9469 10517 9503
rect 10551 9469 10563 9503
rect 10505 9463 10563 9469
rect 10428 9432 10456 9463
rect 10612 9444 10640 9540
rect 11977 9537 11989 9540
rect 12023 9537 12035 9571
rect 12618 9568 12624 9580
rect 12579 9540 12624 9568
rect 11977 9531 12035 9537
rect 12618 9528 12624 9540
rect 12676 9528 12682 9580
rect 12802 9568 12808 9580
rect 12763 9540 12808 9568
rect 12802 9528 12808 9540
rect 12860 9528 12866 9580
rect 14921 9571 14979 9577
rect 14921 9537 14933 9571
rect 14967 9568 14979 9571
rect 17313 9571 17371 9577
rect 17313 9568 17325 9571
rect 14967 9540 15001 9568
rect 16776 9540 17325 9568
rect 14967 9537 14979 9540
rect 14921 9531 14979 9537
rect 10778 9460 10784 9512
rect 10836 9500 10842 9512
rect 10873 9503 10931 9509
rect 10873 9500 10885 9503
rect 10836 9472 10885 9500
rect 10836 9460 10842 9472
rect 10873 9469 10885 9472
rect 10919 9500 10931 9503
rect 11517 9503 11575 9509
rect 11517 9500 11529 9503
rect 10919 9472 11529 9500
rect 10919 9469 10931 9472
rect 10873 9463 10931 9469
rect 11517 9469 11529 9472
rect 11563 9469 11575 9503
rect 11517 9463 11575 9469
rect 11885 9503 11943 9509
rect 11885 9469 11897 9503
rect 11931 9469 11943 9503
rect 11885 9463 11943 9469
rect 14461 9503 14519 9509
rect 14461 9469 14473 9503
rect 14507 9500 14519 9503
rect 14936 9500 14964 9531
rect 15286 9500 15292 9512
rect 14507 9472 15292 9500
rect 14507 9469 14519 9472
rect 14461 9463 14519 9469
rect 10594 9432 10600 9444
rect 10428 9404 10600 9432
rect 10594 9392 10600 9404
rect 10652 9392 10658 9444
rect 11900 9432 11928 9463
rect 15286 9460 15292 9472
rect 15344 9460 15350 9512
rect 13262 9432 13268 9444
rect 11900 9404 13268 9432
rect 13262 9392 13268 9404
rect 13320 9392 13326 9444
rect 15194 9392 15200 9444
rect 15252 9432 15258 9444
rect 16776 9441 16804 9540
rect 17313 9537 17325 9540
rect 17359 9537 17371 9571
rect 17313 9531 17371 9537
rect 20162 9528 20168 9580
rect 20220 9568 20226 9580
rect 22373 9571 22431 9577
rect 22373 9568 22385 9571
rect 20220 9540 22385 9568
rect 20220 9528 20226 9540
rect 22373 9537 22385 9540
rect 22419 9537 22431 9571
rect 22373 9531 22431 9537
rect 22462 9528 22468 9580
rect 22520 9568 22526 9580
rect 22557 9571 22615 9577
rect 22557 9568 22569 9571
rect 22520 9540 22569 9568
rect 22520 9528 22526 9540
rect 22557 9537 22569 9540
rect 22603 9537 22615 9571
rect 22738 9568 22744 9580
rect 22699 9540 22744 9568
rect 22557 9531 22615 9537
rect 22738 9528 22744 9540
rect 22796 9528 22802 9580
rect 24489 9571 24547 9577
rect 24489 9537 24501 9571
rect 24535 9568 24547 9571
rect 25240 9568 25268 9676
rect 25774 9664 25780 9676
rect 25832 9664 25838 9716
rect 29638 9704 29644 9716
rect 29599 9676 29644 9704
rect 29638 9664 29644 9676
rect 29696 9664 29702 9716
rect 30834 9664 30840 9716
rect 30892 9704 30898 9716
rect 31570 9704 31576 9716
rect 30892 9676 31576 9704
rect 30892 9664 30898 9676
rect 31570 9664 31576 9676
rect 31628 9664 31634 9716
rect 37829 9707 37887 9713
rect 37829 9673 37841 9707
rect 37875 9704 37887 9707
rect 38102 9704 38108 9716
rect 37875 9676 38108 9704
rect 37875 9673 37887 9676
rect 37829 9667 37887 9673
rect 38102 9664 38108 9676
rect 38160 9664 38166 9716
rect 25317 9639 25375 9645
rect 25317 9605 25329 9639
rect 25363 9636 25375 9639
rect 26326 9636 26332 9648
rect 25363 9608 26332 9636
rect 25363 9605 25375 9608
rect 25317 9599 25375 9605
rect 26326 9596 26332 9608
rect 26384 9596 26390 9648
rect 29822 9636 29828 9648
rect 28276 9608 29828 9636
rect 28276 9577 28304 9608
rect 29822 9596 29828 9608
rect 29880 9596 29886 9648
rect 31846 9596 31852 9648
rect 31904 9636 31910 9648
rect 32858 9636 32864 9648
rect 31904 9608 32444 9636
rect 31904 9596 31910 9608
rect 28534 9577 28540 9580
rect 24535 9540 25268 9568
rect 25501 9571 25559 9577
rect 24535 9537 24547 9540
rect 24489 9531 24547 9537
rect 25501 9537 25513 9571
rect 25547 9537 25559 9571
rect 25501 9531 25559 9537
rect 28261 9571 28319 9577
rect 28261 9537 28273 9571
rect 28307 9537 28319 9571
rect 28528 9568 28540 9577
rect 28495 9540 28540 9568
rect 28261 9531 28319 9537
rect 28528 9531 28540 9540
rect 19061 9503 19119 9509
rect 19061 9469 19073 9503
rect 19107 9500 19119 9503
rect 19242 9500 19248 9512
rect 19107 9472 19248 9500
rect 19107 9469 19119 9472
rect 19061 9463 19119 9469
rect 19242 9460 19248 9472
rect 19300 9460 19306 9512
rect 16761 9435 16819 9441
rect 16761 9432 16773 9435
rect 15252 9404 16773 9432
rect 15252 9392 15258 9404
rect 16761 9401 16773 9404
rect 16807 9401 16819 9435
rect 22922 9432 22928 9444
rect 22883 9404 22928 9432
rect 16761 9395 16819 9401
rect 22922 9392 22928 9404
rect 22980 9392 22986 9444
rect 24673 9435 24731 9441
rect 24673 9401 24685 9435
rect 24719 9432 24731 9435
rect 25516 9432 25544 9531
rect 28534 9528 28540 9531
rect 28592 9528 28598 9580
rect 29840 9568 29868 9596
rect 30466 9577 30472 9580
rect 30193 9571 30251 9577
rect 30193 9568 30205 9571
rect 29840 9540 30205 9568
rect 30193 9537 30205 9540
rect 30239 9537 30251 9571
rect 30460 9568 30472 9577
rect 30427 9540 30472 9568
rect 30193 9531 30251 9537
rect 30460 9531 30472 9540
rect 30466 9528 30472 9531
rect 30524 9528 30530 9580
rect 32030 9528 32036 9580
rect 32088 9568 32094 9580
rect 32125 9571 32183 9577
rect 32125 9568 32137 9571
rect 32088 9540 32137 9568
rect 32088 9528 32094 9540
rect 32125 9537 32137 9540
rect 32171 9537 32183 9571
rect 32306 9568 32312 9580
rect 32267 9540 32312 9568
rect 32125 9531 32183 9537
rect 32306 9528 32312 9540
rect 32364 9528 32370 9580
rect 32416 9577 32444 9608
rect 32508 9608 32864 9636
rect 32508 9577 32536 9608
rect 32858 9596 32864 9608
rect 32916 9636 32922 9648
rect 33229 9639 33287 9645
rect 33229 9636 33241 9639
rect 32916 9608 33241 9636
rect 32916 9596 32922 9608
rect 33229 9605 33241 9608
rect 33275 9605 33287 9639
rect 33229 9599 33287 9605
rect 34790 9596 34796 9648
rect 34848 9636 34854 9648
rect 38930 9636 38936 9648
rect 34848 9608 38936 9636
rect 34848 9596 34854 9608
rect 38930 9596 38936 9608
rect 38988 9636 38994 9648
rect 38988 9608 39712 9636
rect 38988 9596 38994 9608
rect 32401 9571 32459 9577
rect 32401 9537 32413 9571
rect 32447 9537 32459 9571
rect 32401 9531 32459 9537
rect 32493 9571 32551 9577
rect 32493 9537 32505 9571
rect 32539 9537 32551 9571
rect 32493 9531 32551 9537
rect 34698 9528 34704 9580
rect 34756 9568 34762 9580
rect 35253 9571 35311 9577
rect 35253 9568 35265 9571
rect 34756 9540 35265 9568
rect 34756 9528 34762 9540
rect 35253 9537 35265 9540
rect 35299 9568 35311 9571
rect 35437 9571 35495 9577
rect 35299 9540 35388 9568
rect 35299 9537 35311 9540
rect 35253 9531 35311 9537
rect 25774 9432 25780 9444
rect 24719 9404 25780 9432
rect 24719 9401 24731 9404
rect 24673 9395 24731 9401
rect 25774 9392 25780 9404
rect 25832 9392 25838 9444
rect 34514 9432 34520 9444
rect 31726 9404 34520 9432
rect 2314 9364 2320 9376
rect 2056 9336 2320 9364
rect 2314 9324 2320 9336
rect 2372 9324 2378 9376
rect 3418 9364 3424 9376
rect 3379 9336 3424 9364
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 6270 9324 6276 9376
rect 6328 9364 6334 9376
rect 6365 9367 6423 9373
rect 6365 9364 6377 9367
rect 6328 9336 6377 9364
rect 6328 9324 6334 9336
rect 6365 9333 6377 9336
rect 6411 9333 6423 9367
rect 6365 9327 6423 9333
rect 11698 9324 11704 9376
rect 11756 9364 11762 9376
rect 12161 9367 12219 9373
rect 12161 9364 12173 9367
rect 11756 9336 12173 9364
rect 11756 9324 11762 9336
rect 12161 9333 12173 9336
rect 12207 9333 12219 9367
rect 12161 9327 12219 9333
rect 12989 9367 13047 9373
rect 12989 9333 13001 9367
rect 13035 9364 13047 9367
rect 13078 9364 13084 9376
rect 13035 9336 13084 9364
rect 13035 9333 13047 9336
rect 12989 9327 13047 9333
rect 13078 9324 13084 9336
rect 13136 9324 13142 9376
rect 15654 9364 15660 9376
rect 15615 9336 15660 9364
rect 15654 9324 15660 9336
rect 15712 9324 15718 9376
rect 22738 9324 22744 9376
rect 22796 9364 22802 9376
rect 26234 9364 26240 9376
rect 22796 9336 26240 9364
rect 22796 9324 22802 9336
rect 26234 9324 26240 9336
rect 26292 9324 26298 9376
rect 27062 9324 27068 9376
rect 27120 9364 27126 9376
rect 31726 9364 31754 9404
rect 34514 9392 34520 9404
rect 34572 9432 34578 9444
rect 35250 9432 35256 9444
rect 34572 9404 35256 9432
rect 34572 9392 34578 9404
rect 35250 9392 35256 9404
rect 35308 9392 35314 9444
rect 35360 9432 35388 9540
rect 35437 9537 35449 9571
rect 35483 9568 35495 9571
rect 35618 9568 35624 9580
rect 35483 9540 35624 9568
rect 35483 9537 35495 9540
rect 35437 9531 35495 9537
rect 35618 9528 35624 9540
rect 35676 9528 35682 9580
rect 37461 9571 37519 9577
rect 37461 9537 37473 9571
rect 37507 9568 37519 9571
rect 37550 9568 37556 9580
rect 37507 9540 37556 9568
rect 37507 9537 37519 9540
rect 37461 9531 37519 9537
rect 37550 9528 37556 9540
rect 37608 9528 37614 9580
rect 37645 9571 37703 9577
rect 37645 9537 37657 9571
rect 37691 9537 37703 9571
rect 37645 9531 37703 9537
rect 37366 9460 37372 9512
rect 37424 9500 37430 9512
rect 37660 9500 37688 9531
rect 38838 9528 38844 9580
rect 38896 9568 38902 9580
rect 39684 9577 39712 9608
rect 39402 9571 39460 9577
rect 39402 9568 39414 9571
rect 38896 9540 39414 9568
rect 38896 9528 38902 9540
rect 39402 9537 39414 9540
rect 39448 9537 39460 9571
rect 39402 9531 39460 9537
rect 39669 9571 39727 9577
rect 39669 9537 39681 9571
rect 39715 9537 39727 9571
rect 39669 9531 39727 9537
rect 37424 9472 38332 9500
rect 37424 9460 37430 9472
rect 37734 9432 37740 9444
rect 35360 9404 37740 9432
rect 37734 9392 37740 9404
rect 37792 9392 37798 9444
rect 38304 9441 38332 9472
rect 38289 9435 38347 9441
rect 38289 9401 38301 9435
rect 38335 9401 38347 9435
rect 38289 9395 38347 9401
rect 27120 9336 31754 9364
rect 27120 9324 27126 9336
rect 32674 9324 32680 9376
rect 32732 9364 32738 9376
rect 32769 9367 32827 9373
rect 32769 9364 32781 9367
rect 32732 9336 32781 9364
rect 32732 9324 32738 9336
rect 32769 9333 32781 9336
rect 32815 9333 32827 9367
rect 32769 9327 32827 9333
rect 35434 9324 35440 9376
rect 35492 9364 35498 9376
rect 35621 9367 35679 9373
rect 35621 9364 35633 9367
rect 35492 9336 35633 9364
rect 35492 9324 35498 9336
rect 35621 9333 35633 9336
rect 35667 9333 35679 9367
rect 35621 9327 35679 9333
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 5261 9163 5319 9169
rect 5261 9129 5273 9163
rect 5307 9160 5319 9163
rect 9398 9160 9404 9172
rect 5307 9132 9404 9160
rect 5307 9129 5319 9132
rect 5261 9123 5319 9129
rect 9398 9120 9404 9132
rect 9456 9120 9462 9172
rect 9674 9120 9680 9172
rect 9732 9160 9738 9172
rect 12710 9160 12716 9172
rect 9732 9132 12716 9160
rect 9732 9120 9738 9132
rect 12710 9120 12716 9132
rect 12768 9120 12774 9172
rect 13262 9120 13268 9172
rect 13320 9160 13326 9172
rect 14093 9163 14151 9169
rect 14093 9160 14105 9163
rect 13320 9132 14105 9160
rect 13320 9120 13326 9132
rect 14093 9129 14105 9132
rect 14139 9129 14151 9163
rect 14093 9123 14151 9129
rect 14274 9120 14280 9172
rect 14332 9160 14338 9172
rect 14734 9160 14740 9172
rect 14332 9132 14740 9160
rect 14332 9120 14338 9132
rect 14734 9120 14740 9132
rect 14792 9160 14798 9172
rect 18598 9160 18604 9172
rect 14792 9132 18604 9160
rect 14792 9120 14798 9132
rect 18598 9120 18604 9132
rect 18656 9120 18662 9172
rect 18966 9120 18972 9172
rect 19024 9160 19030 9172
rect 20530 9160 20536 9172
rect 19024 9132 20536 9160
rect 19024 9120 19030 9132
rect 20530 9120 20536 9132
rect 20588 9120 20594 9172
rect 20625 9163 20683 9169
rect 20625 9129 20637 9163
rect 20671 9160 20683 9163
rect 20714 9160 20720 9172
rect 20671 9132 20720 9160
rect 20671 9129 20683 9132
rect 20625 9123 20683 9129
rect 20714 9120 20720 9132
rect 20772 9120 20778 9172
rect 22278 9120 22284 9172
rect 22336 9160 22342 9172
rect 23385 9163 23443 9169
rect 23385 9160 23397 9163
rect 22336 9132 23397 9160
rect 22336 9120 22342 9132
rect 23385 9129 23397 9132
rect 23431 9160 23443 9163
rect 23658 9160 23664 9172
rect 23431 9132 23664 9160
rect 23431 9129 23443 9132
rect 23385 9123 23443 9129
rect 23658 9120 23664 9132
rect 23716 9160 23722 9172
rect 27062 9160 27068 9172
rect 23716 9132 27068 9160
rect 23716 9120 23722 9132
rect 27062 9120 27068 9132
rect 27120 9120 27126 9172
rect 31205 9163 31263 9169
rect 31205 9129 31217 9163
rect 31251 9160 31263 9163
rect 32306 9160 32312 9172
rect 31251 9132 32312 9160
rect 31251 9129 31263 9132
rect 31205 9123 31263 9129
rect 32306 9120 32312 9132
rect 32364 9120 32370 9172
rect 33229 9163 33287 9169
rect 33229 9129 33241 9163
rect 33275 9160 33287 9163
rect 33502 9160 33508 9172
rect 33275 9132 33508 9160
rect 33275 9129 33287 9132
rect 33229 9123 33287 9129
rect 33502 9120 33508 9132
rect 33560 9120 33566 9172
rect 35618 9120 35624 9172
rect 35676 9160 35682 9172
rect 36081 9163 36139 9169
rect 36081 9160 36093 9163
rect 35676 9132 36093 9160
rect 35676 9120 35682 9132
rect 36081 9129 36093 9132
rect 36127 9129 36139 9163
rect 36081 9123 36139 9129
rect 37826 9120 37832 9172
rect 37884 9160 37890 9172
rect 37921 9163 37979 9169
rect 37921 9160 37933 9163
rect 37884 9132 37933 9160
rect 37884 9120 37890 9132
rect 37921 9129 37933 9132
rect 37967 9129 37979 9163
rect 37921 9123 37979 9129
rect 38930 9120 38936 9172
rect 38988 9160 38994 9172
rect 38988 9132 39344 9160
rect 38988 9120 38994 9132
rect 9582 9092 9588 9104
rect 9543 9064 9588 9092
rect 9582 9052 9588 9064
rect 9640 9052 9646 9104
rect 12250 9052 12256 9104
rect 12308 9092 12314 9104
rect 14458 9092 14464 9104
rect 12308 9064 14464 9092
rect 12308 9052 12314 9064
rect 14458 9052 14464 9064
rect 14516 9052 14522 9104
rect 27798 9052 27804 9104
rect 27856 9092 27862 9104
rect 32217 9095 32275 9101
rect 27856 9064 32076 9092
rect 27856 9052 27862 9064
rect 3418 8984 3424 9036
rect 3476 9024 3482 9036
rect 4985 9027 5043 9033
rect 4985 9024 4997 9027
rect 3476 8996 4997 9024
rect 3476 8984 3482 8996
rect 4985 8993 4997 8996
rect 5031 8993 5043 9027
rect 4985 8987 5043 8993
rect 5718 8984 5724 9036
rect 5776 9024 5782 9036
rect 5813 9027 5871 9033
rect 5813 9024 5825 9027
rect 5776 8996 5825 9024
rect 5776 8984 5782 8996
rect 5813 8993 5825 8996
rect 5859 9024 5871 9027
rect 9306 9024 9312 9036
rect 5859 8996 9312 9024
rect 5859 8993 5871 8996
rect 5813 8987 5871 8993
rect 9306 8984 9312 8996
rect 9364 8984 9370 9036
rect 9600 9024 9628 9052
rect 11698 9024 11704 9036
rect 9600 8996 11560 9024
rect 11659 8996 11704 9024
rect 5074 8956 5080 8968
rect 5035 8928 5080 8956
rect 5074 8916 5080 8928
rect 5132 8956 5138 8968
rect 6641 8959 6699 8965
rect 6641 8956 6653 8959
rect 5132 8928 6653 8956
rect 5132 8916 5138 8928
rect 6641 8925 6653 8928
rect 6687 8956 6699 8959
rect 10594 8956 10600 8968
rect 6687 8928 10600 8956
rect 6687 8925 6699 8928
rect 6641 8919 6699 8925
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 11425 8959 11483 8965
rect 11425 8956 11437 8959
rect 11296 8928 11437 8956
rect 11296 8916 11302 8928
rect 11425 8925 11437 8928
rect 11471 8925 11483 8959
rect 11532 8956 11560 8996
rect 11698 8984 11704 8996
rect 11756 8984 11762 9036
rect 11882 9024 11888 9036
rect 11808 8996 11888 9024
rect 11808 8965 11836 8996
rect 11882 8984 11888 8996
rect 11940 8984 11946 9036
rect 21177 9027 21235 9033
rect 21177 8993 21189 9027
rect 21223 9024 21235 9027
rect 21818 9024 21824 9036
rect 21223 8996 21824 9024
rect 21223 8993 21235 8996
rect 21177 8987 21235 8993
rect 21818 8984 21824 8996
rect 21876 9024 21882 9036
rect 22005 9027 22063 9033
rect 22005 9024 22017 9027
rect 21876 8996 22017 9024
rect 21876 8984 21882 8996
rect 22005 8993 22017 8996
rect 22051 8993 22063 9027
rect 22005 8987 22063 8993
rect 22281 9027 22339 9033
rect 22281 8993 22293 9027
rect 22327 9024 22339 9027
rect 22738 9024 22744 9036
rect 22327 8996 22744 9024
rect 22327 8993 22339 8996
rect 22281 8987 22339 8993
rect 22738 8984 22744 8996
rect 22796 8984 22802 9036
rect 26234 8984 26240 9036
rect 26292 9024 26298 9036
rect 28460 9033 28488 9064
rect 28169 9027 28227 9033
rect 28169 9024 28181 9027
rect 26292 8996 28181 9024
rect 26292 8984 26298 8996
rect 28169 8993 28181 8996
rect 28215 8993 28227 9027
rect 28169 8987 28227 8993
rect 28445 9027 28503 9033
rect 28445 8993 28457 9027
rect 28491 8993 28503 9027
rect 28445 8987 28503 8993
rect 11609 8959 11667 8965
rect 11609 8956 11621 8959
rect 11532 8928 11621 8956
rect 11425 8919 11483 8925
rect 11609 8925 11621 8928
rect 11655 8925 11667 8959
rect 11609 8919 11667 8925
rect 11793 8959 11851 8965
rect 11793 8925 11805 8959
rect 11839 8925 11851 8959
rect 11793 8919 11851 8925
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8956 12035 8959
rect 12250 8956 12256 8968
rect 12023 8928 12256 8956
rect 12023 8925 12035 8928
rect 11977 8919 12035 8925
rect 4617 8891 4675 8897
rect 4617 8857 4629 8891
rect 4663 8888 4675 8891
rect 5534 8888 5540 8900
rect 4663 8860 5540 8888
rect 4663 8857 4675 8860
rect 4617 8851 4675 8857
rect 5534 8848 5540 8860
rect 5592 8848 5598 8900
rect 6457 8891 6515 8897
rect 6457 8857 6469 8891
rect 6503 8888 6515 8891
rect 6914 8888 6920 8900
rect 6503 8860 6920 8888
rect 6503 8857 6515 8860
rect 6457 8851 6515 8857
rect 6914 8848 6920 8860
rect 6972 8888 6978 8900
rect 7466 8888 7472 8900
rect 6972 8860 7472 8888
rect 6972 8848 6978 8860
rect 7466 8848 7472 8860
rect 7524 8848 7530 8900
rect 8754 8848 8760 8900
rect 8812 8888 8818 8900
rect 9214 8888 9220 8900
rect 8812 8860 9220 8888
rect 8812 8848 8818 8860
rect 9214 8848 9220 8860
rect 9272 8888 9278 8900
rect 9401 8891 9459 8897
rect 9401 8888 9413 8891
rect 9272 8860 9413 8888
rect 9272 8848 9278 8860
rect 9401 8857 9413 8860
rect 9447 8857 9459 8891
rect 11624 8888 11652 8919
rect 12250 8916 12256 8928
rect 12308 8916 12314 8968
rect 13078 8956 13084 8968
rect 13039 8928 13084 8956
rect 13078 8916 13084 8928
rect 13136 8916 13142 8968
rect 15378 8916 15384 8968
rect 15436 8956 15442 8968
rect 15473 8959 15531 8965
rect 15473 8956 15485 8959
rect 15436 8928 15485 8956
rect 15436 8916 15442 8928
rect 15473 8925 15485 8928
rect 15519 8956 15531 8959
rect 17313 8959 17371 8965
rect 17313 8956 17325 8959
rect 15519 8928 17325 8956
rect 15519 8925 15531 8928
rect 15473 8919 15531 8925
rect 17313 8925 17325 8928
rect 17359 8956 17371 8959
rect 19242 8956 19248 8968
rect 17359 8928 19248 8956
rect 17359 8925 17371 8928
rect 17313 8919 17371 8925
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 20622 8916 20628 8968
rect 20680 8956 20686 8968
rect 21085 8959 21143 8965
rect 21085 8956 21097 8959
rect 20680 8928 21097 8956
rect 20680 8916 20686 8928
rect 21085 8925 21097 8928
rect 21131 8925 21143 8959
rect 21085 8919 21143 8925
rect 21266 8916 21272 8968
rect 21324 8956 21330 8968
rect 21726 8956 21732 8968
rect 21324 8928 21732 8956
rect 21324 8916 21330 8928
rect 21726 8916 21732 8928
rect 21784 8916 21790 8968
rect 28184 8956 28212 8987
rect 31570 8984 31576 9036
rect 31628 9024 31634 9036
rect 32048 9024 32076 9064
rect 32217 9061 32229 9095
rect 32263 9092 32275 9095
rect 33870 9092 33876 9104
rect 32263 9064 33876 9092
rect 32263 9061 32275 9064
rect 32217 9055 32275 9061
rect 33870 9052 33876 9064
rect 33928 9052 33934 9104
rect 32582 9024 32588 9036
rect 31628 8996 31984 9024
rect 31628 8984 31634 8996
rect 28810 8956 28816 8968
rect 28184 8928 28816 8956
rect 28810 8916 28816 8928
rect 28868 8916 28874 8968
rect 30742 8916 30748 8968
rect 30800 8956 30806 8968
rect 30837 8959 30895 8965
rect 30837 8956 30849 8959
rect 30800 8928 30849 8956
rect 30800 8916 30806 8928
rect 30837 8925 30849 8928
rect 30883 8925 30895 8959
rect 31662 8956 31668 8968
rect 31623 8928 31668 8956
rect 30837 8919 30895 8925
rect 31662 8916 31668 8928
rect 31720 8916 31726 8968
rect 31956 8965 31984 8996
rect 32048 8996 32588 9024
rect 32048 8965 32076 8996
rect 32582 8984 32588 8996
rect 32640 9024 32646 9036
rect 32640 8996 33088 9024
rect 32640 8984 32646 8996
rect 31941 8959 31999 8965
rect 31941 8925 31953 8959
rect 31987 8925 31999 8959
rect 31941 8919 31999 8925
rect 32033 8959 32091 8965
rect 32033 8925 32045 8959
rect 32079 8925 32091 8959
rect 32033 8919 32091 8925
rect 32398 8916 32404 8968
rect 32456 8956 32462 8968
rect 32677 8959 32735 8965
rect 32677 8956 32689 8959
rect 32456 8928 32689 8956
rect 32456 8916 32462 8928
rect 32677 8925 32689 8928
rect 32723 8925 32735 8959
rect 32950 8956 32956 8968
rect 32911 8928 32956 8956
rect 32677 8919 32735 8925
rect 32950 8916 32956 8928
rect 33008 8916 33014 8968
rect 33060 8965 33088 8996
rect 35802 8984 35808 9036
rect 35860 9024 35866 9036
rect 39316 9033 39344 9132
rect 39301 9027 39359 9033
rect 35860 8996 37412 9024
rect 35860 8984 35866 8996
rect 33045 8959 33103 8965
rect 33045 8925 33057 8959
rect 33091 8925 33103 8959
rect 33045 8919 33103 8925
rect 34701 8959 34759 8965
rect 34701 8925 34713 8959
rect 34747 8956 34759 8959
rect 34790 8956 34796 8968
rect 34747 8928 34796 8956
rect 34747 8925 34759 8928
rect 34701 8919 34759 8925
rect 34790 8916 34796 8928
rect 34848 8916 34854 8968
rect 36262 8916 36268 8968
rect 36320 8956 36326 8968
rect 36817 8959 36875 8965
rect 36817 8956 36829 8959
rect 36320 8928 36829 8956
rect 36320 8916 36326 8928
rect 36817 8925 36829 8928
rect 36863 8925 36875 8959
rect 36998 8956 37004 8968
rect 36959 8928 37004 8956
rect 36817 8919 36875 8925
rect 36998 8916 37004 8928
rect 37056 8916 37062 8968
rect 37108 8965 37136 8996
rect 37093 8959 37151 8965
rect 37093 8925 37105 8959
rect 37139 8925 37151 8959
rect 37093 8919 37151 8925
rect 37185 8959 37243 8965
rect 37185 8925 37197 8959
rect 37231 8956 37243 8959
rect 37274 8956 37280 8968
rect 37231 8928 37280 8956
rect 37231 8925 37243 8928
rect 37185 8919 37243 8925
rect 37274 8916 37280 8928
rect 37332 8916 37338 8968
rect 37384 8956 37412 8996
rect 39301 8993 39313 9027
rect 39347 8993 39359 9027
rect 39301 8987 39359 8993
rect 38746 8956 38752 8968
rect 37384 8928 38752 8956
rect 38746 8916 38752 8928
rect 38804 8916 38810 8968
rect 58158 8956 58164 8968
rect 58119 8928 58164 8956
rect 58158 8916 58164 8928
rect 58216 8916 58222 8968
rect 11882 8888 11888 8900
rect 11624 8860 11888 8888
rect 9401 8851 9459 8857
rect 11882 8848 11888 8860
rect 11940 8848 11946 8900
rect 15206 8891 15264 8897
rect 15206 8888 15218 8891
rect 13280 8860 15218 8888
rect 3234 8820 3240 8832
rect 3195 8792 3240 8820
rect 3234 8780 3240 8792
rect 3292 8780 3298 8832
rect 4157 8823 4215 8829
rect 4157 8789 4169 8823
rect 4203 8820 4215 8823
rect 4798 8820 4804 8832
rect 4203 8792 4804 8820
rect 4203 8789 4215 8792
rect 4157 8783 4215 8789
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 7190 8820 7196 8832
rect 7151 8792 7196 8820
rect 7190 8780 7196 8792
rect 7248 8780 7254 8832
rect 7745 8823 7803 8829
rect 7745 8789 7757 8823
rect 7791 8820 7803 8823
rect 8110 8820 8116 8832
rect 7791 8792 8116 8820
rect 7791 8789 7803 8792
rect 7745 8783 7803 8789
rect 8110 8780 8116 8792
rect 8168 8780 8174 8832
rect 9582 8780 9588 8832
rect 9640 8820 9646 8832
rect 10045 8823 10103 8829
rect 10045 8820 10057 8823
rect 9640 8792 10057 8820
rect 9640 8780 9646 8792
rect 10045 8789 10057 8792
rect 10091 8789 10103 8823
rect 10045 8783 10103 8789
rect 11241 8823 11299 8829
rect 11241 8789 11253 8823
rect 11287 8820 11299 8823
rect 12710 8820 12716 8832
rect 11287 8792 12716 8820
rect 11287 8789 11299 8792
rect 11241 8783 11299 8789
rect 12710 8780 12716 8792
rect 12768 8780 12774 8832
rect 13280 8829 13308 8860
rect 15206 8857 15218 8860
rect 15252 8857 15264 8891
rect 15206 8851 15264 8857
rect 17580 8891 17638 8897
rect 17580 8857 17592 8891
rect 17626 8888 17638 8891
rect 17678 8888 17684 8900
rect 17626 8860 17684 8888
rect 17626 8857 17638 8860
rect 17580 8851 17638 8857
rect 17678 8848 17684 8860
rect 17736 8848 17742 8900
rect 18782 8848 18788 8900
rect 18840 8888 18846 8900
rect 19490 8891 19548 8897
rect 19490 8888 19502 8891
rect 18840 8860 19502 8888
rect 18840 8848 18846 8860
rect 19490 8857 19502 8860
rect 19536 8857 19548 8891
rect 19490 8851 19548 8857
rect 31021 8891 31079 8897
rect 31021 8857 31033 8891
rect 31067 8888 31079 8891
rect 31386 8888 31392 8900
rect 31067 8860 31392 8888
rect 31067 8857 31079 8860
rect 31021 8851 31079 8857
rect 31386 8848 31392 8860
rect 31444 8848 31450 8900
rect 31849 8891 31907 8897
rect 31849 8888 31861 8891
rect 31726 8860 31861 8888
rect 13265 8823 13323 8829
rect 13265 8789 13277 8823
rect 13311 8789 13323 8823
rect 13265 8783 13323 8789
rect 16301 8823 16359 8829
rect 16301 8789 16313 8823
rect 16347 8820 16359 8823
rect 16390 8820 16396 8832
rect 16347 8792 16396 8820
rect 16347 8789 16359 8792
rect 16301 8783 16359 8789
rect 16390 8780 16396 8792
rect 16448 8780 16454 8832
rect 16853 8823 16911 8829
rect 16853 8789 16865 8823
rect 16899 8820 16911 8823
rect 17954 8820 17960 8832
rect 16899 8792 17960 8820
rect 16899 8789 16911 8792
rect 16853 8783 16911 8789
rect 17954 8780 17960 8792
rect 18012 8780 18018 8832
rect 18693 8823 18751 8829
rect 18693 8789 18705 8823
rect 18739 8820 18751 8823
rect 20162 8820 20168 8832
rect 18739 8792 20168 8820
rect 18739 8789 18751 8792
rect 18693 8783 18751 8789
rect 20162 8780 20168 8792
rect 20220 8780 20226 8832
rect 28258 8780 28264 8832
rect 28316 8820 28322 8832
rect 31726 8820 31754 8860
rect 31849 8857 31861 8860
rect 31895 8888 31907 8891
rect 32306 8888 32312 8900
rect 31895 8860 32312 8888
rect 31895 8857 31907 8860
rect 31849 8851 31907 8857
rect 32306 8848 32312 8860
rect 32364 8888 32370 8900
rect 34974 8897 34980 8900
rect 32861 8891 32919 8897
rect 32861 8888 32873 8891
rect 32364 8860 32873 8888
rect 32364 8848 32370 8860
rect 32861 8857 32873 8860
rect 32907 8857 32919 8891
rect 32861 8851 32919 8857
rect 34968 8851 34980 8897
rect 35032 8888 35038 8900
rect 37461 8891 37519 8897
rect 35032 8860 35068 8888
rect 34974 8848 34980 8851
rect 35032 8848 35038 8860
rect 37461 8857 37473 8891
rect 37507 8888 37519 8891
rect 39034 8891 39092 8897
rect 39034 8888 39046 8891
rect 37507 8860 39046 8888
rect 37507 8857 37519 8860
rect 37461 8851 37519 8857
rect 39034 8857 39046 8860
rect 39080 8857 39092 8891
rect 39034 8851 39092 8857
rect 28316 8792 31754 8820
rect 28316 8780 28322 8792
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 4982 8576 4988 8628
rect 5040 8616 5046 8628
rect 8202 8616 8208 8628
rect 5040 8588 8208 8616
rect 5040 8576 5046 8588
rect 8202 8576 8208 8588
rect 8260 8616 8266 8628
rect 8757 8619 8815 8625
rect 8757 8616 8769 8619
rect 8260 8588 8769 8616
rect 8260 8576 8266 8588
rect 8757 8585 8769 8588
rect 8803 8585 8815 8619
rect 9674 8616 9680 8628
rect 9635 8588 9680 8616
rect 8757 8579 8815 8585
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 10134 8616 10140 8628
rect 10095 8588 10140 8616
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 13354 8576 13360 8628
rect 13412 8616 13418 8628
rect 13449 8619 13507 8625
rect 13449 8616 13461 8619
rect 13412 8588 13461 8616
rect 13412 8576 13418 8588
rect 13449 8585 13461 8588
rect 13495 8585 13507 8619
rect 13449 8579 13507 8585
rect 14185 8619 14243 8625
rect 14185 8585 14197 8619
rect 14231 8616 14243 8619
rect 14274 8616 14280 8628
rect 14231 8588 14280 8616
rect 14231 8585 14243 8588
rect 14185 8579 14243 8585
rect 7006 8508 7012 8560
rect 7064 8548 7070 8560
rect 9766 8548 9772 8560
rect 7064 8520 9772 8548
rect 7064 8508 7070 8520
rect 9766 8508 9772 8520
rect 9824 8508 9830 8560
rect 5626 8440 5632 8492
rect 5684 8480 5690 8492
rect 6638 8480 6644 8492
rect 5684 8452 6644 8480
rect 5684 8440 5690 8452
rect 6638 8440 6644 8452
rect 6696 8480 6702 8492
rect 8754 8480 8760 8492
rect 6696 8452 8760 8480
rect 6696 8440 6702 8452
rect 8754 8440 8760 8452
rect 8812 8440 8818 8492
rect 10152 8480 10180 8576
rect 12802 8548 12808 8560
rect 12084 8520 12808 8548
rect 8956 8452 10180 8480
rect 5813 8415 5871 8421
rect 5813 8381 5825 8415
rect 5859 8412 5871 8415
rect 5902 8412 5908 8424
rect 5859 8384 5908 8412
rect 5859 8381 5871 8384
rect 5813 8375 5871 8381
rect 5902 8372 5908 8384
rect 5960 8412 5966 8424
rect 6362 8412 6368 8424
rect 5960 8384 6368 8412
rect 5960 8372 5966 8384
rect 6362 8372 6368 8384
rect 6420 8372 6426 8424
rect 8570 8412 8576 8424
rect 8531 8384 8576 8412
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 8956 8421 8984 8452
rect 10870 8440 10876 8492
rect 10928 8480 10934 8492
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 10928 8452 11713 8480
rect 10928 8440 10934 8452
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 11882 8480 11888 8492
rect 11843 8452 11888 8480
rect 11701 8443 11759 8449
rect 11882 8440 11888 8452
rect 11940 8440 11946 8492
rect 12084 8489 12112 8520
rect 12802 8508 12808 8520
rect 12860 8508 12866 8560
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8449 12127 8483
rect 12250 8480 12256 8492
rect 12211 8452 12256 8480
rect 12069 8443 12127 8449
rect 12250 8440 12256 8452
rect 12308 8440 12314 8492
rect 13464 8480 13492 8579
rect 14274 8576 14280 8588
rect 14332 8576 14338 8628
rect 14458 8576 14464 8628
rect 14516 8616 14522 8628
rect 17126 8616 17132 8628
rect 14516 8588 17132 8616
rect 14516 8576 14522 8588
rect 17126 8576 17132 8588
rect 17184 8616 17190 8628
rect 17497 8619 17555 8625
rect 17497 8616 17509 8619
rect 17184 8588 17509 8616
rect 17184 8576 17190 8588
rect 17497 8585 17509 8588
rect 17543 8585 17555 8619
rect 17497 8579 17555 8585
rect 18230 8576 18236 8628
rect 18288 8616 18294 8628
rect 18693 8619 18751 8625
rect 18288 8588 18368 8616
rect 18288 8576 18294 8588
rect 15470 8548 15476 8560
rect 14108 8520 15476 8548
rect 13998 8480 14004 8492
rect 13464 8452 14004 8480
rect 13998 8440 14004 8452
rect 14056 8440 14062 8492
rect 8941 8415 8999 8421
rect 8941 8381 8953 8415
rect 8987 8381 8999 8415
rect 8941 8375 8999 8381
rect 9306 8372 9312 8424
rect 9364 8412 9370 8424
rect 11790 8412 11796 8424
rect 9364 8384 11796 8412
rect 9364 8372 9370 8384
rect 11790 8372 11796 8384
rect 11848 8372 11854 8424
rect 11974 8372 11980 8424
rect 12032 8412 12038 8424
rect 12802 8412 12808 8424
rect 12032 8384 12077 8412
rect 12715 8384 12808 8412
rect 12032 8372 12038 8384
rect 12802 8372 12808 8384
rect 12860 8412 12866 8424
rect 14108 8412 14136 8520
rect 15470 8508 15476 8520
rect 15528 8508 15534 8560
rect 18138 8548 18144 8560
rect 16960 8520 18144 8548
rect 14737 8483 14795 8489
rect 14737 8449 14749 8483
rect 14783 8480 14795 8483
rect 14826 8480 14832 8492
rect 14783 8452 14832 8480
rect 14783 8449 14795 8452
rect 14737 8443 14795 8449
rect 14826 8440 14832 8452
rect 14884 8440 14890 8492
rect 15010 8489 15016 8492
rect 15004 8443 15016 8489
rect 15068 8480 15074 8492
rect 16960 8489 16988 8520
rect 18138 8508 18144 8520
rect 18196 8508 18202 8560
rect 16945 8483 17003 8489
rect 16945 8480 16957 8483
rect 15068 8452 15104 8480
rect 16040 8452 16957 8480
rect 15010 8440 15016 8443
rect 15068 8440 15074 8452
rect 12860 8384 14136 8412
rect 12860 8372 12866 8384
rect 1578 8344 1584 8356
rect 1539 8316 1584 8344
rect 1578 8304 1584 8316
rect 1636 8304 1642 8356
rect 2130 8344 2136 8356
rect 2091 8316 2136 8344
rect 2130 8304 2136 8316
rect 2188 8304 2194 8356
rect 2590 8304 2596 8356
rect 2648 8344 2654 8356
rect 2685 8347 2743 8353
rect 2685 8344 2697 8347
rect 2648 8316 2697 8344
rect 2648 8304 2654 8316
rect 2685 8313 2697 8316
rect 2731 8313 2743 8347
rect 2685 8307 2743 8313
rect 4249 8347 4307 8353
rect 4249 8313 4261 8347
rect 4295 8344 4307 8347
rect 4614 8344 4620 8356
rect 4295 8316 4620 8344
rect 4295 8313 4307 8316
rect 4249 8307 4307 8313
rect 4614 8304 4620 8316
rect 4672 8304 4678 8356
rect 7558 8304 7564 8356
rect 7616 8344 7622 8356
rect 7653 8347 7711 8353
rect 7653 8344 7665 8347
rect 7616 8316 7665 8344
rect 7616 8304 7622 8316
rect 7653 8313 7665 8316
rect 7699 8313 7711 8347
rect 7653 8307 7711 8313
rect 8754 8304 8760 8356
rect 8812 8344 8818 8356
rect 10686 8344 10692 8356
rect 8812 8316 10548 8344
rect 10647 8316 10692 8344
rect 8812 8304 8818 8316
rect 3421 8279 3479 8285
rect 3421 8245 3433 8279
rect 3467 8276 3479 8279
rect 3878 8276 3884 8288
rect 3467 8248 3884 8276
rect 3467 8245 3479 8248
rect 3421 8239 3479 8245
rect 3878 8236 3884 8248
rect 3936 8236 3942 8288
rect 5534 8276 5540 8288
rect 5493 8248 5540 8276
rect 5534 8236 5540 8248
rect 5592 8285 5598 8288
rect 5592 8279 5641 8285
rect 5592 8245 5595 8279
rect 5629 8276 5641 8279
rect 8018 8276 8024 8288
rect 5629 8248 8024 8276
rect 5629 8245 5641 8248
rect 5592 8239 5641 8245
rect 5592 8236 5598 8239
rect 8018 8236 8024 8248
rect 8076 8236 8082 8288
rect 8846 8236 8852 8288
rect 8904 8276 8910 8288
rect 8941 8279 8999 8285
rect 8941 8276 8953 8279
rect 8904 8248 8953 8276
rect 8904 8236 8910 8248
rect 8941 8245 8953 8248
rect 8987 8276 8999 8279
rect 9674 8276 9680 8288
rect 8987 8248 9680 8276
rect 8987 8245 8999 8248
rect 8941 8239 8999 8245
rect 9674 8236 9680 8248
rect 9732 8236 9738 8288
rect 10520 8276 10548 8316
rect 10686 8304 10692 8316
rect 10744 8304 10750 8356
rect 11517 8347 11575 8353
rect 10796 8316 11468 8344
rect 10796 8276 10824 8316
rect 10520 8248 10824 8276
rect 11440 8276 11468 8316
rect 11517 8313 11529 8347
rect 11563 8344 11575 8347
rect 11606 8344 11612 8356
rect 11563 8316 11612 8344
rect 11563 8313 11575 8316
rect 11517 8307 11575 8313
rect 11606 8304 11612 8316
rect 11664 8304 11670 8356
rect 16040 8344 16068 8452
rect 16945 8449 16957 8452
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 17126 8440 17132 8492
rect 17184 8480 17190 8492
rect 18340 8489 18368 8588
rect 18693 8585 18705 8619
rect 18739 8616 18751 8619
rect 18782 8616 18788 8628
rect 18739 8588 18788 8616
rect 18739 8585 18751 8588
rect 18693 8579 18751 8585
rect 18782 8576 18788 8588
rect 18840 8576 18846 8628
rect 20714 8616 20720 8628
rect 19352 8588 20720 8616
rect 19352 8557 19380 8588
rect 20714 8576 20720 8588
rect 20772 8576 20778 8628
rect 20993 8619 21051 8625
rect 20993 8585 21005 8619
rect 21039 8616 21051 8619
rect 21266 8616 21272 8628
rect 21039 8588 21272 8616
rect 21039 8585 21051 8588
rect 20993 8579 21051 8585
rect 21266 8576 21272 8588
rect 21324 8576 21330 8628
rect 29825 8619 29883 8625
rect 29825 8585 29837 8619
rect 29871 8616 29883 8619
rect 30282 8616 30288 8628
rect 29871 8588 30288 8616
rect 29871 8585 29883 8588
rect 29825 8579 29883 8585
rect 30282 8576 30288 8588
rect 30340 8576 30346 8628
rect 32122 8576 32128 8628
rect 32180 8616 32186 8628
rect 32677 8619 32735 8625
rect 32180 8588 32444 8616
rect 32180 8576 32186 8588
rect 19337 8551 19395 8557
rect 19337 8517 19349 8551
rect 19383 8517 19395 8551
rect 20162 8548 20168 8560
rect 20123 8520 20168 8548
rect 19337 8511 19395 8517
rect 20162 8508 20168 8520
rect 20220 8508 20226 8560
rect 24302 8548 24308 8560
rect 23768 8520 24308 8548
rect 18049 8483 18107 8489
rect 18049 8480 18061 8483
rect 17184 8452 18061 8480
rect 17184 8440 17190 8452
rect 18049 8449 18061 8452
rect 18095 8449 18107 8483
rect 18049 8443 18107 8449
rect 18233 8483 18291 8489
rect 18233 8449 18245 8483
rect 18279 8449 18291 8483
rect 18233 8443 18291 8449
rect 18325 8483 18383 8489
rect 18325 8449 18337 8483
rect 18371 8449 18383 8483
rect 18325 8443 18383 8449
rect 16482 8372 16488 8424
rect 16540 8412 16546 8424
rect 17494 8412 17500 8424
rect 16540 8384 17500 8412
rect 16540 8372 16546 8384
rect 17494 8372 17500 8384
rect 17552 8372 17558 8424
rect 18248 8412 18276 8443
rect 18414 8440 18420 8492
rect 18472 8480 18478 8492
rect 18472 8452 18517 8480
rect 18472 8440 18478 8452
rect 18598 8440 18604 8492
rect 18656 8480 18662 8492
rect 18656 8452 19288 8480
rect 18656 8440 18662 8452
rect 19153 8415 19211 8421
rect 19153 8412 19165 8415
rect 18248 8384 19165 8412
rect 19153 8381 19165 8384
rect 19199 8381 19211 8415
rect 19260 8412 19288 8452
rect 19426 8440 19432 8492
rect 19484 8480 19490 8492
rect 19521 8483 19579 8489
rect 19521 8480 19533 8483
rect 19484 8452 19533 8480
rect 19484 8440 19490 8452
rect 19521 8449 19533 8452
rect 19567 8480 19579 8483
rect 20349 8483 20407 8489
rect 20349 8480 20361 8483
rect 19567 8452 20361 8480
rect 19567 8449 19579 8452
rect 19521 8443 19579 8449
rect 20349 8449 20361 8452
rect 20395 8480 20407 8483
rect 21358 8480 21364 8492
rect 20395 8452 21364 8480
rect 20395 8449 20407 8452
rect 20349 8443 20407 8449
rect 21358 8440 21364 8452
rect 21416 8440 21422 8492
rect 21818 8480 21824 8492
rect 21779 8452 21824 8480
rect 21818 8440 21824 8452
rect 21876 8440 21882 8492
rect 22094 8440 22100 8492
rect 22152 8480 22158 8492
rect 22646 8480 22652 8492
rect 22152 8452 22652 8480
rect 22152 8440 22158 8452
rect 22646 8440 22652 8452
rect 22704 8440 22710 8492
rect 23658 8480 23664 8492
rect 23619 8452 23664 8480
rect 23658 8440 23664 8452
rect 23716 8440 23722 8492
rect 23768 8489 23796 8520
rect 24302 8508 24308 8520
rect 24360 8508 24366 8560
rect 28626 8548 28632 8560
rect 28000 8520 28632 8548
rect 23753 8483 23811 8489
rect 23753 8449 23765 8483
rect 23799 8449 23811 8483
rect 23753 8443 23811 8449
rect 23845 8483 23903 8489
rect 23845 8449 23857 8483
rect 23891 8449 23903 8483
rect 24026 8480 24032 8492
rect 23987 8452 24032 8480
rect 23845 8443 23903 8449
rect 19260 8384 22094 8412
rect 19153 8375 19211 8381
rect 12268 8316 14780 8344
rect 12268 8276 12296 8316
rect 11440 8248 12296 8276
rect 14752 8276 14780 8316
rect 15672 8316 16068 8344
rect 16117 8347 16175 8353
rect 15672 8276 15700 8316
rect 16117 8313 16129 8347
rect 16163 8344 16175 8347
rect 16850 8344 16856 8356
rect 16163 8316 16856 8344
rect 16163 8313 16175 8316
rect 16117 8307 16175 8313
rect 16850 8304 16856 8316
rect 16908 8304 16914 8356
rect 18138 8304 18144 8356
rect 18196 8344 18202 8356
rect 19981 8347 20039 8353
rect 19981 8344 19993 8347
rect 18196 8316 19993 8344
rect 18196 8304 18202 8316
rect 19981 8313 19993 8316
rect 20027 8313 20039 8347
rect 22066 8344 22094 8384
rect 23290 8372 23296 8424
rect 23348 8412 23354 8424
rect 23860 8412 23888 8443
rect 24026 8440 24032 8452
rect 24084 8440 24090 8492
rect 27614 8440 27620 8492
rect 27672 8480 27678 8492
rect 28000 8489 28028 8520
rect 28626 8508 28632 8520
rect 28684 8548 28690 8560
rect 29457 8551 29515 8557
rect 29457 8548 29469 8551
rect 28684 8520 29469 8548
rect 28684 8508 28690 8520
rect 29457 8517 29469 8520
rect 29503 8517 29515 8551
rect 29457 8511 29515 8517
rect 29549 8551 29607 8557
rect 29549 8517 29561 8551
rect 29595 8548 29607 8551
rect 31386 8548 31392 8560
rect 29595 8520 31392 8548
rect 29595 8517 29607 8520
rect 29549 8511 29607 8517
rect 31386 8508 31392 8520
rect 31444 8508 31450 8560
rect 32306 8548 32312 8560
rect 32267 8520 32312 8548
rect 32306 8508 32312 8520
rect 32364 8508 32370 8560
rect 32416 8557 32444 8588
rect 32677 8585 32689 8619
rect 32723 8616 32735 8619
rect 33686 8616 33692 8628
rect 32723 8588 33692 8616
rect 32723 8585 32735 8588
rect 32677 8579 32735 8585
rect 33686 8576 33692 8588
rect 33744 8576 33750 8628
rect 34514 8616 34520 8628
rect 34475 8588 34520 8616
rect 34514 8576 34520 8588
rect 34572 8576 34578 8628
rect 34974 8616 34980 8628
rect 34935 8588 34980 8616
rect 34974 8576 34980 8588
rect 35032 8576 35038 8628
rect 36998 8576 37004 8628
rect 37056 8616 37062 8628
rect 37277 8619 37335 8625
rect 37277 8616 37289 8619
rect 37056 8588 37289 8616
rect 37056 8576 37062 8588
rect 37277 8585 37289 8588
rect 37323 8585 37335 8619
rect 37277 8579 37335 8585
rect 32401 8551 32459 8557
rect 32401 8517 32413 8551
rect 32447 8517 32459 8551
rect 32401 8511 32459 8517
rect 27985 8483 28043 8489
rect 27985 8480 27997 8483
rect 27672 8452 27997 8480
rect 27672 8440 27678 8452
rect 27985 8449 27997 8452
rect 28031 8449 28043 8483
rect 28258 8480 28264 8492
rect 28219 8452 28264 8480
rect 27985 8443 28043 8449
rect 28258 8440 28264 8452
rect 28316 8440 28322 8492
rect 29270 8480 29276 8492
rect 29231 8452 29276 8480
rect 29270 8440 29276 8452
rect 29328 8440 29334 8492
rect 29641 8483 29699 8489
rect 29641 8449 29653 8483
rect 29687 8449 29699 8483
rect 32122 8480 32128 8492
rect 32083 8452 32128 8480
rect 29641 8443 29699 8449
rect 23348 8384 23888 8412
rect 23348 8372 23354 8384
rect 28810 8372 28816 8424
rect 28868 8412 28874 8424
rect 29656 8412 29684 8443
rect 32122 8440 32128 8452
rect 32180 8440 32186 8492
rect 32493 8483 32551 8489
rect 32493 8449 32505 8483
rect 32539 8480 32551 8483
rect 32582 8480 32588 8492
rect 32539 8452 32588 8480
rect 32539 8449 32551 8452
rect 32493 8443 32551 8449
rect 32582 8440 32588 8452
rect 32640 8440 32646 8492
rect 34532 8480 34560 8576
rect 35802 8548 35808 8560
rect 35360 8520 35808 8548
rect 35360 8489 35388 8520
rect 35802 8508 35808 8520
rect 35860 8508 35866 8560
rect 37461 8551 37519 8557
rect 37461 8517 37473 8551
rect 37507 8548 37519 8551
rect 37826 8548 37832 8560
rect 37507 8520 37832 8548
rect 37507 8517 37519 8520
rect 37461 8511 37519 8517
rect 37826 8508 37832 8520
rect 37884 8508 37890 8560
rect 35253 8483 35311 8489
rect 35253 8480 35265 8483
rect 34532 8452 35265 8480
rect 35253 8449 35265 8452
rect 35299 8449 35311 8483
rect 35253 8443 35311 8449
rect 35345 8483 35403 8489
rect 35345 8449 35357 8483
rect 35391 8449 35403 8483
rect 35345 8443 35403 8449
rect 35434 8440 35440 8492
rect 35492 8480 35498 8492
rect 35621 8483 35679 8489
rect 35492 8452 35537 8480
rect 35492 8440 35498 8452
rect 35621 8449 35633 8483
rect 35667 8480 35679 8483
rect 36262 8480 36268 8492
rect 35667 8452 36268 8480
rect 35667 8449 35679 8452
rect 35621 8443 35679 8449
rect 36262 8440 36268 8452
rect 36320 8440 36326 8492
rect 36725 8483 36783 8489
rect 36725 8449 36737 8483
rect 36771 8480 36783 8483
rect 37645 8483 37703 8489
rect 36771 8452 37274 8480
rect 36771 8449 36783 8452
rect 36725 8443 36783 8449
rect 28868 8384 29684 8412
rect 28868 8372 28874 8384
rect 23474 8344 23480 8356
rect 22066 8316 23480 8344
rect 19981 8307 20039 8313
rect 23474 8304 23480 8316
rect 23532 8304 23538 8356
rect 27614 8304 27620 8356
rect 27672 8344 27678 8356
rect 27890 8344 27896 8356
rect 27672 8316 27896 8344
rect 27672 8304 27678 8316
rect 27890 8304 27896 8316
rect 27948 8344 27954 8356
rect 36740 8344 36768 8443
rect 37246 8424 37274 8452
rect 37645 8449 37657 8483
rect 37691 8480 37703 8483
rect 37734 8480 37740 8492
rect 37691 8452 37740 8480
rect 37691 8449 37703 8452
rect 37645 8443 37703 8449
rect 37734 8440 37740 8452
rect 37792 8440 37798 8492
rect 37246 8384 37280 8424
rect 37274 8372 37280 8384
rect 37332 8372 37338 8424
rect 27948 8316 36768 8344
rect 27948 8304 27954 8316
rect 14752 8248 15700 8276
rect 23198 8236 23204 8288
rect 23256 8276 23262 8288
rect 23385 8279 23443 8285
rect 23385 8276 23397 8279
rect 23256 8248 23397 8276
rect 23256 8236 23262 8248
rect 23385 8245 23397 8248
rect 23431 8245 23443 8279
rect 23385 8239 23443 8245
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 9582 8032 9588 8084
rect 9640 8072 9646 8084
rect 10781 8075 10839 8081
rect 9640 8032 9674 8072
rect 10781 8041 10793 8075
rect 10827 8072 10839 8075
rect 11974 8072 11980 8084
rect 10827 8044 11980 8072
rect 10827 8041 10839 8044
rect 10781 8035 10839 8041
rect 11974 8032 11980 8044
rect 12032 8032 12038 8084
rect 14277 8075 14335 8081
rect 14277 8041 14289 8075
rect 14323 8072 14335 8075
rect 17126 8072 17132 8084
rect 14323 8044 16988 8072
rect 17087 8044 17132 8072
rect 14323 8041 14335 8044
rect 14277 8035 14335 8041
rect 3418 7964 3424 8016
rect 3476 8004 3482 8016
rect 4706 8004 4712 8016
rect 3476 7976 4712 8004
rect 3476 7964 3482 7976
rect 4706 7964 4712 7976
rect 4764 7964 4770 8016
rect 5626 8004 5632 8016
rect 5092 7976 5632 8004
rect 3145 7939 3203 7945
rect 3145 7905 3157 7939
rect 3191 7936 3203 7939
rect 4982 7936 4988 7948
rect 3191 7908 4988 7936
rect 3191 7905 3203 7908
rect 3145 7899 3203 7905
rect 4982 7896 4988 7908
rect 5040 7896 5046 7948
rect 5092 7945 5120 7976
rect 5626 7964 5632 7976
rect 5684 7964 5690 8016
rect 7285 8007 7343 8013
rect 7285 7973 7297 8007
rect 7331 8004 7343 8007
rect 7926 8004 7932 8016
rect 7331 7976 7932 8004
rect 7331 7973 7343 7976
rect 7285 7967 7343 7973
rect 7926 7964 7932 7976
rect 7984 8004 7990 8016
rect 9646 8004 9674 8032
rect 13541 8007 13599 8013
rect 7984 7976 8156 8004
rect 9646 7976 10088 8004
rect 7984 7964 7990 7976
rect 5077 7939 5135 7945
rect 5077 7905 5089 7939
rect 5123 7905 5135 7939
rect 5718 7936 5724 7948
rect 5077 7899 5135 7905
rect 5276 7908 5724 7936
rect 2869 7871 2927 7877
rect 2869 7837 2881 7871
rect 2915 7868 2927 7871
rect 3878 7868 3884 7880
rect 2915 7840 3884 7868
rect 2915 7837 2927 7840
rect 2869 7831 2927 7837
rect 3878 7828 3884 7840
rect 3936 7828 3942 7880
rect 4062 7828 4068 7880
rect 4120 7868 4126 7880
rect 5276 7877 5304 7908
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 8128 7945 8156 7976
rect 8113 7939 8171 7945
rect 8113 7905 8125 7939
rect 8159 7905 8171 7939
rect 8113 7899 8171 7905
rect 8389 7939 8447 7945
rect 8389 7905 8401 7939
rect 8435 7936 8447 7939
rect 9401 7939 9459 7945
rect 9401 7936 9413 7939
rect 8435 7908 9413 7936
rect 8435 7905 8447 7908
rect 8389 7899 8447 7905
rect 9401 7905 9413 7908
rect 9447 7905 9459 7939
rect 9401 7899 9459 7905
rect 4893 7871 4951 7877
rect 4893 7868 4905 7871
rect 4120 7840 4905 7868
rect 4120 7828 4126 7840
rect 4893 7837 4905 7840
rect 4939 7837 4951 7871
rect 4893 7831 4951 7837
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7837 5319 7871
rect 5442 7868 5448 7880
rect 5403 7840 5448 7868
rect 5261 7831 5319 7837
rect 2041 7803 2099 7809
rect 2041 7769 2053 7803
rect 2087 7800 2099 7803
rect 2682 7800 2688 7812
rect 2087 7772 2688 7800
rect 2087 7769 2099 7772
rect 2041 7763 2099 7769
rect 2682 7760 2688 7772
rect 2740 7760 2746 7812
rect 5184 7744 5212 7831
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 5905 7871 5963 7877
rect 5905 7837 5917 7871
rect 5951 7868 5963 7871
rect 6730 7868 6736 7880
rect 5951 7840 6736 7868
rect 5951 7837 5963 7840
rect 5905 7831 5963 7837
rect 6730 7828 6736 7840
rect 6788 7828 6794 7880
rect 7466 7828 7472 7880
rect 7524 7868 7530 7880
rect 8205 7871 8263 7877
rect 8205 7868 8217 7871
rect 7524 7840 8217 7868
rect 7524 7828 7530 7840
rect 8205 7837 8217 7840
rect 8251 7837 8263 7871
rect 8205 7831 8263 7837
rect 9125 7871 9183 7877
rect 9125 7837 9137 7871
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 5994 7760 6000 7812
rect 6052 7800 6058 7812
rect 6150 7803 6208 7809
rect 6150 7800 6162 7803
rect 6052 7772 6162 7800
rect 6052 7760 6058 7772
rect 6150 7769 6162 7772
rect 6196 7769 6208 7803
rect 6150 7763 6208 7769
rect 7745 7803 7803 7809
rect 7745 7769 7757 7803
rect 7791 7800 7803 7803
rect 8018 7800 8024 7812
rect 7791 7772 8024 7800
rect 7791 7769 7803 7772
rect 7745 7763 7803 7769
rect 8018 7760 8024 7772
rect 8076 7760 8082 7812
rect 9140 7800 9168 7831
rect 9214 7828 9220 7880
rect 9272 7877 9278 7880
rect 9272 7871 9321 7877
rect 9272 7837 9275 7871
rect 9309 7837 9321 7871
rect 9490 7868 9496 7880
rect 9451 7840 9496 7868
rect 9272 7831 9321 7837
rect 9272 7828 9278 7831
rect 9490 7828 9496 7840
rect 9548 7828 9554 7880
rect 9674 7828 9680 7880
rect 9732 7868 9738 7880
rect 10060 7868 10088 7976
rect 13541 7973 13553 8007
rect 13587 8004 13599 8007
rect 15102 8004 15108 8016
rect 13587 7976 15108 8004
rect 13587 7973 13599 7976
rect 13541 7967 13599 7973
rect 15102 7964 15108 7976
rect 15160 7964 15166 8016
rect 16960 8004 16988 8044
rect 17126 8032 17132 8044
rect 17184 8032 17190 8084
rect 17678 8072 17684 8084
rect 17639 8044 17684 8072
rect 17678 8032 17684 8044
rect 17736 8032 17742 8084
rect 19429 8075 19487 8081
rect 19429 8041 19441 8075
rect 19475 8072 19487 8075
rect 20070 8072 20076 8084
rect 19475 8044 20076 8072
rect 19475 8041 19487 8044
rect 19429 8035 19487 8041
rect 20070 8032 20076 8044
rect 20128 8032 20134 8084
rect 27154 8032 27160 8084
rect 27212 8072 27218 8084
rect 27985 8075 28043 8081
rect 27212 8044 27844 8072
rect 27212 8032 27218 8044
rect 20625 8007 20683 8013
rect 20625 8004 20637 8007
rect 16960 7976 20637 8004
rect 20625 7973 20637 7976
rect 20671 7973 20683 8007
rect 20625 7967 20683 7973
rect 10594 7936 10600 7948
rect 10555 7908 10600 7936
rect 10594 7896 10600 7908
rect 10652 7896 10658 7948
rect 12989 7939 13047 7945
rect 12989 7905 13001 7939
rect 13035 7936 13047 7939
rect 14458 7936 14464 7948
rect 13035 7908 14464 7936
rect 13035 7905 13047 7908
rect 12989 7899 13047 7905
rect 14458 7896 14464 7908
rect 14516 7896 14522 7948
rect 17126 7896 17132 7948
rect 17184 7936 17190 7948
rect 17184 7908 18368 7936
rect 17184 7896 17190 7908
rect 10505 7871 10563 7877
rect 10505 7868 10517 7871
rect 9732 7840 9777 7868
rect 10060 7840 10517 7868
rect 9732 7828 9738 7840
rect 10505 7837 10517 7840
rect 10551 7837 10563 7871
rect 10505 7831 10563 7837
rect 11885 7871 11943 7877
rect 11885 7837 11897 7871
rect 11931 7868 11943 7871
rect 13354 7868 13360 7880
rect 11931 7840 13360 7868
rect 11931 7837 11943 7840
rect 11885 7831 11943 7837
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 14093 7871 14151 7877
rect 14093 7837 14105 7871
rect 14139 7868 14151 7871
rect 14274 7868 14280 7880
rect 14139 7840 14280 7868
rect 14139 7837 14151 7840
rect 14093 7831 14151 7837
rect 14274 7828 14280 7840
rect 14332 7868 14338 7880
rect 14734 7868 14740 7880
rect 14332 7840 14740 7868
rect 14332 7828 14338 7840
rect 14734 7828 14740 7840
rect 14792 7828 14798 7880
rect 14829 7871 14887 7877
rect 14829 7837 14841 7871
rect 14875 7868 14887 7871
rect 14875 7840 15516 7868
rect 14875 7837 14887 7840
rect 14829 7831 14887 7837
rect 10042 7800 10048 7812
rect 9140 7772 10048 7800
rect 10042 7760 10048 7772
rect 10100 7760 10106 7812
rect 12437 7803 12495 7809
rect 12437 7769 12449 7803
rect 12483 7800 12495 7803
rect 13906 7800 13912 7812
rect 12483 7772 13912 7800
rect 12483 7769 12495 7772
rect 12437 7763 12495 7769
rect 13906 7760 13912 7772
rect 13964 7760 13970 7812
rect 15488 7744 15516 7840
rect 17862 7828 17868 7880
rect 17920 7868 17926 7880
rect 17957 7871 18015 7877
rect 17957 7868 17969 7871
rect 17920 7840 17969 7868
rect 17920 7828 17926 7840
rect 17957 7837 17969 7840
rect 18003 7837 18015 7871
rect 17957 7831 18015 7837
rect 18049 7871 18107 7877
rect 18049 7837 18061 7871
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 18064 7800 18092 7831
rect 18138 7828 18144 7880
rect 18196 7868 18202 7880
rect 18340 7877 18368 7908
rect 18325 7871 18383 7877
rect 18196 7840 18241 7868
rect 18196 7828 18202 7840
rect 18325 7837 18337 7871
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 19058 7828 19064 7880
rect 19116 7868 19122 7880
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 19116 7840 19257 7868
rect 19116 7828 19122 7840
rect 19245 7837 19257 7840
rect 19291 7837 19303 7871
rect 20640 7868 20668 7967
rect 25958 7964 25964 8016
rect 26016 8004 26022 8016
rect 26237 8007 26295 8013
rect 26237 8004 26249 8007
rect 26016 7976 26249 8004
rect 26016 7964 26022 7976
rect 26237 7973 26249 7976
rect 26283 8004 26295 8007
rect 27816 8004 27844 8044
rect 27985 8041 27997 8075
rect 28031 8072 28043 8075
rect 28718 8072 28724 8084
rect 28031 8044 28724 8072
rect 28031 8041 28043 8044
rect 27985 8035 28043 8041
rect 28718 8032 28724 8044
rect 28776 8032 28782 8084
rect 35069 8007 35127 8013
rect 35069 8004 35081 8007
rect 26283 7976 27752 8004
rect 27816 7976 35081 8004
rect 26283 7973 26295 7976
rect 26237 7967 26295 7973
rect 20714 7896 20720 7948
rect 20772 7936 20778 7948
rect 20772 7908 22324 7936
rect 20772 7896 20778 7908
rect 20806 7868 20812 7880
rect 20640 7840 20812 7868
rect 19245 7831 19303 7837
rect 20806 7828 20812 7840
rect 20864 7868 20870 7880
rect 21177 7871 21235 7877
rect 21177 7868 21189 7871
rect 20864 7840 21189 7868
rect 20864 7828 20870 7840
rect 21177 7837 21189 7840
rect 21223 7837 21235 7871
rect 21177 7831 21235 7837
rect 21361 7871 21419 7877
rect 21361 7837 21373 7871
rect 21407 7868 21419 7871
rect 22094 7868 22100 7880
rect 21407 7840 22100 7868
rect 21407 7837 21419 7840
rect 21361 7831 21419 7837
rect 22094 7828 22100 7840
rect 22152 7828 22158 7880
rect 18230 7800 18236 7812
rect 18064 7772 18236 7800
rect 18230 7760 18236 7772
rect 18288 7800 18294 7812
rect 18690 7800 18696 7812
rect 18288 7772 18696 7800
rect 18288 7760 18294 7772
rect 18690 7760 18696 7772
rect 18748 7760 18754 7812
rect 22296 7800 22324 7908
rect 23037 7871 23095 7877
rect 23037 7837 23049 7871
rect 23083 7868 23095 7871
rect 23198 7868 23204 7880
rect 23083 7840 23204 7868
rect 23083 7837 23095 7840
rect 23037 7831 23095 7837
rect 23198 7828 23204 7840
rect 23256 7828 23262 7880
rect 23293 7871 23351 7877
rect 23293 7837 23305 7871
rect 23339 7868 23351 7871
rect 24857 7871 24915 7877
rect 24857 7868 24869 7871
rect 23339 7840 24869 7868
rect 23339 7837 23351 7840
rect 23293 7831 23351 7837
rect 24857 7837 24869 7840
rect 24903 7868 24915 7871
rect 24946 7868 24952 7880
rect 24903 7840 24952 7868
rect 24903 7837 24915 7840
rect 24857 7831 24915 7837
rect 24946 7828 24952 7840
rect 25004 7828 25010 7880
rect 27724 7877 27752 7976
rect 35069 7973 35081 7976
rect 35115 7973 35127 8007
rect 35069 7967 35127 7973
rect 35342 7936 35348 7948
rect 35268 7908 35348 7936
rect 27433 7871 27491 7877
rect 27433 7868 27445 7871
rect 25056 7840 27445 7868
rect 25056 7800 25084 7840
rect 27433 7837 27445 7840
rect 27479 7837 27491 7871
rect 27433 7831 27491 7837
rect 27709 7871 27767 7877
rect 27709 7837 27721 7871
rect 27755 7837 27767 7871
rect 27709 7831 27767 7837
rect 27798 7828 27804 7880
rect 27856 7868 27862 7880
rect 30837 7871 30895 7877
rect 27856 7840 27901 7868
rect 27856 7828 27862 7840
rect 30837 7837 30849 7871
rect 30883 7868 30895 7871
rect 31662 7868 31668 7880
rect 30883 7840 31668 7868
rect 30883 7837 30895 7840
rect 30837 7831 30895 7837
rect 31662 7828 31668 7840
rect 31720 7828 31726 7880
rect 35268 7877 35296 7908
rect 35342 7896 35348 7908
rect 35400 7896 35406 7948
rect 35253 7871 35311 7877
rect 35253 7837 35265 7871
rect 35299 7837 35311 7871
rect 35253 7831 35311 7837
rect 35437 7871 35495 7877
rect 35437 7837 35449 7871
rect 35483 7868 35495 7871
rect 35526 7868 35532 7880
rect 35483 7840 35532 7868
rect 35483 7837 35495 7840
rect 35437 7831 35495 7837
rect 35526 7828 35532 7840
rect 35584 7828 35590 7880
rect 35618 7828 35624 7880
rect 35676 7868 35682 7880
rect 58158 7868 58164 7880
rect 35676 7840 35721 7868
rect 58119 7840 58164 7868
rect 35676 7828 35682 7840
rect 58158 7828 58164 7840
rect 58216 7828 58222 7880
rect 22296 7772 25084 7800
rect 25124 7803 25182 7809
rect 25124 7769 25136 7803
rect 25170 7800 25182 7803
rect 25314 7800 25320 7812
rect 25170 7772 25320 7800
rect 25170 7769 25182 7772
rect 25124 7763 25182 7769
rect 25314 7760 25320 7772
rect 25372 7760 25378 7812
rect 27617 7803 27675 7809
rect 27617 7769 27629 7803
rect 27663 7800 27675 7803
rect 28258 7800 28264 7812
rect 27663 7772 28264 7800
rect 27663 7769 27675 7772
rect 27617 7763 27675 7769
rect 28258 7760 28264 7772
rect 28316 7760 28322 7812
rect 31021 7803 31079 7809
rect 31021 7769 31033 7803
rect 31067 7800 31079 7803
rect 31478 7800 31484 7812
rect 31067 7772 31484 7800
rect 31067 7769 31079 7772
rect 31021 7763 31079 7769
rect 31478 7760 31484 7772
rect 31536 7760 31542 7812
rect 35345 7803 35403 7809
rect 35345 7769 35357 7803
rect 35391 7800 35403 7803
rect 37182 7800 37188 7812
rect 35391 7772 37188 7800
rect 35391 7769 35403 7772
rect 35345 7763 35403 7769
rect 37182 7760 37188 7772
rect 37240 7760 37246 7812
rect 1486 7732 1492 7744
rect 1447 7704 1492 7732
rect 1486 7692 1492 7704
rect 1544 7692 1550 7744
rect 2498 7732 2504 7744
rect 2459 7704 2504 7732
rect 2498 7692 2504 7704
rect 2556 7692 2562 7744
rect 2961 7735 3019 7741
rect 2961 7701 2973 7735
rect 3007 7732 3019 7735
rect 3786 7732 3792 7744
rect 3007 7704 3792 7732
rect 3007 7701 3019 7704
rect 2961 7695 3019 7701
rect 3786 7692 3792 7704
rect 3844 7692 3850 7744
rect 3970 7732 3976 7744
rect 3931 7704 3976 7732
rect 3970 7692 3976 7704
rect 4028 7692 4034 7744
rect 4706 7732 4712 7744
rect 4667 7704 4712 7732
rect 4706 7692 4712 7704
rect 4764 7692 4770 7744
rect 5166 7692 5172 7744
rect 5224 7692 5230 7744
rect 8938 7692 8944 7744
rect 8996 7732 9002 7744
rect 8996 7704 9041 7732
rect 8996 7692 9002 7704
rect 9490 7692 9496 7744
rect 9548 7732 9554 7744
rect 10137 7735 10195 7741
rect 10137 7732 10149 7735
rect 9548 7704 10149 7732
rect 9548 7692 9554 7704
rect 10137 7701 10149 7704
rect 10183 7732 10195 7735
rect 10778 7732 10784 7744
rect 10183 7704 10784 7732
rect 10183 7701 10195 7704
rect 10137 7695 10195 7701
rect 10778 7692 10784 7704
rect 10836 7692 10842 7744
rect 11333 7735 11391 7741
rect 11333 7701 11345 7735
rect 11379 7732 11391 7735
rect 12066 7732 12072 7744
rect 11379 7704 12072 7732
rect 11379 7701 11391 7704
rect 11333 7695 11391 7701
rect 12066 7692 12072 7704
rect 12124 7692 12130 7744
rect 14918 7692 14924 7744
rect 14976 7732 14982 7744
rect 15013 7735 15071 7741
rect 15013 7732 15025 7735
rect 14976 7704 15025 7732
rect 14976 7692 14982 7704
rect 15013 7701 15025 7704
rect 15059 7701 15071 7735
rect 15013 7695 15071 7701
rect 15470 7692 15476 7744
rect 15528 7732 15534 7744
rect 15565 7735 15623 7741
rect 15565 7732 15577 7735
rect 15528 7704 15577 7732
rect 15528 7692 15534 7704
rect 15565 7701 15577 7704
rect 15611 7701 15623 7735
rect 16666 7732 16672 7744
rect 16627 7704 16672 7732
rect 15565 7695 15623 7701
rect 16666 7692 16672 7704
rect 16724 7692 16730 7744
rect 21266 7732 21272 7744
rect 21227 7704 21272 7732
rect 21266 7692 21272 7704
rect 21324 7692 21330 7744
rect 21913 7735 21971 7741
rect 21913 7701 21925 7735
rect 21959 7732 21971 7735
rect 22554 7732 22560 7744
rect 21959 7704 22560 7732
rect 21959 7701 21971 7704
rect 21913 7695 21971 7701
rect 22554 7692 22560 7704
rect 22612 7692 22618 7744
rect 24670 7692 24676 7744
rect 24728 7732 24734 7744
rect 26878 7732 26884 7744
rect 24728 7704 26884 7732
rect 24728 7692 24734 7704
rect 26878 7692 26884 7704
rect 26936 7692 26942 7744
rect 30650 7732 30656 7744
rect 30611 7704 30656 7732
rect 30650 7692 30656 7704
rect 30708 7692 30714 7744
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 3053 7531 3111 7537
rect 3053 7528 3065 7531
rect 2746 7500 3065 7528
rect 2222 7392 2228 7404
rect 2183 7364 2228 7392
rect 2222 7352 2228 7364
rect 2280 7352 2286 7404
rect 2409 7395 2467 7401
rect 2409 7361 2421 7395
rect 2455 7392 2467 7395
rect 2746 7392 2774 7500
rect 3053 7497 3065 7500
rect 3099 7497 3111 7531
rect 3510 7528 3516 7540
rect 3471 7500 3516 7528
rect 3053 7491 3111 7497
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 5166 7528 5172 7540
rect 5127 7500 5172 7528
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 7926 7528 7932 7540
rect 7887 7500 7932 7528
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 8018 7488 8024 7540
rect 8076 7528 8082 7540
rect 9490 7528 9496 7540
rect 8076 7500 9496 7528
rect 8076 7488 8082 7500
rect 9490 7488 9496 7500
rect 9548 7488 9554 7540
rect 10134 7488 10140 7540
rect 10192 7528 10198 7540
rect 10318 7528 10324 7540
rect 10192 7500 10324 7528
rect 10192 7488 10198 7500
rect 10318 7488 10324 7500
rect 10376 7528 10382 7540
rect 10873 7531 10931 7537
rect 10873 7528 10885 7531
rect 10376 7500 10885 7528
rect 10376 7488 10382 7500
rect 10873 7497 10885 7500
rect 10919 7497 10931 7531
rect 10873 7491 10931 7497
rect 14461 7531 14519 7537
rect 14461 7497 14473 7531
rect 14507 7528 14519 7531
rect 14550 7528 14556 7540
rect 14507 7500 14556 7528
rect 14507 7497 14519 7500
rect 14461 7491 14519 7497
rect 14550 7488 14556 7500
rect 14608 7488 14614 7540
rect 15010 7528 15016 7540
rect 14971 7500 15016 7528
rect 15010 7488 15016 7500
rect 15068 7488 15074 7540
rect 17589 7531 17647 7537
rect 17589 7528 17601 7531
rect 15120 7500 17601 7528
rect 3421 7463 3479 7469
rect 3421 7429 3433 7463
rect 3467 7460 3479 7463
rect 3970 7460 3976 7472
rect 3467 7432 3976 7460
rect 3467 7429 3479 7432
rect 3421 7423 3479 7429
rect 3970 7420 3976 7432
rect 4028 7420 4034 7472
rect 4525 7463 4583 7469
rect 4525 7429 4537 7463
rect 4571 7460 4583 7463
rect 5534 7460 5540 7472
rect 4571 7432 5540 7460
rect 4571 7429 4583 7432
rect 4525 7423 4583 7429
rect 5534 7420 5540 7432
rect 5592 7420 5598 7472
rect 5644 7432 9536 7460
rect 2455 7364 2774 7392
rect 2455 7361 2467 7364
rect 2409 7355 2467 7361
rect 3786 7352 3792 7404
rect 3844 7392 3850 7404
rect 4893 7395 4951 7401
rect 4893 7392 4905 7395
rect 3844 7364 4905 7392
rect 3844 7352 3850 7364
rect 4893 7361 4905 7364
rect 4939 7361 4951 7395
rect 4893 7355 4951 7361
rect 4985 7395 5043 7401
rect 4985 7361 4997 7395
rect 5031 7392 5043 7395
rect 5074 7392 5080 7404
rect 5031 7364 5080 7392
rect 5031 7361 5043 7364
rect 4985 7355 5043 7361
rect 5074 7352 5080 7364
rect 5132 7352 5138 7404
rect 3694 7324 3700 7336
rect 3655 7296 3700 7324
rect 3694 7284 3700 7296
rect 3752 7284 3758 7336
rect 3878 7284 3884 7336
rect 3936 7324 3942 7336
rect 5644 7324 5672 7432
rect 9508 7404 9536 7432
rect 12710 7420 12716 7472
rect 12768 7469 12774 7472
rect 12768 7460 12780 7469
rect 15120 7460 15148 7500
rect 17589 7497 17601 7500
rect 17635 7528 17647 7531
rect 17862 7528 17868 7540
rect 17635 7500 17868 7528
rect 17635 7497 17647 7500
rect 17589 7491 17647 7497
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 22833 7531 22891 7537
rect 22833 7497 22845 7531
rect 22879 7528 22891 7531
rect 23106 7528 23112 7540
rect 22879 7500 23112 7528
rect 22879 7497 22891 7500
rect 22833 7491 22891 7497
rect 23106 7488 23112 7500
rect 23164 7488 23170 7540
rect 23290 7528 23296 7540
rect 23251 7500 23296 7528
rect 23290 7488 23296 7500
rect 23348 7488 23354 7540
rect 31573 7531 31631 7537
rect 24872 7500 25268 7528
rect 16669 7463 16727 7469
rect 16669 7460 16681 7463
rect 12768 7432 12813 7460
rect 14016 7432 15148 7460
rect 15488 7432 16681 7460
rect 12768 7423 12780 7432
rect 12768 7420 12774 7423
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 7837 7395 7895 7401
rect 6871 7364 7512 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 7009 7327 7067 7333
rect 7009 7324 7021 7327
rect 3936 7296 5672 7324
rect 5736 7296 7021 7324
rect 3936 7284 3942 7296
rect 1765 7259 1823 7265
rect 1765 7225 1777 7259
rect 1811 7256 1823 7259
rect 3142 7256 3148 7268
rect 1811 7228 3148 7256
rect 1811 7225 1823 7228
rect 1765 7219 1823 7225
rect 3142 7216 3148 7228
rect 3200 7216 3206 7268
rect 5736 7200 5764 7296
rect 7009 7293 7021 7296
rect 7055 7324 7067 7327
rect 7098 7324 7104 7336
rect 7055 7296 7104 7324
rect 7055 7293 7067 7296
rect 7009 7287 7067 7293
rect 7098 7284 7104 7296
rect 7156 7284 7162 7336
rect 7484 7265 7512 7364
rect 7837 7361 7849 7395
rect 7883 7361 7895 7395
rect 7837 7355 7895 7361
rect 7469 7259 7527 7265
rect 7469 7225 7481 7259
rect 7515 7225 7527 7259
rect 7469 7219 7527 7225
rect 2593 7191 2651 7197
rect 2593 7157 2605 7191
rect 2639 7188 2651 7191
rect 2958 7188 2964 7200
rect 2639 7160 2964 7188
rect 2639 7157 2651 7160
rect 2593 7151 2651 7157
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 5718 7188 5724 7200
rect 5679 7160 5724 7188
rect 5718 7148 5724 7160
rect 5776 7148 5782 7200
rect 6178 7148 6184 7200
rect 6236 7188 6242 7200
rect 6641 7191 6699 7197
rect 6641 7188 6653 7191
rect 6236 7160 6653 7188
rect 6236 7148 6242 7160
rect 6641 7157 6653 7160
rect 6687 7157 6699 7191
rect 7852 7188 7880 7355
rect 9490 7352 9496 7404
rect 9548 7392 9554 7404
rect 14016 7392 14044 7432
rect 14274 7392 14280 7404
rect 9548 7364 14044 7392
rect 14235 7364 14280 7392
rect 9548 7352 9554 7364
rect 14274 7352 14280 7364
rect 14332 7352 14338 7404
rect 15286 7392 15292 7404
rect 15247 7364 15292 7392
rect 15286 7352 15292 7364
rect 15344 7352 15350 7404
rect 15488 7401 15516 7432
rect 16669 7429 16681 7432
rect 16715 7429 16727 7463
rect 16669 7423 16727 7429
rect 16850 7420 16856 7472
rect 16908 7460 16914 7472
rect 22554 7460 22560 7472
rect 16908 7432 22094 7460
rect 22515 7432 22560 7460
rect 16908 7420 16914 7432
rect 15381 7395 15439 7401
rect 15381 7361 15393 7395
rect 15427 7361 15439 7395
rect 15381 7355 15439 7361
rect 15473 7395 15531 7401
rect 15473 7361 15485 7395
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 15657 7395 15715 7401
rect 15657 7361 15669 7395
rect 15703 7392 15715 7395
rect 16942 7392 16948 7404
rect 15703 7364 16948 7392
rect 15703 7361 15715 7364
rect 15657 7355 15715 7361
rect 8113 7327 8171 7333
rect 8113 7293 8125 7327
rect 8159 7324 8171 7327
rect 8202 7324 8208 7336
rect 8159 7296 8208 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 12989 7327 13047 7333
rect 12989 7293 13001 7327
rect 13035 7324 13047 7327
rect 13814 7324 13820 7336
rect 13035 7296 13820 7324
rect 13035 7293 13047 7296
rect 12989 7287 13047 7293
rect 13814 7284 13820 7296
rect 13872 7324 13878 7336
rect 14826 7324 14832 7336
rect 13872 7296 14832 7324
rect 13872 7284 13878 7296
rect 14826 7284 14832 7296
rect 14884 7284 14890 7336
rect 15396 7268 15424 7355
rect 16942 7352 16948 7364
rect 17000 7352 17006 7404
rect 17034 7352 17040 7404
rect 17092 7392 17098 7404
rect 18877 7395 18935 7401
rect 17092 7364 17137 7392
rect 17092 7352 17098 7364
rect 18877 7361 18889 7395
rect 18923 7392 18935 7395
rect 19334 7392 19340 7404
rect 18923 7364 19340 7392
rect 18923 7361 18935 7364
rect 18877 7355 18935 7361
rect 19334 7352 19340 7364
rect 19392 7352 19398 7404
rect 21085 7395 21143 7401
rect 21085 7361 21097 7395
rect 21131 7361 21143 7395
rect 21085 7355 21143 7361
rect 21269 7395 21327 7401
rect 21269 7361 21281 7395
rect 21315 7392 21327 7395
rect 21358 7392 21364 7404
rect 21315 7364 21364 7392
rect 21315 7361 21327 7364
rect 21269 7355 21327 7361
rect 20349 7327 20407 7333
rect 20349 7324 20361 7327
rect 16960 7296 20361 7324
rect 15378 7216 15384 7268
rect 15436 7216 15442 7268
rect 8202 7188 8208 7200
rect 7852 7160 8208 7188
rect 6641 7151 6699 7157
rect 8202 7148 8208 7160
rect 8260 7188 8266 7200
rect 8665 7191 8723 7197
rect 8665 7188 8677 7191
rect 8260 7160 8677 7188
rect 8260 7148 8266 7160
rect 8665 7157 8677 7160
rect 8711 7188 8723 7191
rect 8754 7188 8760 7200
rect 8711 7160 8760 7188
rect 8711 7157 8723 7160
rect 8665 7151 8723 7157
rect 8754 7148 8760 7160
rect 8812 7148 8818 7200
rect 9214 7188 9220 7200
rect 9175 7160 9220 7188
rect 9214 7148 9220 7160
rect 9272 7148 9278 7200
rect 9766 7188 9772 7200
rect 9727 7160 9772 7188
rect 9766 7148 9772 7160
rect 9824 7148 9830 7200
rect 10410 7188 10416 7200
rect 10371 7160 10416 7188
rect 10410 7148 10416 7160
rect 10468 7148 10474 7200
rect 11238 7148 11244 7200
rect 11296 7188 11302 7200
rect 11609 7191 11667 7197
rect 11609 7188 11621 7191
rect 11296 7160 11621 7188
rect 11296 7148 11302 7160
rect 11609 7157 11621 7160
rect 11655 7157 11667 7191
rect 11609 7151 11667 7157
rect 13817 7191 13875 7197
rect 13817 7157 13829 7191
rect 13863 7188 13875 7191
rect 14274 7188 14280 7200
rect 13863 7160 14280 7188
rect 13863 7157 13875 7160
rect 13817 7151 13875 7157
rect 14274 7148 14280 7160
rect 14332 7148 14338 7200
rect 14550 7148 14556 7200
rect 14608 7188 14614 7200
rect 16960 7188 16988 7296
rect 20349 7293 20361 7296
rect 20395 7324 20407 7327
rect 20901 7327 20959 7333
rect 20901 7324 20913 7327
rect 20395 7296 20913 7324
rect 20395 7293 20407 7296
rect 20349 7287 20407 7293
rect 20901 7293 20913 7296
rect 20947 7293 20959 7327
rect 21100 7324 21128 7355
rect 21358 7352 21364 7364
rect 21416 7352 21422 7404
rect 22066 7392 22094 7432
rect 22554 7420 22560 7432
rect 22612 7460 22618 7472
rect 23477 7463 23535 7469
rect 23477 7460 23489 7463
rect 22612 7432 23489 7460
rect 22612 7420 22618 7432
rect 23477 7429 23489 7432
rect 23523 7429 23535 7463
rect 23658 7460 23664 7472
rect 23619 7432 23664 7460
rect 23477 7423 23535 7429
rect 23658 7420 23664 7432
rect 23716 7420 23722 7472
rect 22281 7395 22339 7401
rect 22281 7392 22293 7395
rect 22066 7364 22293 7392
rect 22281 7361 22293 7364
rect 22327 7361 22339 7395
rect 22281 7355 22339 7361
rect 22465 7395 22523 7401
rect 22465 7361 22477 7395
rect 22511 7361 22523 7395
rect 22646 7392 22652 7404
rect 22607 7364 22652 7392
rect 22465 7355 22523 7361
rect 22094 7324 22100 7336
rect 21100 7296 22100 7324
rect 20901 7287 20959 7293
rect 22094 7284 22100 7296
rect 22152 7324 22158 7336
rect 22480 7324 22508 7355
rect 22646 7352 22652 7364
rect 22704 7392 22710 7404
rect 23382 7392 23388 7404
rect 22704 7364 23388 7392
rect 22704 7352 22710 7364
rect 23382 7352 23388 7364
rect 23440 7352 23446 7404
rect 24026 7352 24032 7404
rect 24084 7392 24090 7404
rect 24673 7395 24731 7401
rect 24673 7392 24685 7395
rect 24084 7364 24685 7392
rect 24084 7352 24090 7364
rect 24673 7361 24685 7364
rect 24719 7392 24731 7395
rect 24762 7392 24768 7404
rect 24719 7364 24768 7392
rect 24719 7361 24731 7364
rect 24673 7355 24731 7361
rect 24762 7352 24768 7364
rect 24820 7352 24826 7404
rect 24872 7401 24900 7500
rect 25240 7460 25268 7500
rect 31573 7497 31585 7531
rect 31619 7528 31631 7531
rect 31662 7528 31668 7540
rect 31619 7500 31668 7528
rect 31619 7497 31631 7500
rect 31573 7491 31631 7497
rect 31662 7488 31668 7500
rect 31720 7488 31726 7540
rect 34606 7488 34612 7540
rect 34664 7528 34670 7540
rect 35069 7531 35127 7537
rect 35069 7528 35081 7531
rect 34664 7500 35081 7528
rect 34664 7488 34670 7500
rect 35069 7497 35081 7500
rect 35115 7497 35127 7531
rect 35618 7528 35624 7540
rect 35069 7491 35127 7497
rect 35176 7500 35624 7528
rect 26145 7463 26203 7469
rect 26145 7460 26157 7463
rect 25240 7432 26157 7460
rect 26145 7429 26157 7432
rect 26191 7429 26203 7463
rect 26145 7423 26203 7429
rect 34425 7463 34483 7469
rect 34425 7429 34437 7463
rect 34471 7460 34483 7463
rect 34698 7460 34704 7472
rect 34471 7432 34704 7460
rect 34471 7429 34483 7432
rect 34425 7423 34483 7429
rect 34698 7420 34704 7432
rect 34756 7460 34762 7472
rect 35176 7460 35204 7500
rect 35618 7488 35624 7500
rect 35676 7488 35682 7540
rect 36357 7531 36415 7537
rect 36357 7497 36369 7531
rect 36403 7528 36415 7531
rect 36630 7528 36636 7540
rect 36403 7500 36636 7528
rect 36403 7497 36415 7500
rect 36357 7491 36415 7497
rect 36630 7488 36636 7500
rect 36688 7528 36694 7540
rect 37090 7528 37096 7540
rect 36688 7500 37096 7528
rect 36688 7488 36694 7500
rect 37090 7488 37096 7500
rect 37148 7528 37154 7540
rect 38013 7531 38071 7537
rect 38013 7528 38025 7531
rect 37148 7500 38025 7528
rect 37148 7488 37154 7500
rect 38013 7497 38025 7500
rect 38059 7528 38071 7531
rect 39022 7528 39028 7540
rect 38059 7500 39028 7528
rect 38059 7497 38071 7500
rect 38013 7491 38071 7497
rect 39022 7488 39028 7500
rect 39080 7488 39086 7540
rect 34756 7432 35204 7460
rect 35437 7463 35495 7469
rect 34756 7420 34762 7432
rect 35437 7429 35449 7463
rect 35483 7460 35495 7463
rect 35526 7460 35532 7472
rect 35483 7432 35532 7460
rect 35483 7429 35495 7432
rect 35437 7423 35495 7429
rect 35526 7420 35532 7432
rect 35584 7420 35590 7472
rect 24857 7395 24915 7401
rect 24857 7361 24869 7395
rect 24903 7361 24915 7395
rect 24857 7355 24915 7361
rect 24949 7395 25007 7401
rect 24949 7361 24961 7395
rect 24995 7361 25007 7395
rect 24949 7355 25007 7361
rect 25041 7395 25099 7401
rect 25041 7361 25053 7395
rect 25087 7361 25099 7395
rect 25774 7392 25780 7404
rect 25735 7364 25780 7392
rect 25041 7355 25099 7361
rect 22738 7324 22744 7336
rect 22152 7296 22744 7324
rect 22152 7284 22158 7296
rect 22738 7284 22744 7296
rect 22796 7284 22802 7336
rect 23934 7284 23940 7336
rect 23992 7324 23998 7336
rect 24302 7324 24308 7336
rect 23992 7296 24308 7324
rect 23992 7284 23998 7296
rect 24302 7284 24308 7296
rect 24360 7324 24366 7336
rect 24964 7324 24992 7355
rect 24360 7296 24992 7324
rect 25056 7324 25084 7355
rect 25774 7352 25780 7364
rect 25832 7352 25838 7404
rect 25958 7392 25964 7404
rect 25919 7364 25964 7392
rect 25958 7352 25964 7364
rect 26016 7352 26022 7404
rect 26878 7352 26884 7404
rect 26936 7392 26942 7404
rect 27617 7395 27675 7401
rect 27617 7392 27629 7395
rect 26936 7364 27629 7392
rect 26936 7352 26942 7364
rect 27617 7361 27629 7364
rect 27663 7361 27675 7395
rect 27617 7355 27675 7361
rect 27706 7395 27764 7401
rect 27706 7361 27718 7395
rect 27752 7361 27764 7395
rect 27706 7355 27764 7361
rect 25314 7324 25320 7336
rect 25056 7296 25167 7324
rect 25275 7296 25320 7324
rect 24360 7284 24366 7296
rect 17034 7216 17040 7268
rect 17092 7256 17098 7268
rect 18693 7259 18751 7265
rect 18693 7256 18705 7259
rect 17092 7228 18705 7256
rect 17092 7216 17098 7228
rect 18693 7225 18705 7228
rect 18739 7256 18751 7259
rect 18782 7256 18788 7268
rect 18739 7228 18788 7256
rect 18739 7225 18751 7228
rect 18693 7219 18751 7225
rect 18782 7216 18788 7228
rect 18840 7216 18846 7268
rect 20070 7216 20076 7268
rect 20128 7256 20134 7268
rect 24121 7259 24179 7265
rect 24121 7256 24133 7259
rect 20128 7228 24133 7256
rect 20128 7216 20134 7228
rect 24121 7225 24133 7228
rect 24167 7225 24179 7259
rect 24121 7219 24179 7225
rect 25139 7256 25167 7296
rect 25314 7284 25320 7296
rect 25372 7284 25378 7336
rect 26234 7284 26240 7336
rect 26292 7324 26298 7336
rect 27721 7324 27749 7355
rect 27798 7352 27804 7404
rect 27856 7401 27862 7404
rect 27856 7392 27864 7401
rect 27856 7364 27901 7392
rect 27856 7355 27864 7364
rect 27856 7352 27862 7355
rect 27982 7352 27988 7404
rect 28040 7392 28046 7404
rect 28040 7364 28085 7392
rect 28040 7352 28046 7364
rect 28166 7352 28172 7404
rect 28224 7392 28230 7404
rect 30466 7401 30472 7404
rect 28445 7395 28503 7401
rect 28445 7392 28457 7395
rect 28224 7364 28457 7392
rect 28224 7352 28230 7364
rect 28445 7361 28457 7364
rect 28491 7361 28503 7395
rect 28445 7355 28503 7361
rect 30460 7355 30472 7401
rect 30524 7392 30530 7404
rect 34609 7395 34667 7401
rect 30524 7364 30560 7392
rect 30466 7352 30472 7355
rect 30524 7352 30530 7364
rect 34609 7361 34621 7395
rect 34655 7392 34667 7395
rect 34790 7392 34796 7404
rect 34655 7364 34796 7392
rect 34655 7361 34667 7364
rect 34609 7355 34667 7361
rect 34790 7352 34796 7364
rect 34848 7352 34854 7404
rect 35250 7392 35256 7404
rect 35211 7364 35256 7392
rect 35250 7352 35256 7364
rect 35308 7352 35314 7404
rect 35345 7395 35403 7401
rect 35345 7361 35357 7395
rect 35391 7361 35403 7395
rect 35345 7355 35403 7361
rect 35621 7395 35679 7401
rect 35621 7361 35633 7395
rect 35667 7392 35679 7395
rect 36170 7392 36176 7404
rect 35667 7364 36176 7392
rect 35667 7361 35679 7364
rect 35621 7355 35679 7361
rect 26292 7296 27749 7324
rect 26292 7284 26298 7296
rect 29822 7284 29828 7336
rect 29880 7324 29886 7336
rect 30193 7327 30251 7333
rect 30193 7324 30205 7327
rect 29880 7296 30205 7324
rect 29880 7284 29886 7296
rect 30193 7293 30205 7296
rect 30239 7293 30251 7327
rect 35360 7324 35388 7355
rect 36170 7352 36176 7364
rect 36228 7352 36234 7404
rect 37642 7352 37648 7404
rect 37700 7392 37706 7404
rect 38565 7395 38623 7401
rect 38565 7392 38577 7395
rect 37700 7364 38577 7392
rect 37700 7352 37706 7364
rect 38565 7361 38577 7364
rect 38611 7361 38623 7395
rect 38565 7355 38623 7361
rect 38749 7395 38807 7401
rect 38749 7361 38761 7395
rect 38795 7361 38807 7395
rect 38749 7355 38807 7361
rect 38764 7324 38792 7355
rect 39666 7324 39672 7336
rect 35360 7296 39672 7324
rect 30193 7287 30251 7293
rect 39666 7284 39672 7296
rect 39724 7284 39730 7336
rect 27614 7256 27620 7268
rect 25139 7228 27620 7256
rect 18138 7188 18144 7200
rect 14608 7160 16988 7188
rect 18099 7160 18144 7188
rect 14608 7148 14614 7160
rect 18138 7148 18144 7160
rect 18196 7188 18202 7200
rect 19058 7188 19064 7200
rect 18196 7160 19064 7188
rect 18196 7148 18202 7160
rect 19058 7148 19064 7160
rect 19116 7188 19122 7200
rect 19337 7191 19395 7197
rect 19337 7188 19349 7191
rect 19116 7160 19349 7188
rect 19116 7148 19122 7160
rect 19337 7157 19349 7160
rect 19383 7157 19395 7191
rect 24136 7188 24164 7219
rect 25139 7188 25167 7228
rect 27614 7216 27620 7228
rect 27672 7216 27678 7268
rect 34241 7259 34299 7265
rect 34241 7225 34253 7259
rect 34287 7256 34299 7259
rect 35342 7256 35348 7268
rect 34287 7228 35348 7256
rect 34287 7225 34299 7228
rect 34241 7219 34299 7225
rect 35342 7216 35348 7228
rect 35400 7216 35406 7268
rect 27338 7188 27344 7200
rect 24136 7160 25167 7188
rect 27299 7160 27344 7188
rect 19337 7151 19395 7157
rect 27338 7148 27344 7160
rect 27396 7148 27402 7200
rect 28626 7188 28632 7200
rect 28587 7160 28632 7188
rect 28626 7148 28632 7160
rect 28684 7148 28690 7200
rect 38838 7148 38844 7200
rect 38896 7188 38902 7200
rect 38933 7191 38991 7197
rect 38933 7188 38945 7191
rect 38896 7160 38945 7188
rect 38896 7148 38902 7160
rect 38933 7157 38945 7160
rect 38979 7157 38991 7191
rect 38933 7151 38991 7157
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 3602 6944 3608 6996
rect 3660 6984 3666 6996
rect 5350 6984 5356 6996
rect 3660 6956 5356 6984
rect 3660 6944 3666 6956
rect 5350 6944 5356 6956
rect 5408 6944 5414 6996
rect 5994 6984 6000 6996
rect 5955 6956 6000 6984
rect 5994 6944 6000 6956
rect 6052 6944 6058 6996
rect 3970 6876 3976 6928
rect 4028 6916 4034 6928
rect 5258 6916 5264 6928
rect 4028 6888 5264 6916
rect 4028 6876 4034 6888
rect 5258 6876 5264 6888
rect 5316 6916 5322 6928
rect 9490 6916 9496 6928
rect 5316 6888 9496 6916
rect 5316 6876 5322 6888
rect 9490 6876 9496 6888
rect 9548 6876 9554 6928
rect 14918 6876 14924 6928
rect 14976 6916 14982 6928
rect 14976 6888 18552 6916
rect 14976 6876 14982 6888
rect 3881 6851 3939 6857
rect 3881 6817 3893 6851
rect 3927 6848 3939 6851
rect 6086 6848 6092 6860
rect 3927 6820 6092 6848
rect 3927 6817 3939 6820
rect 3881 6811 3939 6817
rect 6086 6808 6092 6820
rect 6144 6808 6150 6860
rect 7374 6848 7380 6860
rect 6564 6820 7380 6848
rect 2222 6780 2228 6792
rect 2183 6752 2228 6780
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 2317 6783 2375 6789
rect 2317 6749 2329 6783
rect 2363 6780 2375 6783
rect 2498 6780 2504 6792
rect 2363 6752 2504 6780
rect 2363 6749 2375 6752
rect 2317 6743 2375 6749
rect 2498 6740 2504 6752
rect 2556 6740 2562 6792
rect 2958 6740 2964 6792
rect 3016 6780 3022 6792
rect 3145 6783 3203 6789
rect 3145 6780 3157 6783
rect 3016 6752 3157 6780
rect 3016 6740 3022 6752
rect 3145 6749 3157 6752
rect 3191 6749 3203 6783
rect 5258 6780 5264 6792
rect 3145 6743 3203 6749
rect 4356 6752 5264 6780
rect 1673 6715 1731 6721
rect 1673 6681 1685 6715
rect 1719 6712 1731 6715
rect 4356 6712 4384 6752
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 6178 6780 6184 6792
rect 6139 6752 6184 6780
rect 6178 6740 6184 6752
rect 6236 6740 6242 6792
rect 1719 6684 4384 6712
rect 4433 6715 4491 6721
rect 1719 6681 1731 6684
rect 1673 6675 1731 6681
rect 4433 6681 4445 6715
rect 4479 6712 4491 6715
rect 5810 6712 5816 6724
rect 4479 6684 5816 6712
rect 4479 6681 4491 6684
rect 4433 6675 4491 6681
rect 5810 6672 5816 6684
rect 5868 6672 5874 6724
rect 2222 6604 2228 6656
rect 2280 6644 2286 6656
rect 2501 6647 2559 6653
rect 2501 6644 2513 6647
rect 2280 6616 2513 6644
rect 2280 6604 2286 6616
rect 2501 6613 2513 6616
rect 2547 6613 2559 6647
rect 2958 6644 2964 6656
rect 2919 6616 2964 6644
rect 2501 6607 2559 6613
rect 2958 6604 2964 6616
rect 3016 6604 3022 6656
rect 4982 6644 4988 6656
rect 4943 6616 4988 6644
rect 4982 6604 4988 6616
rect 5040 6604 5046 6656
rect 5537 6647 5595 6653
rect 5537 6613 5549 6647
rect 5583 6644 5595 6647
rect 6564 6644 6592 6820
rect 7374 6808 7380 6820
rect 7432 6808 7438 6860
rect 8754 6848 8760 6860
rect 7944 6820 8760 6848
rect 6641 6783 6699 6789
rect 6641 6749 6653 6783
rect 6687 6749 6699 6783
rect 6641 6743 6699 6749
rect 7469 6783 7527 6789
rect 7469 6749 7481 6783
rect 7515 6780 7527 6783
rect 7558 6780 7564 6792
rect 7515 6752 7564 6780
rect 7515 6749 7527 6752
rect 7469 6743 7527 6749
rect 6656 6712 6684 6743
rect 7558 6740 7564 6752
rect 7616 6740 7622 6792
rect 7944 6789 7972 6820
rect 8754 6808 8760 6820
rect 8812 6808 8818 6860
rect 11885 6851 11943 6857
rect 11885 6817 11897 6851
rect 11931 6848 11943 6851
rect 13814 6848 13820 6860
rect 11931 6820 13820 6848
rect 11931 6817 11943 6820
rect 11885 6811 11943 6817
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 13998 6808 14004 6860
rect 14056 6848 14062 6860
rect 14277 6851 14335 6857
rect 14277 6848 14289 6851
rect 14056 6820 14289 6848
rect 14056 6808 14062 6820
rect 14277 6817 14289 6820
rect 14323 6817 14335 6851
rect 14277 6811 14335 6817
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 8386 6740 8392 6792
rect 8444 6780 8450 6792
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 8444 6752 9137 6780
rect 8444 6740 8450 6752
rect 9125 6749 9137 6752
rect 9171 6780 9183 6783
rect 9214 6780 9220 6792
rect 9171 6752 9220 6780
rect 9171 6749 9183 6752
rect 9125 6743 9183 6749
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 11606 6740 11612 6792
rect 11664 6789 11670 6792
rect 11664 6780 11676 6789
rect 12621 6783 12679 6789
rect 11664 6752 11709 6780
rect 11664 6743 11676 6752
rect 12621 6749 12633 6783
rect 12667 6780 12679 6783
rect 14918 6780 14924 6792
rect 12667 6752 14924 6780
rect 12667 6749 12679 6752
rect 12621 6743 12679 6749
rect 11664 6740 11670 6743
rect 14918 6740 14924 6752
rect 14976 6740 14982 6792
rect 15933 6783 15991 6789
rect 15580 6752 15884 6780
rect 8570 6712 8576 6724
rect 6656 6684 8576 6712
rect 5583 6616 6592 6644
rect 6825 6647 6883 6653
rect 5583 6613 5595 6616
rect 5537 6607 5595 6613
rect 6825 6613 6837 6647
rect 6871 6644 6883 6647
rect 7098 6644 7104 6656
rect 6871 6616 7104 6644
rect 6871 6613 6883 6616
rect 6825 6607 6883 6613
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 7300 6653 7328 6684
rect 8570 6672 8576 6684
rect 8628 6672 8634 6724
rect 10045 6715 10103 6721
rect 10045 6681 10057 6715
rect 10091 6712 10103 6715
rect 13078 6712 13084 6724
rect 10091 6684 13084 6712
rect 10091 6681 10103 6684
rect 10045 6675 10103 6681
rect 13078 6672 13084 6684
rect 13136 6672 13142 6724
rect 13541 6715 13599 6721
rect 13541 6681 13553 6715
rect 13587 6712 13599 6715
rect 15580 6712 15608 6752
rect 15746 6712 15752 6724
rect 13587 6684 15608 6712
rect 15707 6684 15752 6712
rect 13587 6681 13599 6684
rect 13541 6675 13599 6681
rect 15746 6672 15752 6684
rect 15804 6672 15810 6724
rect 15856 6712 15884 6752
rect 15933 6749 15945 6783
rect 15979 6780 15991 6783
rect 17034 6780 17040 6792
rect 15979 6752 17040 6780
rect 15979 6749 15991 6752
rect 15933 6743 15991 6749
rect 17034 6740 17040 6752
rect 17092 6740 17098 6792
rect 18417 6783 18475 6789
rect 18417 6749 18429 6783
rect 18463 6749 18475 6783
rect 18524 6780 18552 6888
rect 38672 6888 38884 6916
rect 18690 6808 18696 6860
rect 18748 6848 18754 6860
rect 21266 6848 21272 6860
rect 18748 6820 21272 6848
rect 18748 6808 18754 6820
rect 21266 6808 21272 6820
rect 21324 6848 21330 6860
rect 25961 6851 26019 6857
rect 25961 6848 25973 6851
rect 21324 6820 21956 6848
rect 21324 6808 21330 6820
rect 18524 6752 21128 6780
rect 18417 6743 18475 6749
rect 16850 6712 16856 6724
rect 15856 6684 16856 6712
rect 16850 6672 16856 6684
rect 16908 6672 16914 6724
rect 18432 6712 18460 6743
rect 18506 6712 18512 6724
rect 18432 6684 18512 6712
rect 18506 6672 18512 6684
rect 18564 6672 18570 6724
rect 18690 6672 18696 6724
rect 18748 6712 18754 6724
rect 20993 6715 21051 6721
rect 20993 6712 21005 6715
rect 18748 6684 21005 6712
rect 18748 6672 18754 6684
rect 20993 6681 21005 6684
rect 21039 6681 21051 6715
rect 21100 6712 21128 6752
rect 21726 6740 21732 6792
rect 21784 6780 21790 6792
rect 21821 6783 21879 6789
rect 21821 6780 21833 6783
rect 21784 6752 21833 6780
rect 21784 6740 21790 6752
rect 21821 6749 21833 6752
rect 21867 6749 21879 6783
rect 21928 6780 21956 6820
rect 22066 6820 25973 6848
rect 22066 6780 22094 6820
rect 25961 6817 25973 6820
rect 26007 6817 26019 6851
rect 38672 6848 38700 6888
rect 25961 6811 26019 6817
rect 30024 6820 32536 6848
rect 30024 6792 30052 6820
rect 32508 6792 32536 6820
rect 35360 6820 38700 6848
rect 38856 6848 38884 6888
rect 39853 6851 39911 6857
rect 39853 6848 39865 6851
rect 38856 6820 39865 6848
rect 21928 6752 22094 6780
rect 22143 6783 22201 6789
rect 21821 6743 21879 6749
rect 22143 6749 22155 6783
rect 22189 6780 22201 6783
rect 22462 6780 22468 6792
rect 22189 6752 22468 6780
rect 22189 6749 22201 6752
rect 22143 6743 22201 6749
rect 22462 6740 22468 6752
rect 22520 6740 22526 6792
rect 23474 6780 23480 6792
rect 23435 6752 23480 6780
rect 23474 6740 23480 6752
rect 23532 6740 23538 6792
rect 23569 6783 23627 6789
rect 23569 6749 23581 6783
rect 23615 6749 23627 6783
rect 23569 6743 23627 6749
rect 23584 6712 23612 6743
rect 23658 6740 23664 6792
rect 23716 6780 23722 6792
rect 23845 6783 23903 6789
rect 23716 6752 23761 6780
rect 23716 6740 23722 6752
rect 23845 6749 23857 6783
rect 23891 6780 23903 6783
rect 24026 6780 24032 6792
rect 23891 6752 24032 6780
rect 23891 6749 23903 6752
rect 23845 6743 23903 6749
rect 24026 6740 24032 6752
rect 24084 6740 24090 6792
rect 24302 6740 24308 6792
rect 24360 6780 24366 6792
rect 24578 6780 24584 6792
rect 24360 6752 24584 6780
rect 24360 6740 24366 6752
rect 24578 6740 24584 6752
rect 24636 6780 24642 6792
rect 24673 6783 24731 6789
rect 24673 6780 24685 6783
rect 24636 6752 24685 6780
rect 24636 6740 24642 6752
rect 24673 6749 24685 6752
rect 24719 6749 24731 6783
rect 24673 6743 24731 6749
rect 24765 6783 24823 6789
rect 24765 6749 24777 6783
rect 24811 6749 24823 6783
rect 24765 6743 24823 6749
rect 23934 6712 23940 6724
rect 21100 6684 23520 6712
rect 23584 6684 23940 6712
rect 20993 6675 21051 6681
rect 7285 6647 7343 6653
rect 7285 6613 7297 6647
rect 7331 6613 7343 6647
rect 7285 6607 7343 6613
rect 8018 6604 8024 6656
rect 8076 6644 8082 6656
rect 8113 6647 8171 6653
rect 8113 6644 8125 6647
rect 8076 6616 8125 6644
rect 8076 6604 8082 6616
rect 8113 6613 8125 6616
rect 8159 6613 8171 6647
rect 8938 6644 8944 6656
rect 8899 6616 8944 6644
rect 8113 6607 8171 6613
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 10505 6647 10563 6653
rect 10505 6613 10517 6647
rect 10551 6644 10563 6647
rect 10870 6644 10876 6656
rect 10551 6616 10876 6644
rect 10551 6613 10563 6616
rect 10505 6607 10563 6613
rect 10870 6604 10876 6616
rect 10928 6604 10934 6656
rect 14734 6604 14740 6656
rect 14792 6644 14798 6656
rect 14829 6647 14887 6653
rect 14829 6644 14841 6647
rect 14792 6616 14841 6644
rect 14792 6604 14798 6616
rect 14829 6613 14841 6616
rect 14875 6644 14887 6647
rect 15286 6644 15292 6656
rect 14875 6616 15292 6644
rect 14875 6613 14887 6616
rect 14829 6607 14887 6613
rect 15286 6604 15292 6616
rect 15344 6604 15350 6656
rect 15562 6644 15568 6656
rect 15523 6616 15568 6644
rect 15562 6604 15568 6616
rect 15620 6604 15626 6656
rect 16574 6644 16580 6656
rect 16535 6616 16580 6644
rect 16574 6604 16580 6616
rect 16632 6604 16638 6656
rect 17402 6644 17408 6656
rect 17363 6616 17408 6644
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 19058 6604 19064 6656
rect 19116 6644 19122 6656
rect 19245 6647 19303 6653
rect 19245 6644 19257 6647
rect 19116 6616 19257 6644
rect 19116 6604 19122 6616
rect 19245 6613 19257 6616
rect 19291 6613 19303 6647
rect 19978 6644 19984 6656
rect 19939 6616 19984 6644
rect 19245 6607 19303 6613
rect 19978 6604 19984 6616
rect 20036 6604 20042 6656
rect 20438 6644 20444 6656
rect 20399 6616 20444 6644
rect 20438 6604 20444 6616
rect 20496 6604 20502 6656
rect 23198 6644 23204 6656
rect 23159 6616 23204 6644
rect 23198 6604 23204 6616
rect 23256 6604 23262 6656
rect 23492 6644 23520 6684
rect 23934 6672 23940 6684
rect 23992 6712 23998 6724
rect 24780 6712 24808 6743
rect 24854 6740 24860 6792
rect 24912 6780 24918 6792
rect 25041 6783 25099 6789
rect 24912 6752 24957 6780
rect 24912 6740 24918 6752
rect 25041 6749 25053 6783
rect 25087 6749 25099 6783
rect 26234 6780 26240 6792
rect 26195 6752 26240 6780
rect 25041 6743 25099 6749
rect 23992 6684 24808 6712
rect 23992 6672 23998 6684
rect 24302 6644 24308 6656
rect 23492 6616 24308 6644
rect 24302 6604 24308 6616
rect 24360 6604 24366 6656
rect 24397 6647 24455 6653
rect 24397 6613 24409 6647
rect 24443 6644 24455 6647
rect 24670 6644 24676 6656
rect 24443 6616 24676 6644
rect 24443 6613 24455 6616
rect 24397 6607 24455 6613
rect 24670 6604 24676 6616
rect 24728 6604 24734 6656
rect 24762 6604 24768 6656
rect 24820 6644 24826 6656
rect 25056 6644 25084 6743
rect 26234 6740 26240 6752
rect 26292 6740 26298 6792
rect 27154 6740 27160 6792
rect 27212 6780 27218 6792
rect 27249 6783 27307 6789
rect 27249 6780 27261 6783
rect 27212 6752 27261 6780
rect 27212 6740 27218 6752
rect 27249 6749 27261 6752
rect 27295 6780 27307 6783
rect 29822 6780 29828 6792
rect 27295 6752 29828 6780
rect 27295 6749 27307 6752
rect 27249 6743 27307 6749
rect 29822 6740 29828 6752
rect 29880 6740 29886 6792
rect 30006 6780 30012 6792
rect 29919 6752 30012 6780
rect 30006 6740 30012 6752
rect 30064 6740 30070 6792
rect 32401 6783 32459 6789
rect 32401 6780 32413 6783
rect 31312 6752 32413 6780
rect 27338 6672 27344 6724
rect 27396 6712 27402 6724
rect 27494 6715 27552 6721
rect 27494 6712 27506 6715
rect 27396 6684 27506 6712
rect 27396 6672 27402 6684
rect 27494 6681 27506 6684
rect 27540 6681 27552 6715
rect 27494 6675 27552 6681
rect 24820 6616 25084 6644
rect 28629 6647 28687 6653
rect 24820 6604 24826 6616
rect 28629 6613 28641 6647
rect 28675 6644 28687 6647
rect 29270 6644 29276 6656
rect 28675 6616 29276 6644
rect 28675 6613 28687 6616
rect 28629 6607 28687 6613
rect 29270 6604 29276 6616
rect 29328 6604 29334 6656
rect 29840 6644 29868 6740
rect 31202 6644 31208 6656
rect 29840 6616 31208 6644
rect 31202 6604 31208 6616
rect 31260 6644 31266 6656
rect 31312 6653 31340 6752
rect 32401 6749 32413 6752
rect 32447 6749 32459 6783
rect 32401 6743 32459 6749
rect 32490 6740 32496 6792
rect 32548 6740 32554 6792
rect 32674 6789 32680 6792
rect 32668 6780 32680 6789
rect 32635 6752 32680 6780
rect 32668 6743 32680 6752
rect 32674 6740 32680 6743
rect 32732 6740 32738 6792
rect 34330 6740 34336 6792
rect 34388 6780 34394 6792
rect 35360 6789 35388 6820
rect 35345 6783 35403 6789
rect 35345 6780 35357 6783
rect 34388 6752 35357 6780
rect 34388 6740 34394 6752
rect 35345 6749 35357 6752
rect 35391 6749 35403 6783
rect 35345 6743 35403 6749
rect 35437 6783 35495 6789
rect 35437 6749 35449 6783
rect 35483 6749 35495 6783
rect 35437 6743 35495 6749
rect 35452 6712 35480 6743
rect 35526 6740 35532 6792
rect 35584 6780 35590 6792
rect 35713 6783 35771 6789
rect 35584 6752 35629 6780
rect 35584 6740 35590 6752
rect 35713 6749 35725 6783
rect 35759 6780 35771 6783
rect 35894 6780 35900 6792
rect 35759 6752 35900 6780
rect 35759 6749 35771 6752
rect 35713 6743 35771 6749
rect 35894 6740 35900 6752
rect 35952 6780 35958 6792
rect 36262 6780 36268 6792
rect 35952 6752 36268 6780
rect 35952 6740 35958 6752
rect 36262 6740 36268 6752
rect 36320 6740 36326 6792
rect 36630 6780 36636 6792
rect 36591 6752 36636 6780
rect 36630 6740 36636 6752
rect 36688 6740 36694 6792
rect 36814 6780 36820 6792
rect 36775 6752 36820 6780
rect 36814 6740 36820 6752
rect 36872 6740 36878 6792
rect 36909 6783 36967 6789
rect 36909 6749 36921 6783
rect 36955 6749 36967 6783
rect 36909 6743 36967 6749
rect 35802 6712 35808 6724
rect 35452 6684 35808 6712
rect 35802 6672 35808 6684
rect 35860 6672 35866 6724
rect 36924 6712 36952 6743
rect 36998 6740 37004 6792
rect 37056 6780 37062 6792
rect 38672 6789 38700 6820
rect 39853 6817 39865 6820
rect 39899 6817 39911 6851
rect 39853 6811 39911 6817
rect 37737 6783 37795 6789
rect 37737 6780 37749 6783
rect 37056 6752 37749 6780
rect 37056 6740 37062 6752
rect 37737 6749 37749 6752
rect 37783 6749 37795 6783
rect 37737 6743 37795 6749
rect 38657 6783 38715 6789
rect 38657 6749 38669 6783
rect 38703 6749 38715 6783
rect 38657 6743 38715 6749
rect 38749 6783 38807 6789
rect 38749 6749 38761 6783
rect 38795 6749 38807 6783
rect 38749 6743 38807 6749
rect 38764 6712 38792 6743
rect 38838 6740 38844 6792
rect 38896 6780 38902 6792
rect 38896 6752 38941 6780
rect 38896 6740 38902 6752
rect 39022 6740 39028 6792
rect 39080 6780 39086 6792
rect 39080 6752 39125 6780
rect 39080 6740 39086 6752
rect 38930 6712 38936 6724
rect 36924 6684 38936 6712
rect 38930 6672 38936 6684
rect 38988 6672 38994 6724
rect 31297 6647 31355 6653
rect 31297 6644 31309 6647
rect 31260 6616 31309 6644
rect 31260 6604 31266 6616
rect 31297 6613 31309 6616
rect 31343 6613 31355 6647
rect 31297 6607 31355 6613
rect 31386 6604 31392 6656
rect 31444 6644 31450 6656
rect 33781 6647 33839 6653
rect 33781 6644 33793 6647
rect 31444 6616 33793 6644
rect 31444 6604 31450 6616
rect 33781 6613 33793 6616
rect 33827 6613 33839 6647
rect 33781 6607 33839 6613
rect 35069 6647 35127 6653
rect 35069 6613 35081 6647
rect 35115 6644 35127 6647
rect 35434 6644 35440 6656
rect 35115 6616 35440 6644
rect 35115 6613 35127 6616
rect 35069 6607 35127 6613
rect 35434 6604 35440 6616
rect 35492 6604 35498 6656
rect 37274 6644 37280 6656
rect 37235 6616 37280 6644
rect 37274 6604 37280 6616
rect 37332 6604 37338 6656
rect 38378 6644 38384 6656
rect 38339 6616 38384 6644
rect 38378 6604 38384 6616
rect 38436 6604 38442 6656
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 3510 6400 3516 6452
rect 3568 6440 3574 6452
rect 3697 6443 3755 6449
rect 3697 6440 3709 6443
rect 3568 6412 3709 6440
rect 3568 6400 3574 6412
rect 3697 6409 3709 6412
rect 3743 6409 3755 6443
rect 9214 6440 9220 6452
rect 3697 6403 3755 6409
rect 6564 6412 9220 6440
rect 2584 6375 2642 6381
rect 2584 6341 2596 6375
rect 2630 6372 2642 6375
rect 2958 6372 2964 6384
rect 2630 6344 2964 6372
rect 2630 6341 2642 6344
rect 2584 6335 2642 6341
rect 2958 6332 2964 6344
rect 3016 6332 3022 6384
rect 6454 6372 6460 6384
rect 4908 6344 6460 6372
rect 4908 6313 4936 6344
rect 6454 6332 6460 6344
rect 6512 6332 6518 6384
rect 4893 6307 4951 6313
rect 4893 6273 4905 6307
rect 4939 6273 4951 6307
rect 4893 6267 4951 6273
rect 5077 6307 5135 6313
rect 5077 6273 5089 6307
rect 5123 6304 5135 6307
rect 5442 6304 5448 6316
rect 5123 6276 5448 6304
rect 5123 6273 5135 6276
rect 5077 6267 5135 6273
rect 5442 6264 5448 6276
rect 5500 6264 5506 6316
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 5994 6304 6000 6316
rect 5859 6276 6000 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 2314 6236 2320 6248
rect 2275 6208 2320 6236
rect 2314 6196 2320 6208
rect 2372 6196 2378 6248
rect 4433 6239 4491 6245
rect 4433 6205 4445 6239
rect 4479 6236 4491 6239
rect 5828 6236 5856 6267
rect 5994 6264 6000 6276
rect 6052 6264 6058 6316
rect 4479 6208 5856 6236
rect 4479 6205 4491 6208
rect 4433 6199 4491 6205
rect 3418 6128 3424 6180
rect 3476 6168 3482 6180
rect 6564 6168 6592 6412
rect 9214 6400 9220 6412
rect 9272 6400 9278 6452
rect 16574 6400 16580 6452
rect 16632 6440 16638 6452
rect 21266 6440 21272 6452
rect 16632 6412 21272 6440
rect 16632 6400 16638 6412
rect 21266 6400 21272 6412
rect 21324 6400 21330 6452
rect 23661 6443 23719 6449
rect 23661 6409 23673 6443
rect 23707 6440 23719 6443
rect 24210 6440 24216 6452
rect 23707 6412 24216 6440
rect 23707 6409 23719 6412
rect 23661 6403 23719 6409
rect 24210 6400 24216 6412
rect 24268 6400 24274 6452
rect 27798 6400 27804 6452
rect 27856 6440 27862 6452
rect 28261 6443 28319 6449
rect 28261 6440 28273 6443
rect 27856 6412 28273 6440
rect 27856 6400 27862 6412
rect 28261 6409 28273 6412
rect 28307 6409 28319 6443
rect 28261 6403 28319 6409
rect 29454 6400 29460 6452
rect 29512 6440 29518 6452
rect 29641 6443 29699 6449
rect 29641 6440 29653 6443
rect 29512 6412 29653 6440
rect 29512 6400 29518 6412
rect 29641 6409 29653 6412
rect 29687 6440 29699 6443
rect 30098 6440 30104 6452
rect 29687 6412 30104 6440
rect 29687 6409 29699 6412
rect 29641 6403 29699 6409
rect 30098 6400 30104 6412
rect 30156 6400 30162 6452
rect 30193 6443 30251 6449
rect 30193 6409 30205 6443
rect 30239 6440 30251 6443
rect 30466 6440 30472 6452
rect 30239 6412 30472 6440
rect 30239 6409 30251 6412
rect 30193 6403 30251 6409
rect 30466 6400 30472 6412
rect 30524 6400 30530 6452
rect 32217 6443 32275 6449
rect 32217 6409 32229 6443
rect 32263 6440 32275 6443
rect 32490 6440 32496 6452
rect 32263 6412 32496 6440
rect 32263 6409 32275 6412
rect 32217 6403 32275 6409
rect 32490 6400 32496 6412
rect 32548 6400 32554 6452
rect 35526 6400 35532 6452
rect 35584 6440 35590 6452
rect 35989 6443 36047 6449
rect 35989 6440 36001 6443
rect 35584 6412 36001 6440
rect 35584 6400 35590 6412
rect 35989 6409 36001 6412
rect 36035 6409 36047 6443
rect 35989 6403 36047 6409
rect 36814 6400 36820 6452
rect 36872 6440 36878 6452
rect 37277 6443 37335 6449
rect 37277 6440 37289 6443
rect 36872 6412 37289 6440
rect 36872 6400 36878 6412
rect 37277 6409 37289 6412
rect 37323 6409 37335 6443
rect 38746 6440 38752 6452
rect 37277 6403 37335 6409
rect 37476 6412 38752 6440
rect 6730 6332 6736 6384
rect 6788 6372 6794 6384
rect 13909 6375 13967 6381
rect 6788 6344 8984 6372
rect 6788 6332 6794 6344
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6273 6699 6307
rect 6641 6267 6699 6273
rect 7653 6307 7711 6313
rect 7653 6273 7665 6307
rect 7699 6304 7711 6307
rect 8478 6304 8484 6316
rect 7699 6276 8484 6304
rect 7699 6273 7711 6276
rect 7653 6267 7711 6273
rect 6656 6236 6684 6267
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 8956 6313 8984 6344
rect 13909 6341 13921 6375
rect 13955 6372 13967 6375
rect 14369 6375 14427 6381
rect 14369 6372 14381 6375
rect 13955 6344 14381 6372
rect 13955 6341 13967 6344
rect 13909 6335 13967 6341
rect 14369 6341 14381 6344
rect 14415 6372 14427 6375
rect 15194 6372 15200 6384
rect 14415 6344 15200 6372
rect 14415 6341 14427 6344
rect 14369 6335 14427 6341
rect 15194 6332 15200 6344
rect 15252 6332 15258 6384
rect 18782 6372 18788 6384
rect 18743 6344 18788 6372
rect 18782 6332 18788 6344
rect 18840 6372 18846 6384
rect 19245 6375 19303 6381
rect 19245 6372 19257 6375
rect 18840 6344 19257 6372
rect 18840 6332 18846 6344
rect 19245 6341 19257 6344
rect 19291 6341 19303 6375
rect 19245 6335 19303 6341
rect 19429 6375 19487 6381
rect 19429 6341 19441 6375
rect 19475 6372 19487 6375
rect 20714 6372 20720 6384
rect 19475 6344 20720 6372
rect 19475 6341 19487 6344
rect 19429 6335 19487 6341
rect 20714 6332 20720 6344
rect 20772 6332 20778 6384
rect 23385 6375 23443 6381
rect 23385 6341 23397 6375
rect 23431 6372 23443 6375
rect 24762 6372 24768 6384
rect 23431 6344 24768 6372
rect 23431 6341 23443 6344
rect 23385 6335 23443 6341
rect 24762 6332 24768 6344
rect 24820 6332 24826 6384
rect 25961 6375 26019 6381
rect 25961 6341 25973 6375
rect 26007 6372 26019 6375
rect 26142 6372 26148 6384
rect 26007 6344 26148 6372
rect 26007 6341 26019 6344
rect 25961 6335 26019 6341
rect 26142 6332 26148 6344
rect 26200 6372 26206 6384
rect 30006 6372 30012 6384
rect 26200 6344 30012 6372
rect 26200 6332 26206 6344
rect 30006 6332 30012 6344
rect 30064 6332 30070 6384
rect 34330 6372 34336 6384
rect 30208 6344 30880 6372
rect 30208 6316 30236 6344
rect 8941 6307 8999 6313
rect 8941 6273 8953 6307
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 9030 6264 9036 6316
rect 9088 6304 9094 6316
rect 9197 6307 9255 6313
rect 9197 6304 9209 6307
rect 9088 6276 9209 6304
rect 9088 6264 9094 6276
rect 9197 6273 9209 6276
rect 9243 6273 9255 6307
rect 9197 6267 9255 6273
rect 9490 6264 9496 6316
rect 9548 6304 9554 6316
rect 14734 6304 14740 6316
rect 9548 6276 14740 6304
rect 9548 6264 9554 6276
rect 14734 6264 14740 6276
rect 14792 6264 14798 6316
rect 16942 6304 16948 6316
rect 15856 6276 16804 6304
rect 16903 6276 16948 6304
rect 6822 6236 6828 6248
rect 6656 6208 6828 6236
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 6917 6239 6975 6245
rect 6917 6205 6929 6239
rect 6963 6236 6975 6239
rect 7282 6236 7288 6248
rect 6963 6208 7288 6236
rect 6963 6205 6975 6208
rect 6917 6199 6975 6205
rect 7282 6196 7288 6208
rect 7340 6196 7346 6248
rect 13262 6196 13268 6248
rect 13320 6236 13326 6248
rect 15856 6236 15884 6276
rect 16022 6236 16028 6248
rect 13320 6208 15884 6236
rect 15983 6208 16028 6236
rect 13320 6196 13326 6208
rect 16022 6196 16028 6208
rect 16080 6196 16086 6248
rect 16574 6196 16580 6248
rect 16632 6236 16638 6248
rect 16669 6239 16727 6245
rect 16669 6236 16681 6239
rect 16632 6208 16681 6236
rect 16632 6196 16638 6208
rect 16669 6205 16681 6208
rect 16715 6205 16727 6239
rect 16776 6236 16804 6276
rect 16942 6264 16948 6276
rect 17000 6264 17006 6316
rect 18598 6304 18604 6316
rect 18559 6276 18604 6304
rect 18598 6264 18604 6276
rect 18656 6264 18662 6316
rect 23109 6307 23167 6313
rect 23109 6304 23121 6307
rect 22066 6276 23121 6304
rect 18138 6236 18144 6248
rect 16776 6208 18144 6236
rect 16669 6199 16727 6205
rect 18138 6196 18144 6208
rect 18196 6236 18202 6248
rect 18782 6236 18788 6248
rect 18196 6208 18788 6236
rect 18196 6196 18202 6208
rect 18782 6196 18788 6208
rect 18840 6196 18846 6248
rect 21726 6196 21732 6248
rect 21784 6236 21790 6248
rect 21821 6239 21879 6245
rect 21821 6236 21833 6239
rect 21784 6208 21833 6236
rect 21784 6196 21790 6208
rect 21821 6205 21833 6208
rect 21867 6205 21879 6239
rect 22066 6236 22094 6276
rect 23109 6273 23121 6276
rect 23155 6273 23167 6307
rect 23109 6267 23167 6273
rect 23293 6307 23351 6313
rect 23293 6273 23305 6307
rect 23339 6273 23351 6307
rect 23474 6304 23480 6316
rect 23435 6276 23480 6304
rect 23293 6267 23351 6273
rect 21821 6199 21879 6205
rect 21928 6208 22094 6236
rect 22143 6239 22201 6245
rect 3476 6140 6592 6168
rect 6733 6171 6791 6177
rect 3476 6128 3482 6140
rect 6733 6137 6745 6171
rect 6779 6168 6791 6171
rect 7006 6168 7012 6180
rect 6779 6140 7012 6168
rect 6779 6137 6791 6140
rect 6733 6131 6791 6137
rect 7006 6128 7012 6140
rect 7064 6168 7070 6180
rect 7837 6171 7895 6177
rect 7837 6168 7849 6171
rect 7064 6140 7849 6168
rect 7064 6128 7070 6140
rect 7837 6137 7849 6140
rect 7883 6137 7895 6171
rect 7837 6131 7895 6137
rect 10042 6128 10048 6180
rect 10100 6168 10106 6180
rect 10321 6171 10379 6177
rect 10321 6168 10333 6171
rect 10100 6140 10333 6168
rect 10100 6128 10106 6140
rect 10321 6137 10333 6140
rect 10367 6168 10379 6171
rect 11054 6168 11060 6180
rect 10367 6140 11060 6168
rect 10367 6137 10379 6140
rect 10321 6131 10379 6137
rect 11054 6128 11060 6140
rect 11112 6128 11118 6180
rect 11793 6171 11851 6177
rect 11793 6137 11805 6171
rect 11839 6168 11851 6171
rect 13814 6168 13820 6180
rect 11839 6140 13820 6168
rect 11839 6137 11851 6140
rect 11793 6131 11851 6137
rect 13814 6128 13820 6140
rect 13872 6128 13878 6180
rect 15746 6128 15752 6180
rect 15804 6168 15810 6180
rect 21928 6168 21956 6208
rect 22143 6205 22155 6239
rect 22189 6236 22201 6239
rect 22738 6236 22744 6248
rect 22189 6208 22744 6236
rect 22189 6205 22201 6208
rect 22143 6199 22201 6205
rect 22738 6196 22744 6208
rect 22796 6236 22802 6248
rect 23308 6236 23336 6267
rect 23474 6264 23480 6276
rect 23532 6264 23538 6316
rect 27249 6307 27307 6313
rect 24504 6276 27016 6304
rect 22796 6208 23336 6236
rect 22796 6196 22802 6208
rect 24504 6168 24532 6276
rect 24578 6196 24584 6248
rect 24636 6236 24642 6248
rect 24636 6208 25176 6236
rect 24636 6196 24642 6208
rect 15804 6140 21956 6168
rect 22066 6140 24532 6168
rect 25148 6168 25176 6208
rect 26878 6196 26884 6248
rect 26936 6236 26942 6248
rect 26988 6245 27016 6276
rect 27249 6273 27261 6307
rect 27295 6304 27307 6307
rect 27982 6304 27988 6316
rect 27295 6276 27988 6304
rect 27295 6273 27307 6276
rect 27249 6267 27307 6273
rect 27982 6264 27988 6276
rect 28040 6264 28046 6316
rect 28445 6307 28503 6313
rect 28445 6273 28457 6307
rect 28491 6273 28503 6307
rect 28445 6267 28503 6273
rect 26973 6239 27031 6245
rect 26973 6236 26985 6239
rect 26936 6208 26985 6236
rect 26936 6196 26942 6208
rect 26973 6205 26985 6208
rect 27019 6205 27031 6239
rect 28460 6236 28488 6267
rect 28626 6264 28632 6316
rect 28684 6304 28690 6316
rect 28684 6276 29684 6304
rect 28684 6264 28690 6276
rect 29270 6236 29276 6248
rect 28460 6208 29276 6236
rect 26973 6199 27031 6205
rect 29270 6196 29276 6208
rect 29328 6196 29334 6248
rect 29656 6236 29684 6276
rect 30190 6264 30196 6316
rect 30248 6264 30254 6316
rect 30282 6264 30288 6316
rect 30340 6304 30346 6316
rect 30423 6307 30481 6313
rect 30423 6304 30435 6307
rect 30340 6276 30435 6304
rect 30340 6264 30346 6276
rect 30423 6273 30435 6276
rect 30469 6273 30481 6307
rect 30558 6304 30564 6316
rect 30519 6276 30564 6304
rect 30423 6267 30481 6273
rect 30558 6264 30564 6276
rect 30616 6264 30622 6316
rect 30650 6264 30656 6316
rect 30708 6304 30714 6316
rect 30852 6313 30880 6344
rect 31726 6344 34336 6372
rect 30837 6307 30895 6313
rect 30708 6276 30753 6304
rect 30708 6264 30714 6276
rect 30837 6273 30849 6307
rect 30883 6273 30895 6307
rect 30837 6267 30895 6273
rect 31478 6236 31484 6248
rect 29656 6208 31484 6236
rect 31478 6196 31484 6208
rect 31536 6196 31542 6248
rect 31726 6236 31754 6344
rect 34330 6332 34336 6344
rect 34388 6332 34394 6384
rect 35802 6372 35808 6384
rect 35268 6344 35808 6372
rect 35268 6313 35296 6344
rect 35802 6332 35808 6344
rect 35860 6332 35866 6384
rect 37182 6332 37188 6384
rect 37240 6372 37246 6384
rect 37476 6381 37504 6412
rect 38746 6400 38752 6412
rect 38804 6400 38810 6452
rect 39666 6440 39672 6452
rect 39627 6412 39672 6440
rect 39666 6400 39672 6412
rect 39724 6400 39730 6452
rect 37461 6375 37519 6381
rect 37461 6372 37473 6375
rect 37240 6344 37473 6372
rect 37240 6332 37246 6344
rect 37461 6341 37473 6344
rect 37507 6341 37519 6375
rect 37642 6372 37648 6384
rect 37603 6344 37648 6372
rect 37461 6335 37519 6341
rect 37642 6332 37648 6344
rect 37700 6332 37706 6384
rect 38378 6332 38384 6384
rect 38436 6372 38442 6384
rect 38534 6375 38592 6381
rect 38534 6372 38546 6375
rect 38436 6344 38546 6372
rect 38436 6332 38442 6344
rect 38534 6341 38546 6344
rect 38580 6341 38592 6375
rect 38534 6335 38592 6341
rect 35161 6307 35219 6313
rect 35161 6304 35173 6307
rect 31588 6208 31754 6236
rect 33796 6276 35173 6304
rect 31588 6168 31616 6208
rect 25148 6140 31616 6168
rect 15804 6128 15810 6140
rect 1854 6100 1860 6112
rect 1815 6072 1860 6100
rect 1854 6060 1860 6072
rect 1912 6060 1918 6112
rect 5074 6100 5080 6112
rect 5035 6072 5080 6100
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 5626 6100 5632 6112
rect 5587 6072 5632 6100
rect 5626 6060 5632 6072
rect 5684 6060 5690 6112
rect 6638 6100 6644 6112
rect 6599 6072 6644 6100
rect 6638 6060 6644 6072
rect 6696 6060 6702 6112
rect 8481 6103 8539 6109
rect 8481 6069 8493 6103
rect 8527 6100 8539 6103
rect 9950 6100 9956 6112
rect 8527 6072 9956 6100
rect 8527 6069 8539 6072
rect 8481 6063 8539 6069
rect 9950 6060 9956 6072
rect 10008 6060 10014 6112
rect 10502 6060 10508 6112
rect 10560 6100 10566 6112
rect 10781 6103 10839 6109
rect 10781 6100 10793 6103
rect 10560 6072 10793 6100
rect 10560 6060 10566 6072
rect 10781 6069 10793 6072
rect 10827 6069 10839 6103
rect 10781 6063 10839 6069
rect 12158 6060 12164 6112
rect 12216 6100 12222 6112
rect 12253 6103 12311 6109
rect 12253 6100 12265 6103
rect 12216 6072 12265 6100
rect 12216 6060 12222 6072
rect 12253 6069 12265 6072
rect 12299 6069 12311 6103
rect 12253 6063 12311 6069
rect 13265 6103 13323 6109
rect 13265 6069 13277 6103
rect 13311 6100 13323 6103
rect 15286 6100 15292 6112
rect 13311 6072 15292 6100
rect 13311 6069 13323 6072
rect 13265 6063 13323 6069
rect 15286 6060 15292 6072
rect 15344 6060 15350 6112
rect 18138 6060 18144 6112
rect 18196 6100 18202 6112
rect 18417 6103 18475 6109
rect 18417 6100 18429 6103
rect 18196 6072 18429 6100
rect 18196 6060 18202 6072
rect 18417 6069 18429 6072
rect 18463 6069 18475 6103
rect 18417 6063 18475 6069
rect 19334 6060 19340 6112
rect 19392 6100 19398 6112
rect 19613 6103 19671 6109
rect 19613 6100 19625 6103
rect 19392 6072 19625 6100
rect 19392 6060 19398 6072
rect 19613 6069 19625 6072
rect 19659 6069 19671 6103
rect 20162 6100 20168 6112
rect 20123 6072 20168 6100
rect 19613 6063 19671 6069
rect 20162 6060 20168 6072
rect 20220 6060 20226 6112
rect 20622 6100 20628 6112
rect 20583 6072 20628 6100
rect 20622 6060 20628 6072
rect 20680 6060 20686 6112
rect 20714 6060 20720 6112
rect 20772 6100 20778 6112
rect 21177 6103 21235 6109
rect 21177 6100 21189 6103
rect 20772 6072 21189 6100
rect 20772 6060 20778 6072
rect 21177 6069 21189 6072
rect 21223 6069 21235 6103
rect 21177 6063 21235 6069
rect 21266 6060 21272 6112
rect 21324 6100 21330 6112
rect 22066 6100 22094 6140
rect 21324 6072 22094 6100
rect 24673 6103 24731 6109
rect 21324 6060 21330 6072
rect 24673 6069 24685 6103
rect 24719 6100 24731 6103
rect 24946 6100 24952 6112
rect 24719 6072 24952 6100
rect 24719 6069 24731 6072
rect 24673 6063 24731 6069
rect 24946 6060 24952 6072
rect 25004 6060 25010 6112
rect 30098 6060 30104 6112
rect 30156 6100 30162 6112
rect 33796 6109 33824 6276
rect 34716 6168 34744 6276
rect 35161 6273 35173 6276
rect 35207 6273 35219 6307
rect 35161 6267 35219 6273
rect 35250 6307 35308 6313
rect 35250 6273 35262 6307
rect 35296 6273 35308 6307
rect 35250 6267 35308 6273
rect 35342 6264 35348 6316
rect 35400 6304 35406 6316
rect 35529 6307 35587 6313
rect 35400 6276 35445 6304
rect 35400 6264 35406 6276
rect 35529 6273 35541 6307
rect 35575 6304 35587 6307
rect 35894 6304 35900 6316
rect 35575 6276 35900 6304
rect 35575 6273 35587 6276
rect 35529 6267 35587 6273
rect 35894 6264 35900 6276
rect 35952 6264 35958 6316
rect 36170 6304 36176 6316
rect 36131 6276 36176 6304
rect 36170 6264 36176 6276
rect 36228 6264 36234 6316
rect 36357 6307 36415 6313
rect 36357 6273 36369 6307
rect 36403 6273 36415 6307
rect 36357 6267 36415 6273
rect 34790 6196 34796 6248
rect 34848 6236 34854 6248
rect 36372 6236 36400 6267
rect 38286 6236 38292 6248
rect 34848 6208 36400 6236
rect 38247 6208 38292 6236
rect 34848 6196 34854 6208
rect 38286 6196 38292 6208
rect 38344 6196 38350 6248
rect 36998 6168 37004 6180
rect 34716 6140 37004 6168
rect 36998 6128 37004 6140
rect 37056 6128 37062 6180
rect 58158 6168 58164 6180
rect 58119 6140 58164 6168
rect 58158 6128 58164 6140
rect 58216 6128 58222 6180
rect 33781 6103 33839 6109
rect 33781 6100 33793 6103
rect 30156 6072 33793 6100
rect 30156 6060 30162 6072
rect 33781 6069 33793 6072
rect 33827 6069 33839 6103
rect 33781 6063 33839 6069
rect 34885 6103 34943 6109
rect 34885 6069 34897 6103
rect 34931 6100 34943 6103
rect 35802 6100 35808 6112
rect 34931 6072 35808 6100
rect 34931 6069 34943 6072
rect 34885 6063 34943 6069
rect 35802 6060 35808 6072
rect 35860 6060 35866 6112
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 2314 5856 2320 5908
rect 2372 5896 2378 5908
rect 4617 5899 4675 5905
rect 4617 5896 4629 5899
rect 2372 5868 4629 5896
rect 2372 5856 2378 5868
rect 4617 5865 4629 5868
rect 4663 5896 4675 5899
rect 6730 5896 6736 5908
rect 4663 5868 6736 5896
rect 4663 5865 4675 5868
rect 4617 5859 4675 5865
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 7742 5896 7748 5908
rect 7703 5868 7748 5896
rect 7742 5856 7748 5868
rect 7800 5896 7806 5908
rect 13262 5896 13268 5908
rect 7800 5868 13268 5896
rect 7800 5856 7806 5868
rect 13262 5856 13268 5868
rect 13320 5856 13326 5908
rect 15470 5896 15476 5908
rect 13464 5868 15476 5896
rect 4982 5788 4988 5840
rect 5040 5828 5046 5840
rect 9030 5828 9036 5840
rect 5040 5800 9036 5828
rect 5040 5788 5046 5800
rect 9030 5788 9036 5800
rect 9088 5788 9094 5840
rect 9214 5788 9220 5840
rect 9272 5828 9278 5840
rect 13464 5837 13492 5868
rect 15470 5856 15476 5868
rect 15528 5896 15534 5908
rect 15657 5899 15715 5905
rect 15528 5868 15608 5896
rect 15528 5856 15534 5868
rect 13449 5831 13507 5837
rect 13449 5828 13461 5831
rect 9272 5800 13461 5828
rect 9272 5788 9278 5800
rect 13449 5797 13461 5800
rect 13495 5797 13507 5831
rect 13449 5791 13507 5797
rect 9125 5763 9183 5769
rect 9125 5729 9137 5763
rect 9171 5760 9183 5763
rect 12986 5760 12992 5772
rect 9171 5732 12992 5760
rect 9171 5729 9183 5732
rect 9125 5723 9183 5729
rect 12986 5720 12992 5732
rect 13044 5720 13050 5772
rect 15580 5760 15608 5868
rect 15657 5865 15669 5899
rect 15703 5896 15715 5899
rect 15746 5896 15752 5908
rect 15703 5868 15752 5896
rect 15703 5865 15715 5868
rect 15657 5859 15715 5865
rect 15746 5856 15752 5868
rect 15804 5856 15810 5908
rect 18598 5856 18604 5908
rect 18656 5896 18662 5908
rect 20625 5899 20683 5905
rect 20625 5896 20637 5899
rect 18656 5868 20637 5896
rect 18656 5856 18662 5868
rect 20625 5865 20637 5868
rect 20671 5896 20683 5899
rect 20671 5868 22094 5896
rect 20671 5865 20683 5868
rect 20625 5859 20683 5865
rect 17770 5828 17776 5840
rect 17420 5800 17776 5828
rect 15580 5732 16436 5760
rect 2222 5692 2228 5704
rect 2183 5664 2228 5692
rect 2222 5652 2228 5664
rect 2280 5652 2286 5704
rect 5810 5652 5816 5704
rect 5868 5692 5874 5704
rect 5905 5695 5963 5701
rect 5905 5692 5917 5695
rect 5868 5664 5917 5692
rect 5868 5652 5874 5664
rect 5905 5661 5917 5664
rect 5951 5661 5963 5695
rect 6914 5692 6920 5704
rect 6875 5664 6920 5692
rect 5905 5655 5963 5661
rect 6914 5652 6920 5664
rect 6972 5652 6978 5704
rect 7006 5652 7012 5704
rect 7064 5692 7070 5704
rect 7064 5664 7109 5692
rect 7064 5652 7070 5664
rect 7374 5652 7380 5704
rect 7432 5692 7438 5704
rect 7561 5695 7619 5701
rect 7561 5692 7573 5695
rect 7432 5664 7573 5692
rect 7432 5652 7438 5664
rect 7561 5661 7573 5664
rect 7607 5661 7619 5695
rect 7561 5655 7619 5661
rect 8846 5652 8852 5704
rect 8904 5692 8910 5704
rect 9214 5692 9220 5704
rect 8904 5664 9220 5692
rect 8904 5652 8910 5664
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 9769 5695 9827 5701
rect 9769 5661 9781 5695
rect 9815 5692 9827 5695
rect 10226 5692 10232 5704
rect 9815 5664 10232 5692
rect 9815 5661 9827 5664
rect 9769 5655 9827 5661
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 10413 5695 10471 5701
rect 10413 5661 10425 5695
rect 10459 5692 10471 5695
rect 10778 5692 10784 5704
rect 10459 5664 10784 5692
rect 10459 5661 10471 5664
rect 10413 5655 10471 5661
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 11057 5695 11115 5701
rect 11057 5661 11069 5695
rect 11103 5692 11115 5695
rect 11330 5692 11336 5704
rect 11103 5664 11336 5692
rect 11103 5661 11115 5664
rect 11057 5655 11115 5661
rect 11330 5652 11336 5664
rect 11388 5652 11394 5704
rect 11701 5695 11759 5701
rect 11701 5661 11713 5695
rect 11747 5692 11759 5695
rect 11882 5692 11888 5704
rect 11747 5664 11888 5692
rect 11747 5661 11759 5664
rect 11701 5655 11759 5661
rect 11882 5652 11888 5664
rect 11940 5652 11946 5704
rect 12345 5695 12403 5701
rect 12345 5661 12357 5695
rect 12391 5692 12403 5695
rect 12434 5692 12440 5704
rect 12391 5664 12440 5692
rect 12391 5661 12403 5664
rect 12345 5655 12403 5661
rect 12434 5652 12440 5664
rect 12492 5652 12498 5704
rect 12710 5652 12716 5704
rect 12768 5692 12774 5704
rect 12805 5695 12863 5701
rect 12805 5692 12817 5695
rect 12768 5664 12817 5692
rect 12768 5652 12774 5664
rect 12805 5661 12817 5664
rect 12851 5661 12863 5695
rect 12805 5655 12863 5661
rect 14277 5695 14335 5701
rect 14277 5661 14289 5695
rect 14323 5692 14335 5695
rect 14826 5692 14832 5704
rect 14323 5664 14832 5692
rect 14323 5661 14335 5664
rect 14277 5655 14335 5661
rect 14826 5652 14832 5664
rect 14884 5692 14890 5704
rect 16022 5692 16028 5704
rect 14884 5664 16028 5692
rect 14884 5652 14890 5664
rect 16022 5652 16028 5664
rect 16080 5652 16086 5704
rect 16408 5701 16436 5732
rect 17310 5720 17316 5772
rect 17368 5760 17374 5772
rect 17420 5769 17448 5800
rect 17770 5788 17776 5800
rect 17828 5828 17834 5840
rect 17828 5800 18460 5828
rect 17828 5788 17834 5800
rect 17405 5763 17463 5769
rect 17405 5760 17417 5763
rect 17368 5732 17417 5760
rect 17368 5720 17374 5732
rect 17405 5729 17417 5732
rect 17451 5729 17463 5763
rect 17405 5723 17463 5729
rect 16393 5695 16451 5701
rect 16393 5661 16405 5695
rect 16439 5661 16451 5695
rect 16393 5655 16451 5661
rect 16485 5695 16543 5701
rect 16485 5661 16497 5695
rect 16531 5661 16543 5695
rect 16485 5655 16543 5661
rect 3237 5627 3295 5633
rect 3237 5593 3249 5627
rect 3283 5624 3295 5627
rect 6822 5624 6828 5636
rect 3283 5596 6828 5624
rect 3283 5593 3295 5596
rect 3237 5587 3295 5593
rect 6822 5584 6828 5596
rect 6880 5584 6886 5636
rect 8389 5627 8447 5633
rect 8389 5593 8401 5627
rect 8435 5624 8447 5627
rect 13170 5624 13176 5636
rect 8435 5596 13176 5624
rect 8435 5593 8447 5596
rect 8389 5587 8447 5593
rect 13170 5584 13176 5596
rect 13228 5584 13234 5636
rect 14550 5633 14556 5636
rect 14544 5587 14556 5633
rect 14608 5624 14614 5636
rect 14608 5596 14644 5624
rect 14550 5584 14556 5587
rect 14608 5584 14614 5596
rect 15378 5584 15384 5636
rect 15436 5624 15442 5636
rect 16500 5624 16528 5655
rect 16574 5652 16580 5704
rect 16632 5692 16638 5704
rect 16632 5664 16677 5692
rect 16632 5652 16638 5664
rect 16758 5652 16764 5704
rect 16816 5692 16822 5704
rect 16942 5692 16948 5704
rect 16816 5664 16948 5692
rect 16816 5652 16822 5664
rect 16942 5652 16948 5664
rect 17000 5692 17006 5704
rect 17862 5692 17868 5704
rect 17000 5664 17868 5692
rect 17000 5652 17006 5664
rect 17862 5652 17868 5664
rect 17920 5692 17926 5704
rect 17957 5695 18015 5701
rect 17957 5692 17969 5695
rect 17920 5664 17969 5692
rect 17920 5652 17926 5664
rect 17957 5661 17969 5664
rect 18003 5661 18015 5695
rect 18138 5692 18144 5704
rect 18099 5664 18144 5692
rect 17957 5655 18015 5661
rect 18138 5652 18144 5664
rect 18196 5652 18202 5704
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5661 18291 5695
rect 18233 5655 18291 5661
rect 18325 5695 18383 5701
rect 18325 5661 18337 5695
rect 18371 5692 18383 5695
rect 18432 5692 18460 5800
rect 19242 5760 19248 5772
rect 19203 5732 19248 5760
rect 19242 5720 19248 5732
rect 19300 5720 19306 5772
rect 22066 5760 22094 5868
rect 23658 5856 23664 5908
rect 23716 5896 23722 5908
rect 24949 5899 25007 5905
rect 24949 5896 24961 5899
rect 23716 5868 24961 5896
rect 23716 5856 23722 5868
rect 24949 5865 24961 5868
rect 24995 5865 25007 5899
rect 26142 5896 26148 5908
rect 26103 5868 26148 5896
rect 24949 5859 25007 5865
rect 26142 5856 26148 5868
rect 26200 5856 26206 5908
rect 26878 5896 26884 5908
rect 26839 5868 26884 5896
rect 26878 5856 26884 5868
rect 26936 5856 26942 5908
rect 30282 5856 30288 5908
rect 30340 5896 30346 5908
rect 31389 5899 31447 5905
rect 31389 5896 31401 5899
rect 30340 5868 31401 5896
rect 30340 5856 30346 5868
rect 31389 5865 31401 5868
rect 31435 5865 31447 5899
rect 31389 5859 31447 5865
rect 32490 5856 32496 5908
rect 32548 5896 32554 5908
rect 36541 5899 36599 5905
rect 36541 5896 36553 5899
rect 32548 5868 36553 5896
rect 32548 5856 32554 5868
rect 36541 5865 36553 5868
rect 36587 5865 36599 5899
rect 36541 5859 36599 5865
rect 23109 5831 23167 5837
rect 23109 5797 23121 5831
rect 23155 5828 23167 5831
rect 23750 5828 23756 5840
rect 23155 5800 23756 5828
rect 23155 5797 23167 5800
rect 23109 5791 23167 5797
rect 23750 5788 23756 5800
rect 23808 5788 23814 5840
rect 24489 5831 24547 5837
rect 24489 5797 24501 5831
rect 24535 5828 24547 5831
rect 24578 5828 24584 5840
rect 24535 5800 24584 5828
rect 24535 5797 24547 5800
rect 24489 5791 24547 5797
rect 24578 5788 24584 5800
rect 24636 5788 24642 5840
rect 32585 5831 32643 5837
rect 32585 5828 32597 5831
rect 30484 5800 32597 5828
rect 27430 5760 27436 5772
rect 22066 5732 27436 5760
rect 27430 5720 27436 5732
rect 27488 5720 27494 5772
rect 30098 5760 30104 5772
rect 27540 5732 30104 5760
rect 22557 5695 22615 5701
rect 22557 5692 22569 5695
rect 18371 5664 18460 5692
rect 22066 5664 22569 5692
rect 18371 5661 18383 5664
rect 18325 5655 18383 5661
rect 18248 5624 18276 5655
rect 18506 5624 18512 5636
rect 15436 5596 18512 5624
rect 15436 5584 15442 5596
rect 18506 5584 18512 5596
rect 18564 5584 18570 5636
rect 18601 5627 18659 5633
rect 18601 5593 18613 5627
rect 18647 5624 18659 5627
rect 19490 5627 19548 5633
rect 19490 5624 19502 5627
rect 18647 5596 19502 5624
rect 18647 5593 18659 5596
rect 18601 5587 18659 5593
rect 19490 5593 19502 5596
rect 19536 5593 19548 5627
rect 22066 5624 22094 5664
rect 22557 5661 22569 5664
rect 22603 5661 22615 5695
rect 22738 5692 22744 5704
rect 22699 5664 22744 5692
rect 22557 5655 22615 5661
rect 22738 5652 22744 5664
rect 22796 5652 22802 5704
rect 22925 5695 22983 5701
rect 22925 5661 22937 5695
rect 22971 5692 22983 5695
rect 23382 5692 23388 5704
rect 22971 5664 23388 5692
rect 22971 5661 22983 5664
rect 22925 5655 22983 5661
rect 23382 5652 23388 5664
rect 23440 5652 23446 5704
rect 24762 5652 24768 5704
rect 24820 5692 24826 5704
rect 25133 5695 25191 5701
rect 25133 5692 25145 5695
rect 24820 5664 25145 5692
rect 24820 5652 24826 5664
rect 25133 5661 25145 5664
rect 25179 5661 25191 5695
rect 25133 5655 25191 5661
rect 25314 5652 25320 5704
rect 25372 5692 25378 5704
rect 25774 5692 25780 5704
rect 25372 5664 25780 5692
rect 25372 5652 25378 5664
rect 25774 5652 25780 5664
rect 25832 5652 25838 5704
rect 19490 5587 19548 5593
rect 19628 5596 22094 5624
rect 22833 5627 22891 5633
rect 1762 5556 1768 5568
rect 1723 5528 1768 5556
rect 1762 5516 1768 5528
rect 1820 5516 1826 5568
rect 2409 5559 2467 5565
rect 2409 5525 2421 5559
rect 2455 5556 2467 5559
rect 2498 5556 2504 5568
rect 2455 5528 2504 5556
rect 2455 5525 2467 5528
rect 2409 5519 2467 5525
rect 2498 5516 2504 5528
rect 2556 5516 2562 5568
rect 6730 5556 6736 5568
rect 6691 5528 6736 5556
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 15286 5516 15292 5568
rect 15344 5556 15350 5568
rect 15470 5556 15476 5568
rect 15344 5528 15476 5556
rect 15344 5516 15350 5528
rect 15470 5516 15476 5528
rect 15528 5516 15534 5568
rect 16114 5556 16120 5568
rect 16075 5528 16120 5556
rect 16114 5516 16120 5528
rect 16172 5516 16178 5568
rect 17586 5516 17592 5568
rect 17644 5556 17650 5568
rect 19628 5556 19656 5596
rect 22833 5593 22845 5627
rect 22879 5624 22891 5627
rect 24578 5624 24584 5636
rect 22879 5596 24584 5624
rect 22879 5593 22891 5596
rect 22833 5587 22891 5593
rect 24578 5584 24584 5596
rect 24636 5584 24642 5636
rect 21358 5556 21364 5568
rect 17644 5528 19656 5556
rect 21319 5528 21364 5556
rect 17644 5516 17650 5528
rect 21358 5516 21364 5528
rect 21416 5516 21422 5568
rect 21910 5556 21916 5568
rect 21871 5528 21916 5556
rect 21910 5516 21916 5528
rect 21968 5516 21974 5568
rect 23566 5516 23572 5568
rect 23624 5556 23630 5568
rect 23661 5559 23719 5565
rect 23661 5556 23673 5559
rect 23624 5528 23673 5556
rect 23624 5516 23630 5528
rect 23661 5525 23673 5528
rect 23707 5556 23719 5559
rect 27540 5556 27568 5732
rect 30098 5720 30104 5732
rect 30156 5720 30162 5772
rect 28169 5695 28227 5701
rect 28169 5661 28181 5695
rect 28215 5692 28227 5695
rect 28442 5692 28448 5704
rect 28215 5664 28448 5692
rect 28215 5661 28227 5664
rect 28169 5655 28227 5661
rect 28442 5652 28448 5664
rect 28500 5652 28506 5704
rect 30190 5652 30196 5704
rect 30248 5692 30254 5704
rect 30484 5701 30512 5800
rect 32585 5797 32597 5800
rect 32631 5797 32643 5831
rect 34698 5828 34704 5840
rect 34659 5800 34704 5828
rect 32585 5791 32643 5797
rect 34698 5788 34704 5800
rect 34756 5788 34762 5840
rect 30285 5695 30343 5701
rect 30285 5692 30297 5695
rect 30248 5664 30297 5692
rect 30248 5652 30254 5664
rect 30285 5661 30297 5664
rect 30331 5661 30343 5695
rect 30285 5655 30343 5661
rect 30469 5695 30527 5701
rect 30469 5661 30481 5695
rect 30515 5661 30527 5695
rect 30469 5655 30527 5661
rect 30561 5695 30619 5701
rect 30561 5661 30573 5695
rect 30607 5661 30619 5695
rect 30561 5655 30619 5661
rect 28353 5627 28411 5633
rect 28353 5593 28365 5627
rect 28399 5624 28411 5627
rect 28626 5624 28632 5636
rect 28399 5596 28632 5624
rect 28399 5593 28411 5596
rect 28353 5587 28411 5593
rect 28626 5584 28632 5596
rect 28684 5584 28690 5636
rect 30576 5624 30604 5655
rect 30650 5652 30656 5704
rect 30708 5701 30714 5704
rect 30708 5695 30731 5701
rect 30719 5661 30731 5695
rect 30708 5655 30731 5661
rect 31573 5695 31631 5701
rect 31573 5661 31585 5695
rect 31619 5692 31631 5695
rect 32122 5692 32128 5704
rect 31619 5664 32128 5692
rect 31619 5661 31631 5664
rect 31573 5655 31631 5661
rect 30708 5652 30714 5655
rect 32122 5652 32128 5664
rect 32180 5652 32186 5704
rect 32398 5692 32404 5704
rect 32359 5664 32404 5692
rect 32398 5652 32404 5664
rect 32456 5652 32462 5704
rect 35802 5652 35808 5704
rect 35860 5701 35866 5704
rect 35860 5692 35872 5701
rect 36081 5695 36139 5701
rect 35860 5664 35905 5692
rect 35860 5655 35872 5664
rect 36081 5661 36093 5695
rect 36127 5661 36139 5695
rect 36081 5655 36139 5661
rect 35860 5652 35866 5655
rect 30576 5596 30788 5624
rect 23707 5528 27568 5556
rect 23707 5525 23719 5528
rect 23661 5519 23719 5525
rect 27798 5516 27804 5568
rect 27856 5556 27862 5568
rect 27985 5559 28043 5565
rect 27985 5556 27997 5559
rect 27856 5528 27997 5556
rect 27856 5516 27862 5528
rect 27985 5525 27997 5528
rect 28031 5525 28043 5559
rect 27985 5519 28043 5525
rect 29546 5516 29552 5568
rect 29604 5556 29610 5568
rect 29733 5559 29791 5565
rect 29733 5556 29745 5559
rect 29604 5528 29745 5556
rect 29604 5516 29610 5528
rect 29733 5525 29745 5528
rect 29779 5525 29791 5559
rect 29733 5519 29791 5525
rect 30650 5516 30656 5568
rect 30708 5556 30714 5568
rect 30760 5556 30788 5596
rect 31478 5584 31484 5636
rect 31536 5624 31542 5636
rect 31757 5627 31815 5633
rect 31757 5624 31769 5627
rect 31536 5596 31769 5624
rect 31536 5584 31542 5596
rect 31757 5593 31769 5596
rect 31803 5624 31815 5627
rect 32217 5627 32275 5633
rect 32217 5624 32229 5627
rect 31803 5596 32229 5624
rect 31803 5593 31815 5596
rect 31757 5587 31815 5593
rect 32217 5593 32229 5596
rect 32263 5593 32275 5627
rect 32217 5587 32275 5593
rect 35894 5584 35900 5636
rect 35952 5624 35958 5636
rect 36096 5624 36124 5655
rect 35952 5596 36124 5624
rect 36556 5624 36584 5859
rect 37093 5627 37151 5633
rect 37093 5624 37105 5627
rect 36556 5596 37105 5624
rect 35952 5584 35958 5596
rect 30926 5556 30932 5568
rect 30708 5528 30788 5556
rect 30887 5528 30932 5556
rect 30708 5516 30714 5528
rect 30926 5516 30932 5528
rect 30984 5516 30990 5568
rect 36096 5556 36124 5596
rect 37093 5593 37105 5596
rect 37139 5593 37151 5627
rect 37093 5587 37151 5593
rect 37366 5556 37372 5568
rect 36096 5528 37372 5556
rect 37366 5516 37372 5528
rect 37424 5556 37430 5568
rect 38286 5556 38292 5568
rect 37424 5528 38292 5556
rect 37424 5516 37430 5528
rect 38286 5516 38292 5528
rect 38344 5556 38350 5568
rect 38381 5559 38439 5565
rect 38381 5556 38393 5559
rect 38344 5528 38393 5556
rect 38344 5516 38350 5528
rect 38381 5525 38393 5528
rect 38427 5525 38439 5559
rect 38381 5519 38439 5525
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 3605 5355 3663 5361
rect 3605 5321 3617 5355
rect 3651 5352 3663 5355
rect 3786 5352 3792 5364
rect 3651 5324 3792 5352
rect 3651 5321 3663 5324
rect 3605 5315 3663 5321
rect 3786 5312 3792 5324
rect 3844 5312 3850 5364
rect 5074 5312 5080 5364
rect 5132 5352 5138 5364
rect 6549 5355 6607 5361
rect 6549 5352 6561 5355
rect 5132 5324 6561 5352
rect 5132 5312 5138 5324
rect 6549 5321 6561 5324
rect 6595 5321 6607 5355
rect 8846 5352 8852 5364
rect 6549 5315 6607 5321
rect 6656 5324 8852 5352
rect 1765 5287 1823 5293
rect 1765 5253 1777 5287
rect 1811 5284 1823 5287
rect 5166 5284 5172 5296
rect 1811 5256 5172 5284
rect 1811 5253 1823 5256
rect 1765 5247 1823 5253
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5216 2283 5219
rect 2314 5216 2320 5228
rect 2271 5188 2320 5216
rect 2271 5185 2283 5188
rect 2225 5179 2283 5185
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 2498 5225 2504 5228
rect 2492 5216 2504 5225
rect 2459 5188 2504 5216
rect 2492 5179 2504 5188
rect 2498 5176 2504 5179
rect 2556 5176 2562 5228
rect 4172 5225 4200 5256
rect 5166 5244 5172 5256
rect 5224 5244 5230 5296
rect 6362 5284 6368 5296
rect 6323 5256 6368 5284
rect 6362 5244 6368 5256
rect 6420 5244 6426 5296
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5185 4215 5219
rect 4157 5179 4215 5185
rect 4801 5219 4859 5225
rect 4801 5185 4813 5219
rect 4847 5216 4859 5219
rect 4890 5216 4896 5228
rect 4847 5188 4896 5216
rect 4847 5185 4859 5188
rect 4801 5179 4859 5185
rect 4890 5176 4896 5188
rect 4948 5216 4954 5228
rect 5350 5216 5356 5228
rect 4948 5188 5356 5216
rect 4948 5176 4954 5188
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 5537 5219 5595 5225
rect 5537 5185 5549 5219
rect 5583 5185 5595 5219
rect 5537 5179 5595 5185
rect 3786 5108 3792 5160
rect 3844 5148 3850 5160
rect 5552 5148 5580 5179
rect 5994 5176 6000 5228
rect 6052 5216 6058 5228
rect 6656 5216 6684 5324
rect 8846 5312 8852 5324
rect 8904 5312 8910 5364
rect 9214 5352 9220 5364
rect 9175 5324 9220 5352
rect 9214 5312 9220 5324
rect 9272 5312 9278 5364
rect 12253 5355 12311 5361
rect 12253 5321 12265 5355
rect 12299 5352 12311 5355
rect 14182 5352 14188 5364
rect 12299 5324 14188 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 14182 5312 14188 5324
rect 14240 5312 14246 5364
rect 14550 5352 14556 5364
rect 14511 5324 14556 5352
rect 14550 5312 14556 5324
rect 14608 5312 14614 5364
rect 15378 5352 15384 5364
rect 14936 5324 15384 5352
rect 6730 5244 6736 5296
rect 6788 5284 6794 5296
rect 7101 5287 7159 5293
rect 7101 5284 7113 5287
rect 6788 5256 7113 5284
rect 6788 5244 6794 5256
rect 7101 5253 7113 5256
rect 7147 5253 7159 5287
rect 8757 5287 8815 5293
rect 8757 5284 8769 5287
rect 7101 5247 7159 5253
rect 7668 5256 8769 5284
rect 7668 5228 7696 5256
rect 8757 5253 8769 5256
rect 8803 5253 8815 5287
rect 8757 5247 8815 5253
rect 6052 5188 6684 5216
rect 6052 5176 6058 5188
rect 7006 5176 7012 5228
rect 7064 5216 7070 5228
rect 7650 5216 7656 5228
rect 7064 5188 7656 5216
rect 7064 5176 7070 5188
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 7834 5176 7840 5228
rect 7892 5216 7898 5228
rect 8113 5219 8171 5225
rect 8113 5216 8125 5219
rect 7892 5188 8125 5216
rect 7892 5176 7898 5188
rect 8113 5185 8125 5188
rect 8159 5216 8171 5219
rect 9033 5219 9091 5225
rect 9033 5216 9045 5219
rect 8159 5188 9045 5216
rect 8159 5185 8171 5188
rect 8113 5179 8171 5185
rect 9033 5185 9045 5188
rect 9079 5185 9091 5219
rect 9033 5179 9091 5185
rect 11422 5176 11428 5228
rect 11480 5216 11486 5228
rect 11701 5219 11759 5225
rect 11701 5216 11713 5219
rect 11480 5188 11713 5216
rect 11480 5176 11486 5188
rect 11701 5185 11713 5188
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 12069 5219 12127 5225
rect 12069 5185 12081 5219
rect 12115 5185 12127 5219
rect 12069 5179 12127 5185
rect 3844 5120 5580 5148
rect 3844 5108 3850 5120
rect 6546 5108 6552 5160
rect 6604 5148 6610 5160
rect 6641 5151 6699 5157
rect 6641 5148 6653 5151
rect 6604 5120 6653 5148
rect 6604 5108 6610 5120
rect 6641 5117 6653 5120
rect 6687 5117 6699 5151
rect 7929 5151 7987 5157
rect 7929 5148 7941 5151
rect 6641 5111 6699 5117
rect 7116 5120 7941 5148
rect 6270 5040 6276 5092
rect 6328 5080 6334 5092
rect 7116 5089 7144 5120
rect 7929 5117 7941 5120
rect 7975 5148 7987 5151
rect 8849 5151 8907 5157
rect 8849 5148 8861 5151
rect 7975 5120 8861 5148
rect 7975 5117 7987 5120
rect 7929 5111 7987 5117
rect 8849 5117 8861 5120
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 11609 5151 11667 5157
rect 11609 5117 11621 5151
rect 11655 5148 11667 5151
rect 11790 5148 11796 5160
rect 11655 5120 11796 5148
rect 11655 5117 11667 5120
rect 11609 5111 11667 5117
rect 11790 5108 11796 5120
rect 11848 5108 11854 5160
rect 7101 5083 7159 5089
rect 7101 5080 7113 5083
rect 6328 5052 7113 5080
rect 6328 5040 6334 5052
rect 7101 5049 7113 5052
rect 7147 5049 7159 5083
rect 7101 5043 7159 5049
rect 8297 5083 8355 5089
rect 8297 5049 8309 5083
rect 8343 5080 8355 5083
rect 10134 5080 10140 5092
rect 8343 5052 10140 5080
rect 8343 5049 8355 5052
rect 8297 5043 8355 5049
rect 10134 5040 10140 5052
rect 10192 5040 10198 5092
rect 10321 5083 10379 5089
rect 10321 5049 10333 5083
rect 10367 5080 10379 5083
rect 11146 5080 11152 5092
rect 10367 5052 11152 5080
rect 10367 5049 10379 5052
rect 10321 5043 10379 5049
rect 11146 5040 11152 5052
rect 11204 5040 11210 5092
rect 11698 5040 11704 5092
rect 11756 5080 11762 5092
rect 12084 5080 12112 5179
rect 13998 5176 14004 5228
rect 14056 5216 14062 5228
rect 14936 5225 14964 5324
rect 15378 5312 15384 5324
rect 15436 5312 15442 5364
rect 16574 5312 16580 5364
rect 16632 5352 16638 5364
rect 16761 5355 16819 5361
rect 16761 5352 16773 5355
rect 16632 5324 16773 5352
rect 16632 5312 16638 5324
rect 16761 5321 16773 5324
rect 16807 5321 16819 5355
rect 16761 5315 16819 5321
rect 24765 5355 24823 5361
rect 24765 5321 24777 5355
rect 24811 5352 24823 5355
rect 24854 5352 24860 5364
rect 24811 5324 24860 5352
rect 24811 5321 24823 5324
rect 24765 5315 24823 5321
rect 24854 5312 24860 5324
rect 24912 5312 24918 5364
rect 30558 5352 30564 5364
rect 30484 5324 30564 5352
rect 15562 5284 15568 5296
rect 15028 5256 15568 5284
rect 15028 5225 15056 5256
rect 15562 5244 15568 5256
rect 15620 5244 15626 5296
rect 17034 5244 17040 5296
rect 17092 5284 17098 5296
rect 17129 5287 17187 5293
rect 17129 5284 17141 5287
rect 17092 5256 17141 5284
rect 17092 5244 17098 5256
rect 17129 5253 17141 5256
rect 17175 5253 17187 5287
rect 19334 5284 19340 5296
rect 17129 5247 17187 5253
rect 18432 5256 19340 5284
rect 14829 5219 14887 5225
rect 14829 5216 14841 5219
rect 14056 5188 14841 5216
rect 14056 5176 14062 5188
rect 14829 5185 14841 5188
rect 14875 5185 14887 5219
rect 14829 5179 14887 5185
rect 14921 5219 14979 5225
rect 14921 5185 14933 5219
rect 14967 5185 14979 5219
rect 14921 5179 14979 5185
rect 15013 5219 15071 5225
rect 15013 5185 15025 5219
rect 15059 5185 15071 5219
rect 15013 5179 15071 5185
rect 15197 5219 15255 5225
rect 15197 5185 15209 5219
rect 15243 5216 15255 5219
rect 16758 5216 16764 5228
rect 15243 5188 16764 5216
rect 15243 5185 15255 5188
rect 15197 5179 15255 5185
rect 16758 5176 16764 5188
rect 16816 5176 16822 5228
rect 16945 5219 17003 5225
rect 16945 5185 16957 5219
rect 16991 5216 17003 5219
rect 17586 5216 17592 5228
rect 16991 5188 17592 5216
rect 16991 5185 17003 5188
rect 16945 5179 17003 5185
rect 17586 5176 17592 5188
rect 17644 5176 17650 5228
rect 17862 5176 17868 5228
rect 17920 5216 17926 5228
rect 18432 5225 18460 5256
rect 19334 5244 19340 5256
rect 19392 5244 19398 5296
rect 20070 5244 20076 5296
rect 20128 5284 20134 5296
rect 21542 5284 21548 5296
rect 20128 5256 21548 5284
rect 20128 5244 20134 5256
rect 21542 5244 21548 5256
rect 21600 5244 21606 5296
rect 24578 5284 24584 5296
rect 24539 5256 24584 5284
rect 24578 5244 24584 5256
rect 24636 5244 24642 5296
rect 26234 5244 26240 5296
rect 26292 5284 26298 5296
rect 30484 5284 30512 5324
rect 30558 5312 30564 5324
rect 30616 5312 30622 5364
rect 38746 5352 38752 5364
rect 38707 5324 38752 5352
rect 38746 5312 38752 5324
rect 38804 5312 38810 5364
rect 26292 5256 30512 5284
rect 26292 5244 26298 5256
rect 18233 5219 18291 5225
rect 18233 5216 18245 5219
rect 17920 5188 18245 5216
rect 17920 5176 17926 5188
rect 18233 5185 18245 5188
rect 18279 5185 18291 5219
rect 18233 5179 18291 5185
rect 18417 5219 18475 5225
rect 18417 5185 18429 5219
rect 18463 5185 18475 5219
rect 18417 5179 18475 5185
rect 18506 5176 18512 5228
rect 18564 5216 18570 5228
rect 18647 5219 18705 5225
rect 18564 5188 18609 5216
rect 18564 5176 18570 5188
rect 18647 5185 18659 5219
rect 18693 5216 18705 5219
rect 18782 5216 18788 5228
rect 18693 5188 18788 5216
rect 18693 5185 18705 5188
rect 18647 5179 18705 5185
rect 18782 5176 18788 5188
rect 18840 5176 18846 5228
rect 24397 5219 24455 5225
rect 24397 5185 24409 5219
rect 24443 5216 24455 5219
rect 25314 5216 25320 5228
rect 24443 5188 25320 5216
rect 24443 5185 24455 5188
rect 24397 5179 24455 5185
rect 25314 5176 25320 5188
rect 25372 5176 25378 5228
rect 26326 5176 26332 5228
rect 26384 5216 26390 5228
rect 26510 5216 26516 5228
rect 26384 5188 26516 5216
rect 26384 5176 26390 5188
rect 26510 5176 26516 5188
rect 26568 5216 26574 5228
rect 27632 5225 27660 5256
rect 27525 5219 27583 5225
rect 27525 5216 27537 5219
rect 26568 5188 27537 5216
rect 26568 5176 26574 5188
rect 27525 5185 27537 5188
rect 27571 5185 27583 5219
rect 27525 5179 27583 5185
rect 27617 5219 27675 5225
rect 27617 5185 27629 5219
rect 27663 5185 27675 5219
rect 27617 5179 27675 5185
rect 27709 5219 27767 5225
rect 27709 5185 27721 5219
rect 27755 5216 27767 5219
rect 27798 5216 27804 5228
rect 27755 5188 27804 5216
rect 27755 5185 27767 5188
rect 27709 5179 27767 5185
rect 27798 5176 27804 5188
rect 27856 5176 27862 5228
rect 27893 5219 27951 5225
rect 27893 5185 27905 5219
rect 27939 5216 27951 5219
rect 27982 5216 27988 5228
rect 27939 5188 27988 5216
rect 27939 5185 27951 5188
rect 27893 5179 27951 5185
rect 27982 5176 27988 5188
rect 28040 5216 28046 5228
rect 30190 5216 30196 5228
rect 28040 5188 30196 5216
rect 28040 5176 28046 5188
rect 30190 5176 30196 5188
rect 30248 5176 30254 5228
rect 30282 5176 30288 5228
rect 30340 5216 30346 5228
rect 30484 5225 30512 5256
rect 37274 5244 37280 5296
rect 37332 5284 37338 5296
rect 37614 5287 37672 5293
rect 37614 5284 37626 5287
rect 37332 5256 37626 5284
rect 37332 5244 37338 5256
rect 37614 5253 37626 5256
rect 37660 5253 37672 5287
rect 37614 5247 37672 5253
rect 30377 5219 30435 5225
rect 30377 5216 30389 5219
rect 30340 5188 30389 5216
rect 30340 5176 30346 5188
rect 30377 5185 30389 5188
rect 30423 5185 30435 5219
rect 30377 5179 30435 5185
rect 30469 5219 30527 5225
rect 30469 5185 30481 5219
rect 30515 5185 30527 5219
rect 30469 5179 30527 5185
rect 30561 5219 30619 5225
rect 30561 5185 30573 5219
rect 30607 5185 30619 5219
rect 37366 5216 37372 5228
rect 37327 5188 37372 5216
rect 30561 5179 30619 5185
rect 22186 5108 22192 5160
rect 22244 5148 22250 5160
rect 23017 5151 23075 5157
rect 23017 5148 23029 5151
rect 22244 5120 23029 5148
rect 22244 5108 22250 5120
rect 23017 5117 23029 5120
rect 23063 5117 23075 5151
rect 29638 5148 29644 5160
rect 29599 5120 29644 5148
rect 23017 5111 23075 5117
rect 29638 5108 29644 5120
rect 29696 5148 29702 5160
rect 30576 5148 30604 5179
rect 37366 5176 37372 5188
rect 37424 5176 37430 5228
rect 29696 5120 30604 5148
rect 29696 5108 29702 5120
rect 53742 5108 53748 5160
rect 53800 5148 53806 5160
rect 54389 5151 54447 5157
rect 54389 5148 54401 5151
rect 53800 5120 54401 5148
rect 53800 5108 53806 5120
rect 54389 5117 54401 5120
rect 54435 5117 54447 5151
rect 54389 5111 54447 5117
rect 11756 5052 12112 5080
rect 11756 5040 11762 5052
rect 22646 5040 22652 5092
rect 22704 5080 22710 5092
rect 23569 5083 23627 5089
rect 23569 5080 23581 5083
rect 22704 5052 23581 5080
rect 22704 5040 22710 5052
rect 23569 5049 23581 5052
rect 23615 5049 23627 5083
rect 23569 5043 23627 5049
rect 54110 5040 54116 5092
rect 54168 5080 54174 5092
rect 55033 5083 55091 5089
rect 55033 5080 55045 5083
rect 54168 5052 55045 5080
rect 54168 5040 54174 5052
rect 55033 5049 55045 5052
rect 55079 5049 55091 5083
rect 55033 5043 55091 5049
rect 4341 5015 4399 5021
rect 4341 4981 4353 5015
rect 4387 5012 4399 5015
rect 4890 5012 4896 5024
rect 4387 4984 4896 5012
rect 4387 4981 4399 4984
rect 4341 4975 4399 4981
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 4982 4972 4988 5024
rect 5040 5012 5046 5024
rect 5718 5012 5724 5024
rect 5040 4984 5085 5012
rect 5679 4984 5724 5012
rect 5040 4972 5046 4984
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 6454 4972 6460 5024
rect 6512 5012 6518 5024
rect 7742 5012 7748 5024
rect 6512 4984 7748 5012
rect 6512 4972 6518 4984
rect 7742 4972 7748 4984
rect 7800 4972 7806 5024
rect 8018 5012 8024 5024
rect 7979 4984 8024 5012
rect 8018 4972 8024 4984
rect 8076 5012 8082 5024
rect 8757 5015 8815 5021
rect 8757 5012 8769 5015
rect 8076 4984 8769 5012
rect 8076 4972 8082 4984
rect 8757 4981 8769 4984
rect 8803 4981 8815 5015
rect 8757 4975 8815 4981
rect 10965 5015 11023 5021
rect 10965 4981 10977 5015
rect 11011 5012 11023 5015
rect 11606 5012 11612 5024
rect 11011 4984 11612 5012
rect 11011 4981 11023 4984
rect 10965 4975 11023 4981
rect 11606 4972 11612 4984
rect 11664 4972 11670 5024
rect 11974 4972 11980 5024
rect 12032 5012 12038 5024
rect 12069 5015 12127 5021
rect 12069 5012 12081 5015
rect 12032 4984 12081 5012
rect 12032 4972 12038 4984
rect 12069 4981 12081 4984
rect 12115 4981 12127 5015
rect 12069 4975 12127 4981
rect 13449 5015 13507 5021
rect 13449 4981 13461 5015
rect 13495 5012 13507 5015
rect 13538 5012 13544 5024
rect 13495 4984 13544 5012
rect 13495 4981 13507 4984
rect 13449 4975 13507 4981
rect 13538 4972 13544 4984
rect 13596 4972 13602 5024
rect 14093 5015 14151 5021
rect 14093 4981 14105 5015
rect 14139 5012 14151 5015
rect 14366 5012 14372 5024
rect 14139 4984 14372 5012
rect 14139 4981 14151 4984
rect 14093 4975 14151 4981
rect 14366 4972 14372 4984
rect 14424 4972 14430 5024
rect 15378 4972 15384 5024
rect 15436 5012 15442 5024
rect 15657 5015 15715 5021
rect 15657 5012 15669 5015
rect 15436 4984 15669 5012
rect 15436 4972 15442 4984
rect 15657 4981 15669 4984
rect 15703 4981 15715 5015
rect 17586 5012 17592 5024
rect 17547 4984 17592 5012
rect 15657 4975 15715 4981
rect 17586 4972 17592 4984
rect 17644 4972 17650 5024
rect 18874 5012 18880 5024
rect 18835 4984 18880 5012
rect 18874 4972 18880 4984
rect 18932 4972 18938 5024
rect 19334 5012 19340 5024
rect 19295 4984 19340 5012
rect 19334 4972 19340 4984
rect 19392 4972 19398 5024
rect 20070 4972 20076 5024
rect 20128 5012 20134 5024
rect 20165 5015 20223 5021
rect 20165 5012 20177 5015
rect 20128 4984 20177 5012
rect 20128 4972 20134 4984
rect 20165 4981 20177 4984
rect 20211 4981 20223 5015
rect 20165 4975 20223 4981
rect 20898 4972 20904 5024
rect 20956 5012 20962 5024
rect 20993 5015 21051 5021
rect 20993 5012 21005 5015
rect 20956 4984 21005 5012
rect 20956 4972 20962 4984
rect 20993 4981 21005 4984
rect 21039 4981 21051 5015
rect 21818 5012 21824 5024
rect 21779 4984 21824 5012
rect 20993 4975 21051 4981
rect 21818 4972 21824 4984
rect 21876 4972 21882 5024
rect 22278 4972 22284 5024
rect 22336 5012 22342 5024
rect 22373 5015 22431 5021
rect 22373 5012 22385 5015
rect 22336 4984 22385 5012
rect 22336 4972 22342 4984
rect 22373 4981 22385 4984
rect 22419 4981 22431 5015
rect 26326 5012 26332 5024
rect 26287 4984 26332 5012
rect 22373 4975 22431 4981
rect 26326 4972 26332 4984
rect 26384 4972 26390 5024
rect 27246 5012 27252 5024
rect 27207 4984 27252 5012
rect 27246 4972 27252 4984
rect 27304 4972 27310 5024
rect 30834 5012 30840 5024
rect 30795 4984 30840 5012
rect 30834 4972 30840 4984
rect 30892 4972 30898 5024
rect 53650 4972 53656 5024
rect 53708 5012 53714 5024
rect 53745 5015 53803 5021
rect 53745 5012 53757 5015
rect 53708 4984 53757 5012
rect 53708 4972 53714 4984
rect 53745 4981 53757 4984
rect 53791 4981 53803 5015
rect 58158 5012 58164 5024
rect 58119 4984 58164 5012
rect 53745 4975 53803 4981
rect 58158 4972 58164 4984
rect 58216 4972 58222 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 1949 4811 2007 4817
rect 1949 4777 1961 4811
rect 1995 4808 2007 4811
rect 5994 4808 6000 4820
rect 1995 4780 6000 4808
rect 1995 4777 2007 4780
rect 1949 4771 2007 4777
rect 5994 4768 6000 4780
rect 6052 4768 6058 4820
rect 6457 4811 6515 4817
rect 6457 4777 6469 4811
rect 6503 4808 6515 4811
rect 6730 4808 6736 4820
rect 6503 4780 6736 4808
rect 6503 4777 6515 4780
rect 6457 4771 6515 4777
rect 6730 4768 6736 4780
rect 6788 4768 6794 4820
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 7929 4811 7987 4817
rect 7929 4808 7941 4811
rect 7708 4780 7941 4808
rect 7708 4768 7714 4780
rect 7929 4777 7941 4780
rect 7975 4777 7987 4811
rect 7929 4771 7987 4777
rect 8297 4811 8355 4817
rect 8297 4777 8309 4811
rect 8343 4808 8355 4811
rect 8662 4808 8668 4820
rect 8343 4780 8668 4808
rect 8343 4777 8355 4780
rect 8297 4771 8355 4777
rect 8662 4768 8668 4780
rect 8720 4768 8726 4820
rect 9953 4811 10011 4817
rect 9953 4777 9965 4811
rect 9999 4808 10011 4811
rect 10042 4808 10048 4820
rect 9999 4780 10048 4808
rect 9999 4777 10011 4780
rect 9953 4771 10011 4777
rect 10042 4768 10048 4780
rect 10100 4768 10106 4820
rect 10318 4808 10324 4820
rect 10279 4780 10324 4808
rect 10318 4768 10324 4780
rect 10376 4768 10382 4820
rect 10962 4808 10968 4820
rect 10923 4780 10968 4808
rect 10962 4768 10968 4780
rect 11020 4768 11026 4820
rect 11698 4808 11704 4820
rect 11072 4780 11704 4808
rect 3970 4700 3976 4752
rect 4028 4740 4034 4752
rect 4525 4743 4583 4749
rect 4525 4740 4537 4743
rect 4028 4712 4537 4740
rect 4028 4700 4034 4712
rect 4525 4709 4537 4712
rect 4571 4709 4583 4743
rect 4525 4703 4583 4709
rect 5353 4743 5411 4749
rect 5353 4709 5365 4743
rect 5399 4740 5411 4743
rect 7006 4740 7012 4752
rect 5399 4712 7012 4740
rect 5399 4709 5411 4712
rect 5353 4703 5411 4709
rect 7006 4700 7012 4712
rect 7064 4700 7070 4752
rect 7742 4700 7748 4752
rect 7800 4740 7806 4752
rect 7800 4712 10088 4740
rect 7800 4700 7806 4712
rect 1762 4632 1768 4684
rect 1820 4672 1826 4684
rect 4154 4672 4160 4684
rect 1820 4644 4160 4672
rect 1820 4632 1826 4644
rect 4154 4632 4160 4644
rect 4212 4632 4218 4684
rect 5074 4632 5080 4684
rect 5132 4672 5138 4684
rect 9858 4681 9864 4684
rect 8021 4675 8079 4681
rect 8021 4672 8033 4675
rect 5132 4644 6040 4672
rect 5132 4632 5138 4644
rect 2409 4607 2467 4613
rect 2409 4573 2421 4607
rect 2455 4604 2467 4607
rect 2498 4604 2504 4616
rect 2455 4576 2504 4604
rect 2455 4573 2467 4576
rect 2409 4567 2467 4573
rect 2498 4564 2504 4576
rect 2556 4564 2562 4616
rect 3050 4604 3056 4616
rect 3011 4576 3056 4604
rect 3050 4564 3056 4576
rect 3108 4564 3114 4616
rect 3881 4607 3939 4613
rect 3881 4573 3893 4607
rect 3927 4604 3939 4607
rect 4614 4604 4620 4616
rect 3927 4576 4620 4604
rect 3927 4573 3939 4576
rect 3881 4567 3939 4573
rect 4614 4564 4620 4576
rect 4672 4604 4678 4616
rect 5258 4604 5264 4616
rect 4672 4576 5264 4604
rect 4672 4564 4678 4576
rect 5258 4564 5264 4576
rect 5316 4564 5322 4616
rect 5534 4604 5540 4616
rect 5495 4576 5540 4604
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 6012 4613 6040 4644
rect 6380 4644 8033 4672
rect 5997 4607 6055 4613
rect 5997 4573 6009 4607
rect 6043 4573 6055 4607
rect 5997 4567 6055 4573
rect 6270 4564 6276 4616
rect 6328 4604 6334 4616
rect 6380 4613 6408 4644
rect 8021 4641 8033 4644
rect 8067 4641 8079 4675
rect 8021 4635 8079 4641
rect 9824 4675 9864 4681
rect 9824 4641 9836 4675
rect 9824 4635 9864 4641
rect 9858 4632 9864 4635
rect 9916 4632 9922 4684
rect 10060 4681 10088 4712
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 11072 4672 11100 4780
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 12713 4811 12771 4817
rect 12713 4777 12725 4811
rect 12759 4808 12771 4811
rect 12759 4780 20760 4808
rect 12759 4777 12771 4780
rect 12713 4771 12771 4777
rect 11333 4743 11391 4749
rect 11333 4709 11345 4743
rect 11379 4709 11391 4743
rect 11333 4703 11391 4709
rect 11241 4675 11299 4681
rect 11241 4672 11253 4675
rect 10091 4644 11253 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 11241 4641 11253 4644
rect 11287 4641 11299 4675
rect 11348 4672 11376 4703
rect 11422 4700 11428 4752
rect 11480 4740 11486 4752
rect 15749 4743 15807 4749
rect 11480 4712 11525 4740
rect 11480 4700 11486 4712
rect 15749 4709 15761 4743
rect 15795 4740 15807 4743
rect 16482 4740 16488 4752
rect 15795 4712 16488 4740
rect 15795 4709 15807 4712
rect 15749 4703 15807 4709
rect 16482 4700 16488 4712
rect 16540 4700 16546 4752
rect 18693 4743 18751 4749
rect 18693 4709 18705 4743
rect 18739 4740 18751 4743
rect 18966 4740 18972 4752
rect 18739 4712 18972 4740
rect 18739 4709 18751 4712
rect 18693 4703 18751 4709
rect 18966 4700 18972 4712
rect 19024 4700 19030 4752
rect 20732 4740 20760 4780
rect 20806 4768 20812 4820
rect 20864 4808 20870 4820
rect 20901 4811 20959 4817
rect 20901 4808 20913 4811
rect 20864 4780 20913 4808
rect 20864 4768 20870 4780
rect 20901 4777 20913 4780
rect 20947 4777 20959 4811
rect 20901 4771 20959 4777
rect 24578 4768 24584 4820
rect 24636 4808 24642 4820
rect 25777 4811 25835 4817
rect 25777 4808 25789 4811
rect 24636 4780 25789 4808
rect 24636 4768 24642 4780
rect 25777 4777 25789 4780
rect 25823 4777 25835 4811
rect 25777 4771 25835 4777
rect 28442 4768 28448 4820
rect 28500 4808 28506 4820
rect 28537 4811 28595 4817
rect 28537 4808 28549 4811
rect 28500 4780 28549 4808
rect 28500 4768 28506 4780
rect 28537 4777 28549 4780
rect 28583 4777 28595 4811
rect 28537 4771 28595 4777
rect 32398 4768 32404 4820
rect 32456 4808 32462 4820
rect 32585 4811 32643 4817
rect 32585 4808 32597 4811
rect 32456 4780 32597 4808
rect 32456 4768 32462 4780
rect 32585 4777 32597 4780
rect 32631 4777 32643 4811
rect 32585 4771 32643 4777
rect 21726 4740 21732 4752
rect 20732 4712 21732 4740
rect 21726 4700 21732 4712
rect 21784 4700 21790 4752
rect 52178 4700 52184 4752
rect 52236 4740 52242 4752
rect 52825 4743 52883 4749
rect 52825 4740 52837 4743
rect 52236 4712 52837 4740
rect 52236 4700 52242 4712
rect 52825 4709 52837 4712
rect 52871 4709 52883 4743
rect 52825 4703 52883 4709
rect 53926 4700 53932 4752
rect 53984 4740 53990 4752
rect 55309 4743 55367 4749
rect 55309 4740 55321 4743
rect 53984 4712 55321 4740
rect 53984 4700 53990 4712
rect 55309 4709 55321 4712
rect 55355 4709 55367 4743
rect 55309 4703 55367 4709
rect 11514 4672 11520 4684
rect 11348 4644 11520 4672
rect 11241 4635 11299 4641
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 12250 4632 12256 4684
rect 12308 4672 12314 4684
rect 12308 4644 12940 4672
rect 12308 4632 12314 4644
rect 6365 4607 6423 4613
rect 6365 4604 6377 4607
rect 6328 4576 6377 4604
rect 6328 4564 6334 4576
rect 6365 4573 6377 4576
rect 6411 4573 6423 4607
rect 6638 4604 6644 4616
rect 6599 4576 6644 4604
rect 6365 4567 6423 4573
rect 6638 4564 6644 4576
rect 6696 4564 6702 4616
rect 7098 4564 7104 4616
rect 7156 4604 7162 4616
rect 7469 4607 7527 4613
rect 7469 4604 7481 4607
rect 7156 4576 7481 4604
rect 7156 4564 7162 4576
rect 7469 4573 7481 4576
rect 7515 4573 7527 4607
rect 7469 4567 7527 4573
rect 7561 4607 7619 4613
rect 7561 4573 7573 4607
rect 7607 4604 7619 4607
rect 7926 4604 7932 4616
rect 7607 4576 7932 4604
rect 7607 4573 7619 4576
rect 7561 4567 7619 4573
rect 3970 4536 3976 4548
rect 2608 4508 3976 4536
rect 2608 4477 2636 4508
rect 3970 4496 3976 4508
rect 4028 4496 4034 4548
rect 4154 4496 4160 4548
rect 4212 4536 4218 4548
rect 4709 4539 4767 4545
rect 4709 4536 4721 4539
rect 4212 4508 4721 4536
rect 4212 4496 4218 4508
rect 4709 4505 4721 4508
rect 4755 4536 4767 4539
rect 6730 4536 6736 4548
rect 4755 4508 6736 4536
rect 4755 4505 4767 4508
rect 4709 4499 4767 4505
rect 6730 4496 6736 4508
rect 6788 4496 6794 4548
rect 7484 4536 7512 4567
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 9122 4564 9128 4616
rect 9180 4604 9186 4616
rect 9217 4607 9275 4613
rect 9217 4604 9229 4607
rect 9180 4576 9229 4604
rect 9180 4564 9186 4576
rect 9217 4573 9229 4576
rect 9263 4573 9275 4607
rect 11422 4604 11428 4616
rect 9217 4567 9275 4573
rect 9692 4576 11428 4604
rect 7834 4536 7840 4548
rect 7484 4508 7840 4536
rect 7834 4496 7840 4508
rect 7892 4496 7898 4548
rect 9692 4545 9720 4576
rect 11422 4564 11428 4576
rect 11480 4564 11486 4616
rect 11790 4604 11796 4616
rect 11751 4576 11796 4604
rect 11790 4564 11796 4576
rect 11848 4564 11854 4616
rect 12912 4613 12940 4644
rect 16022 4632 16028 4684
rect 16080 4672 16086 4684
rect 19521 4675 19579 4681
rect 19521 4672 19533 4675
rect 16080 4644 19533 4672
rect 16080 4632 16086 4644
rect 19521 4641 19533 4644
rect 19567 4641 19579 4675
rect 27154 4672 27160 4684
rect 27115 4644 27160 4672
rect 19521 4635 19579 4641
rect 27154 4632 27160 4644
rect 27212 4632 27218 4684
rect 31202 4672 31208 4684
rect 31163 4644 31208 4672
rect 31202 4632 31208 4644
rect 31260 4632 31266 4684
rect 53190 4632 53196 4684
rect 53248 4672 53254 4684
rect 54113 4675 54171 4681
rect 54113 4672 54125 4675
rect 53248 4644 54125 4672
rect 53248 4632 53254 4644
rect 54113 4641 54125 4644
rect 54159 4641 54171 4675
rect 54113 4635 54171 4641
rect 54294 4632 54300 4684
rect 54352 4672 54358 4684
rect 55953 4675 56011 4681
rect 55953 4672 55965 4675
rect 54352 4644 55965 4672
rect 54352 4632 54358 4644
rect 55953 4641 55965 4644
rect 55999 4641 56011 4675
rect 55953 4635 56011 4641
rect 12713 4607 12771 4613
rect 12713 4604 12725 4607
rect 12406 4576 12725 4604
rect 9677 4539 9735 4545
rect 9677 4536 9689 4539
rect 7944 4508 9689 4536
rect 2593 4471 2651 4477
rect 2593 4437 2605 4471
rect 2639 4437 2651 4471
rect 2593 4431 2651 4437
rect 3145 4471 3203 4477
rect 3145 4437 3157 4471
rect 3191 4468 3203 4471
rect 3694 4468 3700 4480
rect 3191 4440 3700 4468
rect 3191 4437 3203 4440
rect 3145 4431 3203 4437
rect 3694 4428 3700 4440
rect 3752 4428 3758 4480
rect 4065 4471 4123 4477
rect 4065 4437 4077 4471
rect 4111 4468 4123 4471
rect 4614 4468 4620 4480
rect 4111 4440 4620 4468
rect 4111 4437 4123 4440
rect 4065 4431 4123 4437
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 6181 4471 6239 4477
rect 6181 4437 6193 4471
rect 6227 4468 6239 4471
rect 7098 4468 7104 4480
rect 6227 4440 7104 4468
rect 6227 4437 6239 4440
rect 6181 4431 6239 4437
rect 7098 4428 7104 4440
rect 7156 4428 7162 4480
rect 7282 4428 7288 4480
rect 7340 4468 7346 4480
rect 7944 4468 7972 4508
rect 9677 4505 9689 4508
rect 9723 4505 9735 4539
rect 9677 4499 9735 4505
rect 10134 4496 10140 4548
rect 10192 4536 10198 4548
rect 12406 4536 12434 4576
rect 12713 4573 12725 4576
rect 12759 4573 12771 4607
rect 12713 4567 12771 4573
rect 12897 4607 12955 4613
rect 12897 4573 12909 4607
rect 12943 4573 12955 4607
rect 12897 4567 12955 4573
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4604 13599 4607
rect 13998 4604 14004 4616
rect 13587 4576 14004 4604
rect 13587 4573 13599 4576
rect 13541 4567 13599 4573
rect 13998 4564 14004 4576
rect 14056 4564 14062 4616
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 14274 4564 14280 4576
rect 14332 4604 14338 4616
rect 14734 4604 14740 4616
rect 14332 4576 14740 4604
rect 14332 4564 14338 4576
rect 14734 4564 14740 4576
rect 14792 4564 14798 4616
rect 15105 4607 15163 4613
rect 15105 4573 15117 4607
rect 15151 4604 15163 4607
rect 15930 4604 15936 4616
rect 15151 4576 15936 4604
rect 15151 4573 15163 4576
rect 15105 4567 15163 4573
rect 15930 4564 15936 4576
rect 15988 4564 15994 4616
rect 16393 4607 16451 4613
rect 16393 4573 16405 4607
rect 16439 4573 16451 4607
rect 16393 4567 16451 4573
rect 10192 4508 12434 4536
rect 16408 4536 16436 4567
rect 16758 4564 16764 4616
rect 16816 4604 16822 4616
rect 16853 4607 16911 4613
rect 16853 4604 16865 4607
rect 16816 4576 16865 4604
rect 16816 4564 16822 4576
rect 16853 4573 16865 4576
rect 16899 4573 16911 4607
rect 16853 4567 16911 4573
rect 18049 4607 18107 4613
rect 18049 4573 18061 4607
rect 18095 4604 18107 4607
rect 18598 4604 18604 4616
rect 18095 4576 18604 4604
rect 18095 4573 18107 4576
rect 18049 4567 18107 4573
rect 18598 4564 18604 4576
rect 18656 4564 18662 4616
rect 18874 4564 18880 4616
rect 18932 4604 18938 4616
rect 19777 4607 19835 4613
rect 19777 4604 19789 4607
rect 18932 4576 19789 4604
rect 18932 4564 18938 4576
rect 19777 4573 19789 4576
rect 19823 4573 19835 4607
rect 21726 4604 21732 4616
rect 21687 4576 21732 4604
rect 19777 4567 19835 4573
rect 21726 4564 21732 4576
rect 21784 4564 21790 4616
rect 22373 4607 22431 4613
rect 22373 4573 22385 4607
rect 22419 4604 22431 4607
rect 22554 4604 22560 4616
rect 22419 4576 22560 4604
rect 22419 4573 22431 4576
rect 22373 4567 22431 4573
rect 22554 4564 22560 4576
rect 22612 4564 22618 4616
rect 23017 4607 23075 4613
rect 23017 4573 23029 4607
rect 23063 4604 23075 4607
rect 23106 4604 23112 4616
rect 23063 4576 23112 4604
rect 23063 4573 23075 4576
rect 23017 4567 23075 4573
rect 23106 4564 23112 4576
rect 23164 4564 23170 4616
rect 23474 4604 23480 4616
rect 23435 4576 23480 4604
rect 23474 4564 23480 4576
rect 23532 4564 23538 4616
rect 23934 4564 23940 4616
rect 23992 4604 23998 4616
rect 24397 4607 24455 4613
rect 24397 4604 24409 4607
rect 23992 4576 24409 4604
rect 23992 4564 23998 4576
rect 24397 4573 24409 4576
rect 24443 4604 24455 4607
rect 24946 4604 24952 4616
rect 24443 4576 24952 4604
rect 24443 4573 24455 4576
rect 24397 4567 24455 4573
rect 24946 4564 24952 4576
rect 25004 4564 25010 4616
rect 27246 4564 27252 4616
rect 27304 4604 27310 4616
rect 27413 4607 27471 4613
rect 27413 4604 27425 4607
rect 27304 4576 27425 4604
rect 27304 4564 27310 4576
rect 27413 4573 27425 4576
rect 27459 4573 27471 4607
rect 27413 4567 27471 4573
rect 30926 4564 30932 4616
rect 30984 4604 30990 4616
rect 31461 4607 31519 4613
rect 31461 4604 31473 4607
rect 30984 4576 31473 4604
rect 30984 4564 30990 4576
rect 31461 4573 31473 4576
rect 31507 4573 31519 4607
rect 31461 4567 31519 4573
rect 52086 4564 52092 4616
rect 52144 4604 52150 4616
rect 52181 4607 52239 4613
rect 52181 4604 52193 4607
rect 52144 4576 52193 4604
rect 52144 4564 52150 4576
rect 52181 4573 52193 4576
rect 52227 4573 52239 4607
rect 52181 4567 52239 4573
rect 52638 4564 52644 4616
rect 52696 4604 52702 4616
rect 53469 4607 53527 4613
rect 53469 4604 53481 4607
rect 52696 4576 53481 4604
rect 52696 4564 52702 4576
rect 53469 4573 53481 4576
rect 53515 4573 53527 4607
rect 53469 4567 53527 4573
rect 18138 4536 18144 4548
rect 16408 4508 18144 4536
rect 10192 4496 10198 4508
rect 18138 4496 18144 4508
rect 18196 4496 18202 4548
rect 24670 4545 24676 4548
rect 24664 4536 24676 4545
rect 24631 4508 24676 4536
rect 24664 4499 24676 4508
rect 24670 4496 24676 4499
rect 24728 4496 24734 4548
rect 7340 4440 7972 4468
rect 7340 4428 7346 4440
rect 8294 4428 8300 4480
rect 8352 4468 8358 4480
rect 9033 4471 9091 4477
rect 9033 4468 9045 4471
rect 8352 4440 9045 4468
rect 8352 4428 8358 4440
rect 9033 4437 9045 4440
rect 9079 4437 9091 4471
rect 9033 4431 9091 4437
rect 10042 4428 10048 4480
rect 10100 4468 10106 4480
rect 11514 4468 11520 4480
rect 10100 4440 11520 4468
rect 10100 4428 10106 4440
rect 11514 4428 11520 4440
rect 11572 4468 11578 4480
rect 11974 4468 11980 4480
rect 11572 4440 11980 4468
rect 11572 4428 11578 4440
rect 11974 4428 11980 4440
rect 12032 4428 12038 4480
rect 14461 4471 14519 4477
rect 14461 4437 14473 4471
rect 14507 4468 14519 4471
rect 14826 4468 14832 4480
rect 14507 4440 14832 4468
rect 14507 4437 14519 4440
rect 14461 4431 14519 4437
rect 14826 4428 14832 4440
rect 14884 4428 14890 4480
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 3050 4264 3056 4276
rect 3011 4236 3056 4264
rect 3050 4224 3056 4236
rect 3108 4224 3114 4276
rect 3694 4224 3700 4276
rect 3752 4264 3758 4276
rect 5534 4264 5540 4276
rect 3752 4236 5540 4264
rect 3752 4224 3758 4236
rect 5534 4224 5540 4236
rect 5592 4224 5598 4276
rect 5813 4267 5871 4273
rect 5813 4233 5825 4267
rect 5859 4264 5871 4267
rect 6270 4264 6276 4276
rect 5859 4236 6276 4264
rect 5859 4233 5871 4236
rect 5813 4227 5871 4233
rect 6270 4224 6276 4236
rect 6328 4224 6334 4276
rect 6546 4224 6552 4276
rect 6604 4273 6610 4276
rect 6604 4267 6623 4273
rect 6611 4233 6623 4267
rect 6604 4227 6623 4233
rect 6604 4224 6610 4227
rect 7098 4224 7104 4276
rect 7156 4264 7162 4276
rect 7466 4264 7472 4276
rect 7156 4236 7472 4264
rect 7156 4224 7162 4236
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 7650 4224 7656 4276
rect 7708 4264 7714 4276
rect 7708 4236 9904 4264
rect 7708 4224 7714 4236
rect 3602 4156 3608 4208
rect 3660 4196 3666 4208
rect 3660 4168 4384 4196
rect 3660 4156 3666 4168
rect 1765 4131 1823 4137
rect 1765 4097 1777 4131
rect 1811 4097 1823 4131
rect 1765 4091 1823 4097
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4128 2467 4131
rect 2682 4128 2688 4140
rect 2455 4100 2688 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 1780 4060 1808 4091
rect 2682 4088 2688 4100
rect 2740 4088 2746 4140
rect 3142 4088 3148 4140
rect 3200 4128 3206 4140
rect 3237 4131 3295 4137
rect 3237 4128 3249 4131
rect 3200 4100 3249 4128
rect 3200 4088 3206 4100
rect 3237 4097 3249 4100
rect 3283 4128 3295 4131
rect 3878 4128 3884 4140
rect 3283 4100 3884 4128
rect 3283 4097 3295 4100
rect 3237 4091 3295 4097
rect 3878 4088 3884 4100
rect 3936 4088 3942 4140
rect 4356 4137 4384 4168
rect 4890 4156 4896 4208
rect 4948 4196 4954 4208
rect 6365 4199 6423 4205
rect 6365 4196 6377 4199
rect 4948 4168 6377 4196
rect 4948 4156 4954 4168
rect 6365 4165 6377 4168
rect 6411 4165 6423 4199
rect 6365 4159 6423 4165
rect 7484 4168 8064 4196
rect 4341 4131 4399 4137
rect 4341 4097 4353 4131
rect 4387 4097 4399 4131
rect 4341 4091 4399 4097
rect 4985 4131 5043 4137
rect 4985 4097 4997 4131
rect 5031 4128 5043 4131
rect 5629 4131 5687 4137
rect 5031 4100 5580 4128
rect 5031 4097 5043 4100
rect 4985 4091 5043 4097
rect 4801 4063 4859 4069
rect 4801 4060 4813 4063
rect 1780 4032 4813 4060
rect 4801 4029 4813 4032
rect 4847 4029 4859 4063
rect 4801 4023 4859 4029
rect 4890 4020 4896 4072
rect 4948 4060 4954 4072
rect 5169 4063 5227 4069
rect 5169 4060 5181 4063
rect 4948 4032 5181 4060
rect 4948 4020 4954 4032
rect 5169 4029 5181 4032
rect 5215 4029 5227 4063
rect 5552 4060 5580 4100
rect 5629 4097 5641 4131
rect 5675 4128 5687 4131
rect 7484 4128 7512 4168
rect 5675 4100 7512 4128
rect 7561 4131 7619 4137
rect 5675 4097 5687 4100
rect 5629 4091 5687 4097
rect 7561 4097 7573 4131
rect 7607 4128 7619 4131
rect 7926 4128 7932 4140
rect 7607 4100 7932 4128
rect 7607 4097 7619 4100
rect 7561 4091 7619 4097
rect 7926 4088 7932 4100
rect 7984 4088 7990 4140
rect 8036 4128 8064 4168
rect 8036 4100 8156 4128
rect 5810 4060 5816 4072
rect 5552 4032 5816 4060
rect 5169 4023 5227 4029
rect 5810 4020 5816 4032
rect 5868 4060 5874 4072
rect 6546 4060 6552 4072
rect 5868 4032 6552 4060
rect 5868 4020 5874 4032
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 7466 4060 7472 4072
rect 7427 4032 7472 4060
rect 7466 4020 7472 4032
rect 7524 4020 7530 4072
rect 7834 4020 7840 4072
rect 7892 4060 7898 4072
rect 8021 4063 8079 4069
rect 8021 4060 8033 4063
rect 7892 4032 8033 4060
rect 7892 4020 7898 4032
rect 8021 4029 8033 4032
rect 8067 4029 8079 4063
rect 8021 4023 8079 4029
rect 2593 3995 2651 4001
rect 2593 3961 2605 3995
rect 2639 3992 2651 3995
rect 3694 3992 3700 4004
rect 2639 3964 3700 3992
rect 2639 3961 2651 3964
rect 2593 3955 2651 3961
rect 3694 3952 3700 3964
rect 3752 3952 3758 4004
rect 3970 3952 3976 4004
rect 4028 3992 4034 4004
rect 4028 3964 6592 3992
rect 4028 3952 4034 3964
rect 1946 3924 1952 3936
rect 1907 3896 1952 3924
rect 1946 3884 1952 3896
rect 2004 3884 2010 3936
rect 4157 3927 4215 3933
rect 4157 3893 4169 3927
rect 4203 3924 4215 3927
rect 6454 3924 6460 3936
rect 4203 3896 6460 3924
rect 4203 3893 4215 3896
rect 4157 3887 4215 3893
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 6564 3933 6592 3964
rect 6914 3952 6920 4004
rect 6972 3992 6978 4004
rect 7193 3995 7251 4001
rect 7193 3992 7205 3995
rect 6972 3964 7205 3992
rect 6972 3952 6978 3964
rect 7193 3961 7205 3964
rect 7239 3961 7251 3995
rect 7193 3955 7251 3961
rect 6549 3927 6607 3933
rect 6549 3893 6561 3927
rect 6595 3893 6607 3927
rect 6549 3887 6607 3893
rect 6733 3927 6791 3933
rect 6733 3893 6745 3927
rect 6779 3924 6791 3927
rect 7098 3924 7104 3936
rect 6779 3896 7104 3924
rect 6779 3893 6791 3896
rect 6733 3887 6791 3893
rect 7098 3884 7104 3896
rect 7156 3884 7162 3936
rect 7561 3927 7619 3933
rect 7561 3893 7573 3927
rect 7607 3924 7619 3927
rect 7852 3924 7880 4020
rect 7607 3896 7880 3924
rect 8128 3924 8156 4100
rect 9306 4088 9312 4140
rect 9364 4128 9370 4140
rect 9677 4131 9735 4137
rect 9677 4128 9689 4131
rect 9364 4100 9689 4128
rect 9364 4088 9370 4100
rect 9677 4097 9689 4100
rect 9723 4128 9735 4131
rect 9766 4128 9772 4140
rect 9723 4100 9772 4128
rect 9723 4097 9735 4100
rect 9677 4091 9735 4097
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 9876 4128 9904 4236
rect 15562 4224 15568 4276
rect 15620 4264 15626 4276
rect 15838 4264 15844 4276
rect 15620 4236 15844 4264
rect 15620 4224 15626 4236
rect 15838 4224 15844 4236
rect 15896 4224 15902 4276
rect 14476 4168 15700 4196
rect 10965 4131 11023 4137
rect 10965 4128 10977 4131
rect 9876 4100 10977 4128
rect 10965 4097 10977 4100
rect 11011 4097 11023 4131
rect 14476 4128 14504 4168
rect 15672 4137 15700 4168
rect 22094 4156 22100 4208
rect 22152 4196 22158 4208
rect 25133 4199 25191 4205
rect 25133 4196 25145 4199
rect 22152 4168 25145 4196
rect 22152 4156 22158 4168
rect 25133 4165 25145 4168
rect 25179 4165 25191 4199
rect 35894 4196 35900 4208
rect 25133 4159 25191 4165
rect 35360 4168 35900 4196
rect 10965 4091 11023 4097
rect 11256 4100 14504 4128
rect 14553 4131 14611 4137
rect 8478 4060 8484 4072
rect 8404 4032 8484 4060
rect 8404 4001 8432 4032
rect 8478 4020 8484 4032
rect 8536 4020 8542 4072
rect 8573 4063 8631 4069
rect 8573 4029 8585 4063
rect 8619 4029 8631 4063
rect 8573 4023 8631 4029
rect 8389 3995 8447 4001
rect 8389 3961 8401 3995
rect 8435 3961 8447 3995
rect 8588 3992 8616 4023
rect 8662 4020 8668 4072
rect 8720 4060 8726 4072
rect 10229 4063 10287 4069
rect 8720 4032 8765 4060
rect 8720 4020 8726 4032
rect 10229 4029 10241 4063
rect 10275 4060 10287 4063
rect 11256 4060 11284 4100
rect 14553 4097 14565 4131
rect 14599 4128 14611 4131
rect 15657 4131 15715 4137
rect 14599 4100 15608 4128
rect 14599 4097 14611 4100
rect 14553 4091 14611 4097
rect 10275 4032 11284 4060
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 11422 4020 11428 4072
rect 11480 4060 11486 4072
rect 11517 4063 11575 4069
rect 11517 4060 11529 4063
rect 11480 4032 11529 4060
rect 11480 4020 11486 4032
rect 11517 4029 11529 4032
rect 11563 4029 11575 4063
rect 11517 4023 11575 4029
rect 11698 4020 11704 4072
rect 11756 4060 11762 4072
rect 12069 4063 12127 4069
rect 12069 4060 12081 4063
rect 11756 4032 12081 4060
rect 11756 4020 11762 4032
rect 12069 4029 12081 4032
rect 12115 4029 12127 4063
rect 12069 4023 12127 4029
rect 12345 4063 12403 4069
rect 12345 4029 12357 4063
rect 12391 4060 12403 4063
rect 12894 4060 12900 4072
rect 12391 4032 12900 4060
rect 12391 4029 12403 4032
rect 12345 4023 12403 4029
rect 12894 4020 12900 4032
rect 12952 4020 12958 4072
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4060 13323 4063
rect 14642 4060 14648 4072
rect 13311 4032 14648 4060
rect 13311 4029 13323 4032
rect 13265 4023 13323 4029
rect 14642 4020 14648 4032
rect 14700 4020 14706 4072
rect 15580 4060 15608 4100
rect 15657 4097 15669 4131
rect 15703 4128 15715 4131
rect 15746 4128 15752 4140
rect 15703 4100 15752 4128
rect 15703 4097 15715 4100
rect 15657 4091 15715 4097
rect 15746 4088 15752 4100
rect 15804 4088 15810 4140
rect 16666 4088 16672 4140
rect 16724 4128 16730 4140
rect 17218 4128 17224 4140
rect 16724 4100 17224 4128
rect 16724 4088 16730 4100
rect 17218 4088 17224 4100
rect 17276 4128 17282 4140
rect 17313 4131 17371 4137
rect 17313 4128 17325 4131
rect 17276 4100 17325 4128
rect 17276 4088 17282 4100
rect 17313 4097 17325 4100
rect 17359 4097 17371 4131
rect 17313 4091 17371 4097
rect 22916 4131 22974 4137
rect 22916 4097 22928 4131
rect 22962 4128 22974 4131
rect 23198 4128 23204 4140
rect 22962 4100 23204 4128
rect 22962 4097 22974 4100
rect 22916 4091 22974 4097
rect 23198 4088 23204 4100
rect 23256 4088 23262 4140
rect 35161 4131 35219 4137
rect 35161 4097 35173 4131
rect 35207 4128 35219 4131
rect 35360 4128 35388 4168
rect 35894 4156 35900 4168
rect 35952 4156 35958 4208
rect 35434 4137 35440 4140
rect 35207 4100 35388 4128
rect 35207 4097 35219 4100
rect 35161 4091 35219 4097
rect 35428 4091 35440 4137
rect 35492 4128 35498 4140
rect 35492 4100 35528 4128
rect 35434 4088 35440 4091
rect 35492 4088 35498 4100
rect 53006 4088 53012 4140
rect 53064 4128 53070 4140
rect 54665 4131 54723 4137
rect 54665 4128 54677 4131
rect 53064 4100 54677 4128
rect 53064 4088 53070 4100
rect 54665 4097 54677 4100
rect 54711 4097 54723 4131
rect 54665 4091 54723 4097
rect 17862 4060 17868 4072
rect 15580 4032 17868 4060
rect 17862 4020 17868 4032
rect 17920 4020 17926 4072
rect 22649 4063 22707 4069
rect 22649 4029 22661 4063
rect 22695 4029 22707 4063
rect 22649 4023 22707 4029
rect 8754 3992 8760 4004
rect 8588 3964 8760 3992
rect 8389 3955 8447 3961
rect 8754 3952 8760 3964
rect 8812 3952 8818 4004
rect 9490 3992 9496 4004
rect 9451 3964 9496 3992
rect 9490 3952 9496 3964
rect 9548 3952 9554 4004
rect 9858 3952 9864 4004
rect 9916 3992 9922 4004
rect 11974 3992 11980 4004
rect 9916 3964 11744 3992
rect 11935 3964 11980 3992
rect 9916 3952 9922 3964
rect 8481 3927 8539 3933
rect 8481 3924 8493 3927
rect 8128 3896 8493 3924
rect 7607 3893 7619 3896
rect 7561 3887 7619 3893
rect 8481 3893 8493 3896
rect 8527 3924 8539 3927
rect 8938 3924 8944 3936
rect 8527 3896 8944 3924
rect 8527 3893 8539 3896
rect 8481 3887 8539 3893
rect 8938 3884 8944 3896
rect 8996 3924 9002 3936
rect 9214 3924 9220 3936
rect 8996 3896 9220 3924
rect 8996 3884 9002 3896
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 10594 3884 10600 3936
rect 10652 3924 10658 3936
rect 10781 3927 10839 3933
rect 10781 3924 10793 3927
rect 10652 3896 10793 3924
rect 10652 3884 10658 3896
rect 10781 3893 10793 3896
rect 10827 3893 10839 3927
rect 11716 3924 11744 3964
rect 11974 3952 11980 3964
rect 12032 3952 12038 4004
rect 13909 3995 13967 4001
rect 13909 3961 13921 3995
rect 13955 3992 13967 3995
rect 15286 3992 15292 4004
rect 13955 3964 15292 3992
rect 13955 3961 13967 3964
rect 13909 3955 13967 3961
rect 15286 3952 15292 3964
rect 15344 3952 15350 4004
rect 15838 3992 15844 4004
rect 15799 3964 15844 3992
rect 15838 3952 15844 3964
rect 15896 3952 15902 4004
rect 18693 3995 18751 4001
rect 18693 3961 18705 3995
rect 18739 3992 18751 3995
rect 19426 3992 19432 4004
rect 18739 3964 19432 3992
rect 18739 3961 18751 3964
rect 18693 3955 18751 3961
rect 19426 3952 19432 3964
rect 19484 3952 19490 4004
rect 20625 3995 20683 4001
rect 20625 3961 20637 3995
rect 20671 3992 20683 3995
rect 21450 3992 21456 4004
rect 20671 3964 21456 3992
rect 20671 3961 20683 3964
rect 20625 3955 20683 3961
rect 21450 3952 21456 3964
rect 21508 3952 21514 4004
rect 11790 3924 11796 3936
rect 11703 3896 11796 3924
rect 10781 3887 10839 3893
rect 11790 3884 11796 3896
rect 11848 3924 11854 3936
rect 11885 3927 11943 3933
rect 11885 3924 11897 3927
rect 11848 3896 11897 3924
rect 11848 3884 11854 3896
rect 11885 3893 11897 3896
rect 11931 3893 11943 3927
rect 11885 3887 11943 3893
rect 15197 3927 15255 3933
rect 15197 3893 15209 3927
rect 15243 3924 15255 3927
rect 16298 3924 16304 3936
rect 15243 3896 16304 3924
rect 15243 3893 15255 3896
rect 15197 3887 15255 3893
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 16853 3927 16911 3933
rect 16853 3893 16865 3927
rect 16899 3924 16911 3927
rect 17310 3924 17316 3936
rect 16899 3896 17316 3924
rect 16899 3893 16911 3896
rect 16853 3887 16911 3893
rect 17310 3884 17316 3896
rect 17368 3884 17374 3936
rect 17497 3927 17555 3933
rect 17497 3893 17509 3927
rect 17543 3924 17555 3927
rect 18782 3924 18788 3936
rect 17543 3896 18788 3924
rect 17543 3893 17555 3896
rect 17497 3887 17555 3893
rect 18782 3884 18788 3896
rect 18840 3884 18846 3936
rect 19337 3927 19395 3933
rect 19337 3893 19349 3927
rect 19383 3924 19395 3927
rect 19702 3924 19708 3936
rect 19383 3896 19708 3924
rect 19383 3893 19395 3896
rect 19337 3887 19395 3893
rect 19702 3884 19708 3896
rect 19760 3884 19766 3936
rect 19981 3927 20039 3933
rect 19981 3893 19993 3927
rect 20027 3924 20039 3927
rect 20346 3924 20352 3936
rect 20027 3896 20352 3924
rect 20027 3893 20039 3896
rect 19981 3887 20039 3893
rect 20346 3884 20352 3896
rect 20404 3884 20410 3936
rect 21269 3927 21327 3933
rect 21269 3893 21281 3927
rect 21315 3924 21327 3927
rect 22002 3924 22008 3936
rect 21315 3896 22008 3924
rect 21315 3893 21327 3896
rect 21269 3887 21327 3893
rect 22002 3884 22008 3896
rect 22060 3884 22066 3936
rect 22189 3927 22247 3933
rect 22189 3893 22201 3927
rect 22235 3924 22247 3927
rect 22462 3924 22468 3936
rect 22235 3896 22468 3924
rect 22235 3893 22247 3896
rect 22189 3887 22247 3893
rect 22462 3884 22468 3896
rect 22520 3884 22526 3936
rect 22664 3924 22692 4023
rect 24026 4020 24032 4072
rect 24084 4060 24090 4072
rect 24489 4063 24547 4069
rect 24489 4060 24501 4063
rect 24084 4032 24501 4060
rect 24084 4020 24090 4032
rect 24489 4029 24501 4032
rect 24535 4029 24547 4063
rect 24489 4023 24547 4029
rect 51810 4020 51816 4072
rect 51868 4060 51874 4072
rect 52733 4063 52791 4069
rect 52733 4060 52745 4063
rect 51868 4032 52745 4060
rect 51868 4020 51874 4032
rect 52733 4029 52745 4032
rect 52779 4029 52791 4063
rect 52733 4023 52791 4029
rect 54018 4020 54024 4072
rect 54076 4060 54082 4072
rect 55953 4063 56011 4069
rect 55953 4060 55965 4063
rect 54076 4032 55965 4060
rect 54076 4020 54082 4032
rect 55953 4029 55965 4032
rect 55999 4029 56011 4063
rect 55953 4023 56011 4029
rect 24762 3992 24768 4004
rect 24044 3964 24768 3992
rect 23934 3924 23940 3936
rect 22664 3896 23940 3924
rect 23934 3884 23940 3896
rect 23992 3884 23998 3936
rect 24044 3933 24072 3964
rect 24762 3952 24768 3964
rect 24820 3952 24826 4004
rect 36170 3952 36176 4004
rect 36228 3992 36234 4004
rect 36541 3995 36599 4001
rect 36541 3992 36553 3995
rect 36228 3964 36553 3992
rect 36228 3952 36234 3964
rect 36541 3961 36553 3964
rect 36587 3961 36599 3995
rect 36541 3955 36599 3961
rect 52822 3952 52828 4004
rect 52880 3992 52886 4004
rect 52880 3964 54064 3992
rect 52880 3952 52886 3964
rect 24029 3927 24087 3933
rect 24029 3893 24041 3927
rect 24075 3893 24087 3927
rect 25682 3924 25688 3936
rect 25643 3896 25688 3924
rect 24029 3887 24087 3893
rect 25682 3884 25688 3896
rect 25740 3884 25746 3936
rect 26234 3924 26240 3936
rect 26195 3896 26240 3924
rect 26234 3884 26240 3896
rect 26292 3884 26298 3936
rect 51074 3884 51080 3936
rect 51132 3924 51138 3936
rect 51169 3927 51227 3933
rect 51169 3924 51181 3927
rect 51132 3896 51181 3924
rect 51132 3884 51138 3896
rect 51169 3893 51181 3896
rect 51215 3893 51227 3927
rect 51169 3887 51227 3893
rect 51350 3884 51356 3936
rect 51408 3924 51414 3936
rect 51813 3927 51871 3933
rect 51813 3924 51825 3927
rect 51408 3896 51825 3924
rect 51408 3884 51414 3896
rect 51813 3893 51825 3896
rect 51859 3893 51871 3927
rect 51813 3887 51871 3893
rect 52454 3884 52460 3936
rect 52512 3924 52518 3936
rect 54036 3933 54064 3964
rect 53377 3927 53435 3933
rect 53377 3924 53389 3927
rect 52512 3896 53389 3924
rect 52512 3884 52518 3896
rect 53377 3893 53389 3896
rect 53423 3893 53435 3927
rect 53377 3887 53435 3893
rect 54021 3927 54079 3933
rect 54021 3893 54033 3927
rect 54067 3893 54079 3927
rect 55306 3924 55312 3936
rect 55267 3896 55312 3924
rect 54021 3887 54079 3893
rect 55306 3884 55312 3896
rect 55364 3884 55370 3936
rect 58161 3927 58219 3933
rect 58161 3893 58173 3927
rect 58207 3924 58219 3927
rect 58434 3924 58440 3936
rect 58207 3896 58440 3924
rect 58207 3893 58219 3896
rect 58161 3887 58219 3893
rect 58434 3884 58440 3896
rect 58492 3884 58498 3936
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 3694 3680 3700 3732
rect 3752 3720 3758 3732
rect 4890 3720 4896 3732
rect 3752 3692 4896 3720
rect 3752 3680 3758 3692
rect 4890 3680 4896 3692
rect 4948 3680 4954 3732
rect 4982 3680 4988 3732
rect 5040 3720 5046 3732
rect 6270 3720 6276 3732
rect 5040 3692 6276 3720
rect 5040 3680 5046 3692
rect 6270 3680 6276 3692
rect 6328 3680 6334 3732
rect 6362 3680 6368 3732
rect 6420 3680 6426 3732
rect 7466 3680 7472 3732
rect 7524 3720 7530 3732
rect 9858 3720 9864 3732
rect 7524 3692 9864 3720
rect 7524 3680 7530 3692
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 17405 3723 17463 3729
rect 17405 3689 17417 3723
rect 17451 3720 17463 3723
rect 17678 3720 17684 3732
rect 17451 3692 17684 3720
rect 17451 3689 17463 3692
rect 17405 3683 17463 3689
rect 17678 3680 17684 3692
rect 17736 3680 17742 3732
rect 20254 3720 20260 3732
rect 20215 3692 20260 3720
rect 20254 3680 20260 3692
rect 20312 3680 20318 3732
rect 20990 3720 20996 3732
rect 20951 3692 20996 3720
rect 20990 3680 20996 3692
rect 21048 3680 21054 3732
rect 21082 3680 21088 3732
rect 21140 3720 21146 3732
rect 25682 3720 25688 3732
rect 21140 3692 25688 3720
rect 21140 3680 21146 3692
rect 25682 3680 25688 3692
rect 25740 3680 25746 3732
rect 32122 3720 32128 3732
rect 32083 3692 32128 3720
rect 32122 3680 32128 3692
rect 32180 3680 32186 3732
rect 52730 3680 52736 3732
rect 52788 3720 52794 3732
rect 52788 3692 55214 3720
rect 52788 3680 52794 3692
rect 3237 3655 3295 3661
rect 3237 3621 3249 3655
rect 3283 3621 3295 3655
rect 6380 3652 6408 3680
rect 8202 3652 8208 3664
rect 6380 3624 6868 3652
rect 8163 3624 8208 3652
rect 3237 3615 3295 3621
rect 3252 3584 3280 3615
rect 3252 3556 4384 3584
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 2406 3516 2412 3528
rect 1903 3488 2412 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 2406 3476 2412 3488
rect 2464 3516 2470 3528
rect 4249 3519 4307 3525
rect 4249 3516 4261 3519
rect 2464 3488 4261 3516
rect 2464 3476 2470 3488
rect 4249 3485 4261 3488
rect 4295 3485 4307 3519
rect 4356 3516 4384 3556
rect 6086 3544 6092 3596
rect 6144 3584 6150 3596
rect 6362 3584 6368 3596
rect 6144 3556 6368 3584
rect 6144 3544 6150 3556
rect 6362 3544 6368 3556
rect 6420 3584 6426 3596
rect 6840 3593 6868 3624
rect 8202 3612 8208 3624
rect 8260 3612 8266 3664
rect 9398 3652 9404 3664
rect 9359 3624 9404 3652
rect 9398 3612 9404 3624
rect 9456 3612 9462 3664
rect 9674 3612 9680 3664
rect 9732 3652 9738 3664
rect 11517 3655 11575 3661
rect 11517 3652 11529 3655
rect 9732 3624 11529 3652
rect 9732 3612 9738 3624
rect 11517 3621 11529 3624
rect 11563 3621 11575 3655
rect 11517 3615 11575 3621
rect 12253 3655 12311 3661
rect 12253 3621 12265 3655
rect 12299 3652 12311 3655
rect 14829 3655 14887 3661
rect 12299 3624 14320 3652
rect 12299 3621 12311 3624
rect 12253 3615 12311 3621
rect 6549 3587 6607 3593
rect 6549 3584 6561 3587
rect 6420 3556 6561 3584
rect 6420 3544 6426 3556
rect 6549 3553 6561 3556
rect 6595 3553 6607 3587
rect 6549 3547 6607 3553
rect 6825 3587 6883 3593
rect 6825 3553 6837 3587
rect 6871 3553 6883 3587
rect 6825 3547 6883 3553
rect 11054 3544 11060 3596
rect 11112 3584 11118 3596
rect 14182 3584 14188 3596
rect 11112 3556 11376 3584
rect 11112 3544 11118 3556
rect 5350 3516 5356 3528
rect 4356 3488 5356 3516
rect 4249 3479 4307 3485
rect 5350 3476 5356 3488
rect 5408 3476 5414 3528
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 9030 3516 9036 3528
rect 8435 3488 9036 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 9030 3476 9036 3488
rect 9088 3516 9094 3528
rect 9490 3516 9496 3528
rect 9088 3488 9496 3516
rect 9088 3476 9094 3488
rect 9490 3476 9496 3488
rect 9548 3476 9554 3528
rect 9677 3519 9735 3525
rect 9677 3485 9689 3519
rect 9723 3516 9735 3519
rect 9766 3516 9772 3528
rect 9723 3488 9772 3516
rect 9723 3485 9735 3488
rect 9677 3479 9735 3485
rect 9766 3476 9772 3488
rect 9824 3516 9830 3528
rect 10686 3516 10692 3528
rect 9824 3488 10692 3516
rect 9824 3476 9830 3488
rect 10686 3476 10692 3488
rect 10744 3476 10750 3528
rect 10873 3519 10931 3525
rect 10873 3485 10885 3519
rect 10919 3516 10931 3519
rect 11238 3516 11244 3528
rect 10919 3488 11244 3516
rect 10919 3485 10931 3488
rect 10873 3479 10931 3485
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 11348 3525 11376 3556
rect 13372 3556 14188 3584
rect 13372 3528 13400 3556
rect 14182 3544 14188 3556
rect 14240 3544 14246 3596
rect 14292 3593 14320 3624
rect 14829 3621 14841 3655
rect 14875 3621 14887 3655
rect 14829 3615 14887 3621
rect 18693 3655 18751 3661
rect 18693 3621 18705 3655
rect 18739 3652 18751 3655
rect 19150 3652 19156 3664
rect 18739 3624 19156 3652
rect 18739 3621 18751 3624
rect 18693 3615 18751 3621
rect 14277 3587 14335 3593
rect 14277 3553 14289 3587
rect 14323 3553 14335 3587
rect 14277 3547 14335 3553
rect 11333 3519 11391 3525
rect 11333 3485 11345 3519
rect 11379 3485 11391 3519
rect 12066 3516 12072 3528
rect 12027 3488 12072 3516
rect 11333 3479 11391 3485
rect 12066 3476 12072 3488
rect 12124 3476 12130 3528
rect 12897 3519 12955 3525
rect 12897 3485 12909 3519
rect 12943 3516 12955 3519
rect 13262 3516 13268 3528
rect 12943 3488 13268 3516
rect 12943 3485 12955 3488
rect 12897 3479 12955 3485
rect 13262 3476 13268 3488
rect 13320 3476 13326 3528
rect 13354 3476 13360 3528
rect 13412 3516 13418 3528
rect 13412 3488 13457 3516
rect 13412 3476 13418 3488
rect 13630 3476 13636 3528
rect 13688 3516 13694 3528
rect 14844 3516 14872 3615
rect 19150 3612 19156 3624
rect 19208 3612 19214 3664
rect 19242 3612 19248 3664
rect 19300 3652 19306 3664
rect 26234 3652 26240 3664
rect 19300 3624 26240 3652
rect 19300 3612 19306 3624
rect 26234 3612 26240 3624
rect 26292 3612 26298 3664
rect 46290 3612 46296 3664
rect 46348 3652 46354 3664
rect 46937 3655 46995 3661
rect 46937 3652 46949 3655
rect 46348 3624 46949 3652
rect 46348 3612 46354 3624
rect 46937 3621 46949 3624
rect 46983 3621 46995 3655
rect 46937 3615 46995 3621
rect 51442 3612 51448 3664
rect 51500 3652 51506 3664
rect 52825 3655 52883 3661
rect 52825 3652 52837 3655
rect 51500 3624 52837 3652
rect 51500 3612 51506 3624
rect 52825 3621 52837 3624
rect 52871 3621 52883 3655
rect 55186 3652 55214 3692
rect 55309 3655 55367 3661
rect 55309 3652 55321 3655
rect 55186 3624 55321 3652
rect 52825 3615 52883 3621
rect 55309 3621 55321 3624
rect 55355 3621 55367 3655
rect 55309 3615 55367 3621
rect 16022 3584 16028 3596
rect 15983 3556 16028 3584
rect 16022 3544 16028 3556
rect 16080 3544 16086 3596
rect 19613 3587 19671 3593
rect 19613 3553 19625 3587
rect 19659 3584 19671 3587
rect 21174 3584 21180 3596
rect 19659 3556 21180 3584
rect 19659 3553 19671 3556
rect 19613 3547 19671 3553
rect 21174 3544 21180 3556
rect 21232 3544 21238 3596
rect 21542 3544 21548 3596
rect 21600 3584 21606 3596
rect 21729 3587 21787 3593
rect 21729 3584 21741 3587
rect 21600 3556 21741 3584
rect 21600 3544 21606 3556
rect 21729 3553 21741 3556
rect 21775 3553 21787 3587
rect 21729 3547 21787 3553
rect 50798 3544 50804 3596
rect 50856 3584 50862 3596
rect 51537 3587 51595 3593
rect 51537 3584 51549 3587
rect 50856 3556 51549 3584
rect 50856 3544 50862 3556
rect 51537 3553 51549 3556
rect 51583 3553 51595 3587
rect 51537 3547 51595 3553
rect 51626 3544 51632 3596
rect 51684 3584 51690 3596
rect 53469 3587 53527 3593
rect 53469 3584 53481 3587
rect 51684 3556 53481 3584
rect 51684 3544 51690 3556
rect 53469 3553 53481 3556
rect 53515 3553 53527 3587
rect 53469 3547 53527 3553
rect 53834 3544 53840 3596
rect 53892 3584 53898 3596
rect 56597 3587 56655 3593
rect 56597 3584 56609 3587
rect 53892 3556 56609 3584
rect 53892 3544 53898 3556
rect 56597 3553 56609 3556
rect 56643 3553 56655 3587
rect 56597 3547 56655 3553
rect 13688 3488 14872 3516
rect 15565 3519 15623 3525
rect 13688 3476 13694 3488
rect 15565 3485 15577 3519
rect 15611 3485 15623 3519
rect 15565 3479 15623 3485
rect 2124 3451 2182 3457
rect 2124 3417 2136 3451
rect 2170 3448 2182 3451
rect 2590 3448 2596 3460
rect 2170 3420 2596 3448
rect 2170 3417 2182 3420
rect 2124 3411 2182 3417
rect 2590 3408 2596 3420
rect 2648 3408 2654 3460
rect 4516 3451 4574 3457
rect 4516 3417 4528 3451
rect 4562 3448 4574 3451
rect 4706 3448 4712 3460
rect 4562 3420 4712 3448
rect 4562 3417 4574 3420
rect 4516 3411 4574 3417
rect 4706 3408 4712 3420
rect 4764 3408 4770 3460
rect 5166 3408 5172 3460
rect 5224 3448 5230 3460
rect 6086 3448 6092 3460
rect 5224 3420 6092 3448
rect 5224 3408 5230 3420
rect 6086 3408 6092 3420
rect 6144 3408 6150 3460
rect 9122 3408 9128 3460
rect 9180 3448 9186 3460
rect 14369 3451 14427 3457
rect 14369 3448 14381 3451
rect 9180 3420 9536 3448
rect 9180 3408 9186 3420
rect 4062 3340 4068 3392
rect 4120 3380 4126 3392
rect 5629 3383 5687 3389
rect 5629 3380 5641 3383
rect 4120 3352 5641 3380
rect 4120 3340 4126 3352
rect 5629 3349 5641 3352
rect 5675 3349 5687 3383
rect 9508 3380 9536 3420
rect 13556 3420 14381 3448
rect 13556 3389 13584 3420
rect 14369 3417 14381 3420
rect 14415 3417 14427 3451
rect 14826 3448 14832 3460
rect 14787 3420 14832 3448
rect 14369 3411 14427 3417
rect 14826 3408 14832 3420
rect 14884 3408 14890 3460
rect 15580 3448 15608 3479
rect 16114 3476 16120 3528
rect 16172 3516 16178 3528
rect 16281 3519 16339 3525
rect 16281 3516 16293 3519
rect 16172 3488 16293 3516
rect 16172 3476 16178 3488
rect 16281 3485 16293 3488
rect 16327 3485 16339 3519
rect 16281 3479 16339 3485
rect 17402 3476 17408 3528
rect 17460 3516 17466 3528
rect 18322 3516 18328 3528
rect 17460 3488 18328 3516
rect 17460 3476 17466 3488
rect 18322 3476 18328 3488
rect 18380 3516 18386 3528
rect 18509 3519 18567 3525
rect 18509 3516 18521 3519
rect 18380 3488 18521 3516
rect 18380 3476 18386 3488
rect 18509 3485 18521 3488
rect 18555 3485 18567 3519
rect 20162 3516 20168 3528
rect 20123 3488 20168 3516
rect 18509 3479 18567 3485
rect 20162 3476 20168 3488
rect 20220 3476 20226 3528
rect 21634 3476 21640 3528
rect 21692 3516 21698 3528
rect 21818 3516 21824 3528
rect 21692 3488 21824 3516
rect 21692 3476 21698 3488
rect 21818 3476 21824 3488
rect 21876 3516 21882 3528
rect 21913 3519 21971 3525
rect 21913 3516 21925 3519
rect 21876 3488 21925 3516
rect 21876 3476 21882 3488
rect 21913 3485 21925 3488
rect 21959 3485 21971 3519
rect 21913 3479 21971 3485
rect 23201 3519 23259 3525
rect 23201 3485 23213 3519
rect 23247 3516 23259 3519
rect 23658 3516 23664 3528
rect 23247 3488 23664 3516
rect 23247 3485 23259 3488
rect 23201 3479 23259 3485
rect 23658 3476 23664 3488
rect 23716 3476 23722 3528
rect 23845 3519 23903 3525
rect 23845 3485 23857 3519
rect 23891 3516 23903 3519
rect 24210 3516 24216 3528
rect 23891 3488 24216 3516
rect 23891 3485 23903 3488
rect 23845 3479 23903 3485
rect 24210 3476 24216 3488
rect 24268 3476 24274 3528
rect 24762 3476 24768 3528
rect 24820 3516 24826 3528
rect 24857 3519 24915 3525
rect 24857 3516 24869 3519
rect 24820 3488 24869 3516
rect 24820 3476 24826 3488
rect 24857 3485 24869 3488
rect 24903 3485 24915 3519
rect 24857 3479 24915 3485
rect 25590 3476 25596 3528
rect 25648 3516 25654 3528
rect 25685 3519 25743 3525
rect 25685 3516 25697 3519
rect 25648 3488 25697 3516
rect 25648 3476 25654 3488
rect 25685 3485 25697 3488
rect 25731 3485 25743 3519
rect 25685 3479 25743 3485
rect 26694 3476 26700 3528
rect 26752 3516 26758 3528
rect 26789 3519 26847 3525
rect 26789 3516 26801 3519
rect 26752 3488 26801 3516
rect 26752 3476 26758 3488
rect 26789 3485 26801 3488
rect 26835 3485 26847 3519
rect 26789 3479 26847 3485
rect 27522 3476 27528 3528
rect 27580 3516 27586 3528
rect 27617 3519 27675 3525
rect 27617 3516 27629 3519
rect 27580 3488 27629 3516
rect 27580 3476 27586 3488
rect 27617 3485 27629 3488
rect 27663 3485 27675 3519
rect 27617 3479 27675 3485
rect 28626 3476 28632 3528
rect 28684 3516 28690 3528
rect 28721 3519 28779 3525
rect 28721 3516 28733 3519
rect 28684 3488 28733 3516
rect 28684 3476 28690 3488
rect 28721 3485 28733 3488
rect 28767 3485 28779 3519
rect 28721 3479 28779 3485
rect 30745 3519 30803 3525
rect 30745 3485 30757 3519
rect 30791 3516 30803 3519
rect 30791 3488 31248 3516
rect 30791 3485 30803 3488
rect 30745 3479 30803 3485
rect 31220 3460 31248 3488
rect 34698 3476 34704 3528
rect 34756 3516 34762 3528
rect 34793 3519 34851 3525
rect 34793 3516 34805 3519
rect 34756 3488 34805 3516
rect 34756 3476 34762 3488
rect 34793 3485 34805 3488
rect 34839 3485 34851 3519
rect 34793 3479 34851 3485
rect 35342 3476 35348 3528
rect 35400 3516 35406 3528
rect 35437 3519 35495 3525
rect 35437 3516 35449 3519
rect 35400 3488 35449 3516
rect 35400 3476 35406 3488
rect 35437 3485 35449 3488
rect 35483 3485 35495 3519
rect 35437 3479 35495 3485
rect 35802 3476 35808 3528
rect 35860 3516 35866 3528
rect 36081 3519 36139 3525
rect 36081 3516 36093 3519
rect 35860 3488 36093 3516
rect 35860 3476 35866 3488
rect 36081 3485 36093 3488
rect 36127 3485 36139 3519
rect 36081 3479 36139 3485
rect 36630 3476 36636 3528
rect 36688 3516 36694 3528
rect 36725 3519 36783 3525
rect 36725 3516 36737 3519
rect 36688 3488 36737 3516
rect 36688 3476 36694 3488
rect 36725 3485 36737 3488
rect 36771 3485 36783 3519
rect 36725 3479 36783 3485
rect 37458 3476 37464 3528
rect 37516 3516 37522 3528
rect 37553 3519 37611 3525
rect 37553 3516 37565 3519
rect 37516 3488 37565 3516
rect 37516 3476 37522 3488
rect 37553 3485 37565 3488
rect 37599 3485 37611 3519
rect 37553 3479 37611 3485
rect 38562 3476 38568 3528
rect 38620 3516 38626 3528
rect 38657 3519 38715 3525
rect 38657 3516 38669 3519
rect 38620 3488 38669 3516
rect 38620 3476 38626 3488
rect 38657 3485 38669 3488
rect 38703 3485 38715 3519
rect 38657 3479 38715 3485
rect 39942 3476 39948 3528
rect 40000 3516 40006 3528
rect 40037 3519 40095 3525
rect 40037 3516 40049 3519
rect 40000 3488 40049 3516
rect 40000 3476 40006 3488
rect 40037 3485 40049 3488
rect 40083 3485 40095 3519
rect 40037 3479 40095 3485
rect 40494 3476 40500 3528
rect 40552 3516 40558 3528
rect 40681 3519 40739 3525
rect 40681 3516 40693 3519
rect 40552 3488 40693 3516
rect 40552 3476 40558 3488
rect 40681 3485 40693 3488
rect 40727 3485 40739 3519
rect 40681 3479 40739 3485
rect 41046 3476 41052 3528
rect 41104 3516 41110 3528
rect 41325 3519 41383 3525
rect 41325 3516 41337 3519
rect 41104 3488 41337 3516
rect 41104 3476 41110 3488
rect 41325 3485 41337 3488
rect 41371 3485 41383 3519
rect 41325 3479 41383 3485
rect 42426 3476 42432 3528
rect 42484 3516 42490 3528
rect 42521 3519 42579 3525
rect 42521 3516 42533 3519
rect 42484 3488 42533 3516
rect 42484 3476 42490 3488
rect 42521 3485 42533 3488
rect 42567 3485 42579 3519
rect 42521 3479 42579 3485
rect 42702 3476 42708 3528
rect 42760 3516 42766 3528
rect 43165 3519 43223 3525
rect 43165 3516 43177 3519
rect 42760 3488 43177 3516
rect 42760 3476 42766 3488
rect 43165 3485 43177 3488
rect 43211 3485 43223 3519
rect 43165 3479 43223 3485
rect 44358 3476 44364 3528
rect 44416 3516 44422 3528
rect 45005 3519 45063 3525
rect 45005 3516 45017 3519
rect 44416 3488 45017 3516
rect 44416 3476 44422 3488
rect 45005 3485 45017 3488
rect 45051 3485 45063 3519
rect 45005 3479 45063 3485
rect 45186 3476 45192 3528
rect 45244 3516 45250 3528
rect 45649 3519 45707 3525
rect 45649 3516 45661 3519
rect 45244 3488 45661 3516
rect 45244 3476 45250 3488
rect 45649 3485 45661 3488
rect 45695 3485 45707 3519
rect 45649 3479 45707 3485
rect 46014 3476 46020 3528
rect 46072 3516 46078 3528
rect 46293 3519 46351 3525
rect 46293 3516 46305 3519
rect 46072 3488 46305 3516
rect 46072 3476 46078 3488
rect 46293 3485 46305 3488
rect 46339 3485 46351 3519
rect 46293 3479 46351 3485
rect 47670 3476 47676 3528
rect 47728 3516 47734 3528
rect 47765 3519 47823 3525
rect 47765 3516 47777 3519
rect 47728 3488 47777 3516
rect 47728 3476 47734 3488
rect 47765 3485 47777 3488
rect 47811 3485 47823 3519
rect 47765 3479 47823 3485
rect 48222 3476 48228 3528
rect 48280 3516 48286 3528
rect 48409 3519 48467 3525
rect 48409 3516 48421 3519
rect 48280 3488 48421 3516
rect 48280 3476 48286 3488
rect 48409 3485 48421 3488
rect 48455 3485 48467 3519
rect 48409 3479 48467 3485
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50249 3519 50307 3525
rect 50249 3516 50261 3519
rect 50212 3488 50261 3516
rect 50212 3476 50218 3488
rect 50249 3485 50261 3488
rect 50295 3485 50307 3519
rect 50249 3479 50307 3485
rect 50614 3476 50620 3528
rect 50672 3516 50678 3528
rect 50893 3519 50951 3525
rect 50893 3516 50905 3519
rect 50672 3488 50905 3516
rect 50672 3476 50678 3488
rect 50893 3485 50905 3488
rect 50939 3485 50951 3519
rect 50893 3479 50951 3485
rect 51166 3476 51172 3528
rect 51224 3516 51230 3528
rect 52181 3519 52239 3525
rect 52181 3516 52193 3519
rect 51224 3488 52193 3516
rect 51224 3476 51230 3488
rect 52181 3485 52193 3488
rect 52227 3485 52239 3519
rect 52181 3479 52239 3485
rect 52270 3476 52276 3528
rect 52328 3516 52334 3528
rect 54113 3519 54171 3525
rect 54113 3516 54125 3519
rect 52328 3488 54125 3516
rect 52328 3476 52334 3488
rect 54113 3485 54125 3488
rect 54159 3485 54171 3519
rect 55953 3519 56011 3525
rect 55953 3516 55965 3519
rect 54113 3479 54171 3485
rect 55186 3488 55965 3516
rect 17957 3451 18015 3457
rect 15580 3420 17908 3448
rect 10689 3383 10747 3389
rect 10689 3380 10701 3383
rect 9508 3352 10701 3380
rect 5629 3343 5687 3349
rect 10689 3349 10701 3352
rect 10735 3349 10747 3383
rect 10689 3343 10747 3349
rect 13541 3383 13599 3389
rect 13541 3349 13553 3383
rect 13587 3349 13599 3383
rect 14090 3380 14096 3392
rect 14051 3352 14096 3380
rect 13541 3343 13599 3349
rect 14090 3340 14096 3352
rect 14148 3340 14154 3392
rect 15746 3340 15752 3392
rect 15804 3380 15810 3392
rect 16022 3380 16028 3392
rect 15804 3352 16028 3380
rect 15804 3340 15810 3352
rect 16022 3340 16028 3352
rect 16080 3340 16086 3392
rect 17880 3380 17908 3420
rect 17957 3417 17969 3451
rect 18003 3448 18015 3451
rect 20806 3448 20812 3460
rect 18003 3420 20812 3448
rect 18003 3417 18015 3420
rect 17957 3411 18015 3417
rect 20806 3408 20812 3420
rect 20864 3448 20870 3460
rect 21085 3451 21143 3457
rect 21085 3448 21097 3451
rect 20864 3420 21097 3448
rect 20864 3408 20870 3420
rect 21085 3417 21097 3420
rect 21131 3417 21143 3451
rect 21085 3411 21143 3417
rect 30834 3408 30840 3460
rect 30892 3448 30898 3460
rect 30990 3451 31048 3457
rect 30990 3448 31002 3451
rect 30892 3420 31002 3448
rect 30892 3408 30898 3420
rect 30990 3417 31002 3420
rect 31036 3417 31048 3451
rect 30990 3411 31048 3417
rect 31202 3408 31208 3460
rect 31260 3408 31266 3460
rect 53282 3408 53288 3460
rect 53340 3448 53346 3460
rect 55186 3448 55214 3488
rect 55953 3485 55965 3488
rect 55999 3485 56011 3519
rect 57514 3516 57520 3528
rect 57475 3488 57520 3516
rect 55953 3479 56011 3485
rect 57514 3476 57520 3488
rect 57572 3476 57578 3528
rect 58158 3516 58164 3528
rect 58119 3488 58164 3516
rect 58158 3476 58164 3488
rect 58216 3476 58222 3528
rect 53340 3420 55214 3448
rect 53340 3408 53346 3420
rect 18874 3380 18880 3392
rect 17880 3352 18880 3380
rect 18874 3340 18880 3352
rect 18932 3340 18938 3392
rect 19702 3340 19708 3392
rect 19760 3380 19766 3392
rect 20162 3380 20168 3392
rect 19760 3352 20168 3380
rect 19760 3340 19766 3352
rect 20162 3340 20168 3352
rect 20220 3340 20226 3392
rect 22557 3383 22615 3389
rect 22557 3349 22569 3383
rect 22603 3380 22615 3383
rect 22830 3380 22836 3392
rect 22603 3352 22836 3380
rect 22603 3349 22615 3352
rect 22557 3343 22615 3349
rect 22830 3340 22836 3352
rect 22888 3340 22894 3392
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 1857 3179 1915 3185
rect 1857 3145 1869 3179
rect 1903 3176 1915 3179
rect 3418 3176 3424 3188
rect 1903 3148 3424 3176
rect 1903 3145 1915 3148
rect 1857 3139 1915 3145
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 3786 3176 3792 3188
rect 3747 3148 3792 3176
rect 3786 3136 3792 3148
rect 3844 3136 3850 3188
rect 3878 3136 3884 3188
rect 3936 3176 3942 3188
rect 5350 3176 5356 3188
rect 3936 3148 5356 3176
rect 3936 3136 3942 3148
rect 5350 3136 5356 3148
rect 5408 3136 5414 3188
rect 5655 3179 5713 3185
rect 5655 3145 5667 3179
rect 5701 3176 5713 3179
rect 8202 3176 8208 3188
rect 5701 3148 8208 3176
rect 5701 3145 5713 3148
rect 5655 3139 5713 3145
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 9766 3176 9772 3188
rect 8312 3148 9772 3176
rect 1946 3068 1952 3120
rect 2004 3108 2010 3120
rect 2654 3111 2712 3117
rect 2654 3108 2666 3111
rect 2004 3080 2666 3108
rect 2004 3068 2010 3080
rect 2654 3077 2666 3080
rect 2700 3077 2712 3111
rect 2654 3071 2712 3077
rect 4614 3068 4620 3120
rect 4672 3108 4678 3120
rect 5445 3111 5503 3117
rect 5445 3108 5457 3111
rect 4672 3080 5457 3108
rect 4672 3068 4678 3080
rect 5445 3077 5457 3080
rect 5491 3077 5503 3111
rect 5445 3071 5503 3077
rect 1486 3000 1492 3052
rect 1544 3040 1550 3052
rect 1765 3043 1823 3049
rect 1765 3040 1777 3043
rect 1544 3012 1777 3040
rect 1544 3000 1550 3012
rect 1765 3009 1777 3012
rect 1811 3009 1823 3043
rect 2406 3040 2412 3052
rect 2367 3012 2412 3040
rect 1765 3003 1823 3009
rect 1780 2972 1808 3003
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 4985 3043 5043 3049
rect 2516 3012 4016 3040
rect 2516 2972 2544 3012
rect 1780 2944 2544 2972
rect 3988 2972 4016 3012
rect 4985 3009 4997 3043
rect 5031 3040 5043 3043
rect 5074 3040 5080 3052
rect 5031 3012 5080 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 5074 3000 5080 3012
rect 5132 3040 5138 3052
rect 6733 3043 6791 3049
rect 5132 3012 6684 3040
rect 5132 3000 5138 3012
rect 5258 2972 5264 2984
rect 3988 2944 5264 2972
rect 5258 2932 5264 2944
rect 5316 2932 5322 2984
rect 6656 2972 6684 3012
rect 6733 3009 6745 3043
rect 6779 3040 6791 3043
rect 6822 3040 6828 3052
rect 6779 3012 6828 3040
rect 6779 3009 6791 3012
rect 6733 3003 6791 3009
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3040 7067 3043
rect 7282 3040 7288 3052
rect 7055 3012 7288 3040
rect 7055 3009 7067 3012
rect 7009 3003 7067 3009
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 7926 3000 7932 3052
rect 7984 3040 7990 3052
rect 8021 3043 8079 3049
rect 8021 3040 8033 3043
rect 7984 3012 8033 3040
rect 7984 3000 7990 3012
rect 8021 3009 8033 3012
rect 8067 3009 8079 3043
rect 8021 3003 8079 3009
rect 8202 3000 8208 3052
rect 8260 3040 8266 3052
rect 8312 3040 8340 3148
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 13541 3179 13599 3185
rect 13541 3145 13553 3179
rect 13587 3176 13599 3179
rect 13630 3176 13636 3188
rect 13587 3148 13636 3176
rect 13587 3145 13599 3148
rect 13541 3139 13599 3145
rect 13630 3136 13636 3148
rect 13688 3136 13694 3188
rect 14550 3176 14556 3188
rect 14511 3148 14556 3176
rect 14550 3136 14556 3148
rect 14608 3136 14614 3188
rect 15194 3176 15200 3188
rect 15155 3148 15200 3176
rect 15194 3136 15200 3148
rect 15252 3136 15258 3188
rect 15933 3179 15991 3185
rect 15933 3145 15945 3179
rect 15979 3176 15991 3179
rect 16114 3176 16120 3188
rect 15979 3148 16120 3176
rect 15979 3145 15991 3148
rect 15933 3139 15991 3145
rect 16114 3136 16120 3148
rect 16172 3136 16178 3188
rect 17402 3176 17408 3188
rect 17363 3148 17408 3176
rect 17402 3136 17408 3148
rect 17460 3136 17466 3188
rect 17770 3176 17776 3188
rect 17604 3148 17776 3176
rect 8570 3068 8576 3120
rect 8628 3068 8634 3120
rect 8846 3068 8852 3120
rect 8904 3108 8910 3120
rect 10410 3108 10416 3120
rect 8904 3080 9536 3108
rect 10371 3080 10416 3108
rect 8904 3068 8910 3080
rect 8260 3012 8340 3040
rect 8260 3000 8266 3012
rect 7650 2972 7656 2984
rect 5368 2944 5948 2972
rect 6656 2944 7656 2972
rect 5368 2904 5396 2944
rect 5810 2904 5816 2916
rect 4724 2876 5396 2904
rect 5771 2876 5816 2904
rect 2682 2796 2688 2848
rect 2740 2836 2746 2848
rect 4724 2836 4752 2876
rect 5810 2864 5816 2876
rect 5868 2864 5874 2916
rect 5920 2904 5948 2944
rect 7650 2932 7656 2944
rect 7708 2932 7714 2984
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 8478 2972 8484 2984
rect 7800 2944 8484 2972
rect 7800 2932 7806 2944
rect 7834 2904 7840 2916
rect 5920 2876 7840 2904
rect 7834 2864 7840 2876
rect 7892 2864 7898 2916
rect 7944 2904 7972 2944
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 8588 2981 8616 3068
rect 8662 3000 8668 3052
rect 8720 3000 8726 3052
rect 8938 3040 8944 3052
rect 8899 3012 8944 3040
rect 8938 3000 8944 3012
rect 8996 3000 9002 3052
rect 9508 3049 9536 3080
rect 10410 3068 10416 3080
rect 10468 3068 10474 3120
rect 17034 3108 17040 3120
rect 12912 3080 17040 3108
rect 9493 3043 9551 3049
rect 9493 3009 9505 3043
rect 9539 3009 9551 3043
rect 9858 3040 9864 3052
rect 9819 3012 9864 3040
rect 9493 3003 9551 3009
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 10781 3043 10839 3049
rect 10781 3009 10793 3043
rect 10827 3040 10839 3043
rect 10962 3040 10968 3052
rect 10827 3012 10968 3040
rect 10827 3009 10839 3012
rect 10781 3003 10839 3009
rect 10962 3000 10968 3012
rect 11020 3000 11026 3052
rect 11514 3040 11520 3052
rect 11475 3012 11520 3040
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 12912 3049 12940 3080
rect 17034 3068 17040 3080
rect 17092 3068 17098 3120
rect 12897 3043 12955 3049
rect 12897 3009 12909 3043
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 13078 3000 13084 3052
rect 13136 3040 13142 3052
rect 13357 3043 13415 3049
rect 13357 3040 13369 3043
rect 13136 3012 13369 3040
rect 13136 3000 13142 3012
rect 13357 3009 13369 3012
rect 13403 3009 13415 3043
rect 13357 3003 13415 3009
rect 14369 3043 14427 3049
rect 14369 3009 14381 3043
rect 14415 3040 14427 3043
rect 14458 3040 14464 3052
rect 14415 3012 14464 3040
rect 14415 3009 14427 3012
rect 14369 3003 14427 3009
rect 8573 2975 8631 2981
rect 8573 2941 8585 2975
rect 8619 2941 8631 2975
rect 8680 2972 8708 3000
rect 13372 2972 13400 3003
rect 14458 3000 14464 3012
rect 14516 3040 14522 3052
rect 15381 3043 15439 3049
rect 14516 3012 15332 3040
rect 14516 3000 14522 3012
rect 15010 2972 15016 2984
rect 8680 2944 11744 2972
rect 13372 2944 15016 2972
rect 8573 2935 8631 2941
rect 7944 2876 8064 2904
rect 2740 2808 4752 2836
rect 4801 2839 4859 2845
rect 2740 2796 2746 2808
rect 4801 2805 4813 2839
rect 4847 2836 4859 2839
rect 4890 2836 4896 2848
rect 4847 2808 4896 2836
rect 4847 2805 4859 2808
rect 4801 2799 4859 2805
rect 4890 2796 4896 2808
rect 4948 2796 4954 2848
rect 5626 2836 5632 2848
rect 5587 2808 5632 2836
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 7466 2796 7472 2848
rect 7524 2836 7530 2848
rect 7926 2836 7932 2848
rect 7524 2808 7932 2836
rect 7524 2796 7530 2808
rect 7926 2796 7932 2808
rect 7984 2796 7990 2848
rect 8036 2836 8064 2876
rect 9030 2864 9036 2916
rect 9088 2904 9094 2916
rect 9088 2876 9352 2904
rect 9088 2864 9094 2876
rect 8389 2839 8447 2845
rect 8389 2836 8401 2839
rect 8036 2808 8401 2836
rect 8389 2805 8401 2808
rect 8435 2805 8447 2839
rect 8389 2799 8447 2805
rect 8481 2839 8539 2845
rect 8481 2805 8493 2839
rect 8527 2836 8539 2839
rect 9214 2836 9220 2848
rect 8527 2808 9220 2836
rect 8527 2805 8539 2808
rect 8481 2799 8539 2805
rect 9214 2796 9220 2808
rect 9272 2796 9278 2848
rect 9324 2836 9352 2876
rect 9398 2864 9404 2916
rect 9456 2904 9462 2916
rect 11054 2904 11060 2916
rect 9456 2876 11060 2904
rect 9456 2864 9462 2876
rect 11054 2864 11060 2876
rect 11112 2864 11118 2916
rect 11716 2913 11744 2944
rect 15010 2932 15016 2944
rect 15068 2932 15074 2984
rect 15304 2972 15332 3012
rect 15381 3009 15393 3043
rect 15427 3040 15439 3043
rect 15654 3040 15660 3052
rect 15427 3012 15660 3040
rect 15427 3009 15439 3012
rect 15381 3003 15439 3009
rect 15654 3000 15660 3012
rect 15712 3000 15718 3052
rect 16117 3043 16175 3049
rect 16117 3009 16129 3043
rect 16163 3040 16175 3043
rect 16390 3040 16396 3052
rect 16163 3012 16396 3040
rect 16163 3009 16175 3012
rect 16117 3003 16175 3009
rect 16390 3000 16396 3012
rect 16448 3040 16454 3052
rect 16942 3040 16948 3052
rect 16448 3012 16948 3040
rect 16448 3000 16454 3012
rect 16942 3000 16948 3012
rect 17000 3000 17006 3052
rect 17604 3049 17632 3148
rect 17770 3136 17776 3148
rect 17828 3176 17834 3188
rect 21082 3176 21088 3188
rect 17828 3148 21088 3176
rect 17828 3136 17834 3148
rect 21082 3136 21088 3148
rect 21140 3136 21146 3188
rect 23014 3176 23020 3188
rect 22975 3148 23020 3176
rect 23014 3136 23020 3148
rect 23072 3136 23078 3188
rect 18046 3108 18052 3120
rect 18007 3080 18052 3108
rect 18046 3068 18052 3080
rect 18104 3068 18110 3120
rect 18782 3108 18788 3120
rect 18743 3080 18788 3108
rect 18782 3068 18788 3080
rect 18840 3068 18846 3120
rect 18969 3111 19027 3117
rect 18969 3077 18981 3111
rect 19015 3108 19027 3111
rect 19058 3108 19064 3120
rect 19015 3080 19064 3108
rect 19015 3077 19027 3080
rect 18969 3071 19027 3077
rect 19058 3068 19064 3080
rect 19116 3068 19122 3120
rect 20441 3111 20499 3117
rect 20441 3077 20453 3111
rect 20487 3108 20499 3111
rect 20622 3108 20628 3120
rect 20487 3080 20628 3108
rect 20487 3077 20499 3080
rect 20441 3071 20499 3077
rect 20622 3068 20628 3080
rect 20680 3108 20686 3120
rect 20990 3108 20996 3120
rect 20680 3080 20852 3108
rect 20951 3080 20996 3108
rect 20680 3068 20686 3080
rect 17589 3043 17647 3049
rect 17589 3009 17601 3043
rect 17635 3009 17647 3043
rect 17589 3003 17647 3009
rect 18233 3043 18291 3049
rect 18233 3009 18245 3043
rect 18279 3040 18291 3043
rect 18506 3040 18512 3052
rect 18279 3012 18512 3040
rect 18279 3009 18291 3012
rect 18233 3003 18291 3009
rect 18506 3000 18512 3012
rect 18564 3040 18570 3052
rect 18690 3040 18696 3052
rect 18564 3012 18696 3040
rect 18564 3000 18570 3012
rect 18690 3000 18696 3012
rect 18748 3000 18754 3052
rect 19797 3043 19855 3049
rect 19797 3009 19809 3043
rect 19843 3040 19855 3043
rect 19978 3040 19984 3052
rect 19843 3012 19984 3040
rect 19843 3009 19855 3012
rect 19797 3003 19855 3009
rect 19978 3000 19984 3012
rect 20036 3000 20042 3052
rect 15562 2972 15568 2984
rect 15304 2944 15568 2972
rect 15562 2932 15568 2944
rect 15620 2932 15626 2984
rect 11701 2907 11759 2913
rect 11701 2873 11713 2907
rect 11747 2873 11759 2907
rect 11701 2867 11759 2873
rect 12066 2864 12072 2916
rect 12124 2904 12130 2916
rect 14458 2904 14464 2916
rect 12124 2876 14464 2904
rect 12124 2864 12130 2876
rect 14458 2864 14464 2876
rect 14516 2864 14522 2916
rect 15672 2904 15700 3000
rect 19058 2932 19064 2984
rect 19116 2972 19122 2984
rect 19242 2972 19248 2984
rect 19116 2944 19248 2972
rect 19116 2932 19122 2944
rect 19242 2932 19248 2944
rect 19300 2932 19306 2984
rect 19610 2932 19616 2984
rect 19668 2972 19674 2984
rect 20257 2975 20315 2981
rect 20257 2972 20269 2975
rect 19668 2944 20269 2972
rect 19668 2932 19674 2944
rect 20257 2941 20269 2944
rect 20303 2941 20315 2975
rect 20257 2935 20315 2941
rect 20346 2932 20352 2984
rect 20404 2972 20410 2984
rect 20622 2972 20628 2984
rect 20404 2944 20628 2972
rect 20404 2932 20410 2944
rect 20622 2932 20628 2944
rect 20680 2932 20686 2984
rect 16390 2904 16396 2916
rect 15672 2876 16396 2904
rect 16390 2864 16396 2876
rect 16448 2864 16454 2916
rect 19426 2864 19432 2916
rect 19484 2904 19490 2916
rect 19886 2904 19892 2916
rect 19484 2876 19892 2904
rect 19484 2864 19490 2876
rect 19886 2864 19892 2876
rect 19944 2864 19950 2916
rect 10410 2836 10416 2848
rect 9324 2808 10416 2836
rect 10410 2796 10416 2808
rect 10468 2796 10474 2848
rect 15102 2796 15108 2848
rect 15160 2836 15166 2848
rect 16666 2836 16672 2848
rect 15160 2808 16672 2836
rect 15160 2796 15166 2808
rect 16666 2796 16672 2808
rect 16724 2796 16730 2848
rect 16853 2839 16911 2845
rect 16853 2805 16865 2839
rect 16899 2836 16911 2839
rect 18414 2836 18420 2848
rect 16899 2808 18420 2836
rect 16899 2805 16911 2808
rect 16853 2799 16911 2805
rect 18414 2796 18420 2808
rect 18472 2796 18478 2848
rect 19613 2839 19671 2845
rect 19613 2805 19625 2839
rect 19659 2836 19671 2839
rect 19794 2836 19800 2848
rect 19659 2808 19800 2836
rect 19659 2805 19671 2808
rect 19613 2799 19671 2805
rect 19794 2796 19800 2808
rect 19852 2796 19858 2848
rect 20530 2796 20536 2848
rect 20588 2836 20594 2848
rect 20824 2836 20852 3080
rect 20990 3068 20996 3080
rect 21048 3068 21054 3120
rect 21177 3111 21235 3117
rect 21177 3077 21189 3111
rect 21223 3108 21235 3111
rect 21358 3108 21364 3120
rect 21223 3080 21364 3108
rect 21223 3077 21235 3080
rect 21177 3071 21235 3077
rect 21358 3068 21364 3080
rect 21416 3068 21422 3120
rect 22186 3108 22192 3120
rect 22147 3080 22192 3108
rect 22186 3068 22192 3080
rect 22244 3068 22250 3120
rect 22370 3108 22376 3120
rect 22331 3080 22376 3108
rect 22370 3068 22376 3080
rect 22428 3068 22434 3120
rect 51902 3068 51908 3120
rect 51960 3108 51966 3120
rect 51960 3080 54708 3108
rect 51960 3068 51966 3080
rect 22830 3040 22836 3052
rect 22791 3012 22836 3040
rect 22830 3000 22836 3012
rect 22888 3000 22894 3052
rect 51718 3000 51724 3052
rect 51776 3040 51782 3052
rect 54680 3049 54708 3080
rect 54021 3043 54079 3049
rect 54021 3040 54033 3043
rect 51776 3012 54033 3040
rect 51776 3000 51782 3012
rect 54021 3009 54033 3012
rect 54067 3009 54079 3043
rect 54021 3003 54079 3009
rect 54665 3043 54723 3049
rect 54665 3009 54677 3043
rect 54711 3009 54723 3043
rect 54665 3003 54723 3009
rect 54754 3000 54760 3052
rect 54812 3040 54818 3052
rect 55309 3043 55367 3049
rect 55309 3040 55321 3043
rect 54812 3012 55321 3040
rect 54812 3000 54818 3012
rect 55309 3009 55321 3012
rect 55355 3009 55367 3043
rect 55309 3003 55367 3009
rect 23845 2975 23903 2981
rect 23845 2941 23857 2975
rect 23891 2972 23903 2975
rect 24486 2972 24492 2984
rect 23891 2944 24492 2972
rect 23891 2941 23903 2944
rect 23845 2935 23903 2941
rect 24486 2932 24492 2944
rect 24544 2932 24550 2984
rect 32766 2932 32772 2984
rect 32824 2972 32830 2984
rect 33413 2975 33471 2981
rect 33413 2972 33425 2975
rect 32824 2944 33425 2972
rect 32824 2932 32830 2944
rect 33413 2941 33425 2944
rect 33459 2941 33471 2975
rect 33413 2935 33471 2941
rect 38286 2932 38292 2984
rect 38344 2972 38350 2984
rect 39209 2975 39267 2981
rect 39209 2972 39221 2975
rect 38344 2944 39221 2972
rect 38344 2932 38350 2944
rect 39209 2941 39221 2944
rect 39255 2941 39267 2975
rect 39209 2935 39267 2941
rect 42150 2932 42156 2984
rect 42208 2972 42214 2984
rect 43073 2975 43131 2981
rect 43073 2972 43085 2975
rect 42208 2944 43085 2972
rect 42208 2932 42214 2944
rect 43073 2941 43085 2944
rect 43119 2941 43131 2975
rect 43073 2935 43131 2941
rect 53098 2932 53104 2984
rect 53156 2972 53162 2984
rect 55953 2975 56011 2981
rect 55953 2972 55965 2975
rect 53156 2944 55965 2972
rect 53156 2932 53162 2944
rect 55953 2941 55965 2944
rect 55999 2941 56011 2975
rect 56594 2972 56600 2984
rect 56555 2944 56600 2972
rect 55953 2935 56011 2941
rect 56594 2932 56600 2944
rect 56652 2932 56658 2984
rect 33870 2864 33876 2916
rect 33928 2904 33934 2916
rect 34701 2907 34759 2913
rect 34701 2904 34713 2907
rect 33928 2876 34713 2904
rect 33928 2864 33934 2876
rect 34701 2873 34713 2876
rect 34747 2873 34759 2907
rect 34701 2867 34759 2873
rect 37182 2864 37188 2916
rect 37240 2904 37246 2916
rect 37921 2907 37979 2913
rect 37921 2904 37933 2907
rect 37240 2876 37933 2904
rect 37240 2864 37246 2876
rect 37921 2873 37933 2876
rect 37967 2873 37979 2907
rect 37921 2867 37979 2873
rect 39114 2864 39120 2916
rect 39172 2904 39178 2916
rect 39853 2907 39911 2913
rect 39853 2904 39865 2907
rect 39172 2876 39865 2904
rect 39172 2864 39178 2876
rect 39853 2873 39865 2876
rect 39899 2873 39911 2907
rect 39853 2867 39911 2873
rect 40218 2864 40224 2916
rect 40276 2904 40282 2916
rect 41141 2907 41199 2913
rect 41141 2904 41153 2907
rect 40276 2876 41153 2904
rect 40276 2864 40282 2876
rect 41141 2873 41153 2876
rect 41187 2873 41199 2907
rect 41141 2867 41199 2873
rect 42978 2864 42984 2916
rect 43036 2904 43042 2916
rect 43717 2907 43775 2913
rect 43717 2904 43729 2907
rect 43036 2876 43729 2904
rect 43036 2864 43042 2876
rect 43717 2873 43729 2876
rect 43763 2873 43775 2907
rect 43717 2867 43775 2873
rect 44082 2864 44088 2916
rect 44140 2904 44146 2916
rect 45005 2907 45063 2913
rect 45005 2904 45017 2907
rect 44140 2876 45017 2904
rect 44140 2864 44146 2876
rect 45005 2873 45017 2876
rect 45051 2873 45063 2907
rect 45649 2907 45707 2913
rect 45649 2904 45661 2907
rect 45005 2867 45063 2873
rect 45112 2876 45661 2904
rect 20588 2808 20852 2836
rect 20588 2796 20594 2808
rect 22462 2796 22468 2848
rect 22520 2836 22526 2848
rect 22830 2836 22836 2848
rect 22520 2808 22836 2836
rect 22520 2796 22526 2808
rect 22830 2796 22836 2808
rect 22888 2796 22894 2848
rect 24489 2839 24547 2845
rect 24489 2805 24501 2839
rect 24535 2836 24547 2839
rect 25038 2836 25044 2848
rect 24535 2808 25044 2836
rect 24535 2805 24547 2808
rect 24489 2799 24547 2805
rect 25038 2796 25044 2808
rect 25096 2796 25102 2848
rect 25133 2839 25191 2845
rect 25133 2805 25145 2839
rect 25179 2836 25191 2839
rect 25314 2836 25320 2848
rect 25179 2808 25320 2836
rect 25179 2805 25191 2808
rect 25133 2799 25191 2805
rect 25314 2796 25320 2808
rect 25372 2796 25378 2848
rect 25777 2839 25835 2845
rect 25777 2805 25789 2839
rect 25823 2836 25835 2839
rect 26142 2836 26148 2848
rect 25823 2808 26148 2836
rect 25823 2805 25835 2808
rect 25777 2799 25835 2805
rect 26142 2796 26148 2808
rect 26200 2796 26206 2848
rect 26421 2839 26479 2845
rect 26421 2805 26433 2839
rect 26467 2836 26479 2839
rect 26970 2836 26976 2848
rect 26467 2808 26976 2836
rect 26467 2805 26479 2808
rect 26421 2799 26479 2805
rect 26970 2796 26976 2808
rect 27028 2796 27034 2848
rect 27617 2839 27675 2845
rect 27617 2805 27629 2839
rect 27663 2836 27675 2839
rect 27798 2836 27804 2848
rect 27663 2808 27804 2836
rect 27663 2805 27675 2808
rect 27617 2799 27675 2805
rect 27798 2796 27804 2808
rect 27856 2796 27862 2848
rect 28074 2836 28080 2848
rect 28035 2808 28080 2836
rect 28074 2796 28080 2808
rect 28132 2796 28138 2848
rect 28905 2839 28963 2845
rect 28905 2805 28917 2839
rect 28951 2836 28963 2839
rect 29178 2836 29184 2848
rect 28951 2808 29184 2836
rect 28951 2805 28963 2808
rect 28905 2799 28963 2805
rect 29178 2796 29184 2808
rect 29236 2796 29242 2848
rect 29549 2839 29607 2845
rect 29549 2805 29561 2839
rect 29595 2836 29607 2839
rect 29730 2836 29736 2848
rect 29595 2808 29736 2836
rect 29595 2805 29607 2808
rect 29549 2799 29607 2805
rect 29730 2796 29736 2808
rect 29788 2796 29794 2848
rect 30006 2836 30012 2848
rect 29967 2808 30012 2836
rect 30006 2796 30012 2808
rect 30064 2796 30070 2848
rect 30558 2796 30564 2848
rect 30616 2836 30622 2848
rect 30653 2839 30711 2845
rect 30653 2836 30665 2839
rect 30616 2808 30665 2836
rect 30616 2796 30622 2808
rect 30653 2805 30665 2808
rect 30699 2805 30711 2839
rect 30653 2799 30711 2805
rect 31662 2796 31668 2848
rect 31720 2836 31726 2848
rect 32125 2839 32183 2845
rect 32125 2836 32137 2839
rect 31720 2808 32137 2836
rect 31720 2796 31726 2808
rect 32125 2805 32137 2808
rect 32171 2805 32183 2839
rect 32125 2799 32183 2805
rect 32214 2796 32220 2848
rect 32272 2836 32278 2848
rect 32769 2839 32827 2845
rect 32769 2836 32781 2839
rect 32272 2808 32781 2836
rect 32272 2796 32278 2808
rect 32769 2805 32781 2808
rect 32815 2805 32827 2839
rect 32769 2799 32827 2805
rect 33318 2796 33324 2848
rect 33376 2836 33382 2848
rect 34057 2839 34115 2845
rect 34057 2836 34069 2839
rect 33376 2808 34069 2836
rect 33376 2796 33382 2808
rect 34057 2805 34069 2808
rect 34103 2805 34115 2839
rect 34057 2799 34115 2805
rect 34422 2796 34428 2848
rect 34480 2836 34486 2848
rect 35345 2839 35403 2845
rect 35345 2836 35357 2839
rect 34480 2808 35357 2836
rect 34480 2796 34486 2808
rect 35345 2805 35357 2808
rect 35391 2805 35403 2839
rect 35345 2799 35403 2805
rect 35434 2796 35440 2848
rect 35492 2836 35498 2848
rect 35989 2839 36047 2845
rect 35989 2836 36001 2839
rect 35492 2808 36001 2836
rect 35492 2796 35498 2808
rect 35989 2805 36001 2808
rect 36035 2805 36047 2839
rect 35989 2799 36047 2805
rect 36354 2796 36360 2848
rect 36412 2836 36418 2848
rect 37277 2839 37335 2845
rect 37277 2836 37289 2839
rect 36412 2808 37289 2836
rect 36412 2796 36418 2808
rect 37277 2805 37289 2808
rect 37323 2805 37335 2839
rect 37277 2799 37335 2805
rect 37734 2796 37740 2848
rect 37792 2836 37798 2848
rect 38565 2839 38623 2845
rect 38565 2836 38577 2839
rect 37792 2808 38577 2836
rect 37792 2796 37798 2808
rect 38565 2805 38577 2808
rect 38611 2805 38623 2839
rect 38565 2799 38623 2805
rect 39666 2796 39672 2848
rect 39724 2836 39730 2848
rect 40497 2839 40555 2845
rect 40497 2836 40509 2839
rect 39724 2808 40509 2836
rect 39724 2796 39730 2808
rect 40497 2805 40509 2808
rect 40543 2805 40555 2839
rect 40497 2799 40555 2805
rect 41598 2796 41604 2848
rect 41656 2836 41662 2848
rect 42429 2839 42487 2845
rect 42429 2836 42441 2839
rect 41656 2808 42441 2836
rect 41656 2796 41662 2808
rect 42429 2805 42441 2808
rect 42475 2805 42487 2839
rect 42429 2799 42487 2805
rect 43530 2796 43536 2848
rect 43588 2836 43594 2848
rect 44361 2839 44419 2845
rect 44361 2836 44373 2839
rect 43588 2808 44373 2836
rect 43588 2796 43594 2808
rect 44361 2805 44373 2808
rect 44407 2805 44419 2839
rect 44361 2799 44419 2805
rect 44910 2796 44916 2848
rect 44968 2836 44974 2848
rect 45112 2836 45140 2876
rect 45649 2873 45661 2876
rect 45695 2873 45707 2907
rect 45649 2867 45707 2873
rect 47394 2864 47400 2916
rect 47452 2904 47458 2916
rect 48225 2907 48283 2913
rect 48225 2904 48237 2907
rect 47452 2876 48237 2904
rect 47452 2864 47458 2876
rect 48225 2873 48237 2876
rect 48271 2873 48283 2907
rect 48225 2867 48283 2873
rect 48774 2864 48780 2916
rect 48832 2904 48838 2916
rect 49513 2907 49571 2913
rect 49513 2904 49525 2907
rect 48832 2876 49525 2904
rect 48832 2864 48838 2876
rect 49513 2873 49525 2876
rect 49559 2873 49571 2907
rect 49513 2867 49571 2873
rect 49878 2864 49884 2916
rect 49936 2904 49942 2916
rect 50801 2907 50859 2913
rect 50801 2904 50813 2907
rect 49936 2876 50813 2904
rect 49936 2864 49942 2876
rect 50801 2873 50813 2876
rect 50847 2873 50859 2907
rect 50801 2867 50859 2873
rect 50982 2864 50988 2916
rect 51040 2904 51046 2916
rect 52733 2907 52791 2913
rect 52733 2904 52745 2907
rect 51040 2876 52745 2904
rect 51040 2864 51046 2876
rect 52733 2873 52745 2876
rect 52779 2873 52791 2907
rect 52733 2867 52791 2873
rect 54202 2864 54208 2916
rect 54260 2904 54266 2916
rect 57885 2907 57943 2913
rect 57885 2904 57897 2907
rect 54260 2876 57897 2904
rect 54260 2864 54266 2876
rect 57885 2873 57897 2876
rect 57931 2873 57943 2907
rect 57885 2867 57943 2873
rect 44968 2808 45140 2836
rect 44968 2796 44974 2808
rect 45462 2796 45468 2848
rect 45520 2836 45526 2848
rect 46293 2839 46351 2845
rect 46293 2836 46305 2839
rect 45520 2808 46305 2836
rect 45520 2796 45526 2808
rect 46293 2805 46305 2808
rect 46339 2805 46351 2839
rect 46293 2799 46351 2805
rect 46842 2796 46848 2848
rect 46900 2836 46906 2848
rect 47581 2839 47639 2845
rect 47581 2836 47593 2839
rect 46900 2808 47593 2836
rect 46900 2796 46906 2808
rect 47581 2805 47593 2808
rect 47627 2805 47639 2839
rect 47581 2799 47639 2805
rect 47946 2796 47952 2848
rect 48004 2836 48010 2848
rect 48869 2839 48927 2845
rect 48869 2836 48881 2839
rect 48004 2808 48881 2836
rect 48004 2796 48010 2808
rect 48869 2805 48881 2808
rect 48915 2805 48927 2839
rect 48869 2799 48927 2805
rect 49326 2796 49332 2848
rect 49384 2836 49390 2848
rect 50157 2839 50215 2845
rect 50157 2836 50169 2839
rect 49384 2808 50169 2836
rect 49384 2796 49390 2808
rect 50157 2805 50169 2808
rect 50203 2805 50215 2839
rect 50157 2799 50215 2805
rect 50706 2796 50712 2848
rect 50764 2836 50770 2848
rect 51445 2839 51503 2845
rect 51445 2836 51457 2839
rect 50764 2808 51457 2836
rect 50764 2796 50770 2808
rect 51445 2805 51457 2808
rect 51491 2805 51503 2839
rect 51445 2799 51503 2805
rect 51534 2796 51540 2848
rect 51592 2836 51598 2848
rect 53377 2839 53435 2845
rect 53377 2836 53389 2839
rect 51592 2808 53389 2836
rect 51592 2796 51598 2808
rect 53377 2805 53389 2808
rect 53423 2805 53435 2839
rect 53377 2799 53435 2805
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 1765 2635 1823 2641
rect 1765 2601 1777 2635
rect 1811 2632 1823 2635
rect 5166 2632 5172 2644
rect 1811 2604 5172 2632
rect 1811 2601 1823 2604
rect 1765 2595 1823 2601
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 5350 2592 5356 2644
rect 5408 2632 5414 2644
rect 5626 2632 5632 2644
rect 5408 2604 5632 2632
rect 5408 2592 5414 2604
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 6546 2592 6552 2644
rect 6604 2632 6610 2644
rect 6641 2635 6699 2641
rect 6641 2632 6653 2635
rect 6604 2604 6653 2632
rect 6604 2592 6610 2604
rect 6641 2601 6653 2604
rect 6687 2601 6699 2635
rect 10410 2632 10416 2644
rect 10371 2604 10416 2632
rect 6641 2595 6699 2601
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 11701 2635 11759 2641
rect 11701 2632 11713 2635
rect 11112 2604 11713 2632
rect 11112 2592 11118 2604
rect 11701 2601 11713 2604
rect 11747 2601 11759 2635
rect 13446 2632 13452 2644
rect 13407 2604 13452 2632
rect 11701 2595 11759 2601
rect 13446 2592 13452 2604
rect 13504 2592 13510 2644
rect 14550 2632 14556 2644
rect 14511 2604 14556 2632
rect 14550 2592 14556 2604
rect 14608 2592 14614 2644
rect 20346 2632 20352 2644
rect 20307 2604 20352 2632
rect 20346 2592 20352 2604
rect 20404 2592 20410 2644
rect 22741 2635 22799 2641
rect 22741 2601 22753 2635
rect 22787 2632 22799 2635
rect 22922 2632 22928 2644
rect 22787 2604 22928 2632
rect 22787 2601 22799 2604
rect 22741 2595 22799 2601
rect 22922 2592 22928 2604
rect 22980 2592 22986 2644
rect 26973 2635 27031 2641
rect 26973 2632 26985 2635
rect 23032 2604 26985 2632
rect 2038 2524 2044 2576
rect 2096 2564 2102 2576
rect 2225 2567 2283 2573
rect 2225 2564 2237 2567
rect 2096 2536 2237 2564
rect 2096 2524 2102 2536
rect 2225 2533 2237 2536
rect 2271 2533 2283 2567
rect 2225 2527 2283 2533
rect 3053 2567 3111 2573
rect 3053 2533 3065 2567
rect 3099 2564 3111 2567
rect 7374 2564 7380 2576
rect 3099 2536 7380 2564
rect 3099 2533 3111 2536
rect 3053 2527 3111 2533
rect 7374 2524 7380 2536
rect 7432 2524 7438 2576
rect 8570 2524 8576 2576
rect 8628 2564 8634 2576
rect 12437 2567 12495 2573
rect 12437 2564 12449 2567
rect 8628 2536 12449 2564
rect 8628 2524 8634 2536
rect 12437 2533 12449 2536
rect 12483 2533 12495 2567
rect 12437 2527 12495 2533
rect 16117 2567 16175 2573
rect 16117 2533 16129 2567
rect 16163 2564 16175 2567
rect 16206 2564 16212 2576
rect 16163 2536 16212 2564
rect 16163 2533 16175 2536
rect 16117 2527 16175 2533
rect 16206 2524 16212 2536
rect 16264 2524 16270 2576
rect 16853 2567 16911 2573
rect 16853 2533 16865 2567
rect 16899 2564 16911 2567
rect 17494 2564 17500 2576
rect 16899 2536 17500 2564
rect 16899 2533 16911 2536
rect 16853 2527 16911 2533
rect 17494 2524 17500 2536
rect 17552 2524 17558 2576
rect 17678 2564 17684 2576
rect 17639 2536 17684 2564
rect 17678 2524 17684 2536
rect 17736 2524 17742 2576
rect 18693 2567 18751 2573
rect 18693 2533 18705 2567
rect 18739 2564 18751 2567
rect 18782 2564 18788 2576
rect 18739 2536 18788 2564
rect 18739 2533 18751 2536
rect 18693 2527 18751 2533
rect 18782 2524 18788 2536
rect 18840 2524 18846 2576
rect 21266 2564 21272 2576
rect 21227 2536 21272 2564
rect 21266 2524 21272 2536
rect 21324 2524 21330 2576
rect 5258 2456 5264 2508
rect 5316 2496 5322 2508
rect 6546 2496 6552 2508
rect 5316 2468 6552 2496
rect 5316 2456 5322 2468
rect 6546 2456 6552 2468
rect 6604 2456 6610 2508
rect 7561 2499 7619 2505
rect 7561 2465 7573 2499
rect 7607 2496 7619 2499
rect 7926 2496 7932 2508
rect 7607 2468 7932 2496
rect 7607 2465 7619 2468
rect 7561 2459 7619 2465
rect 7926 2456 7932 2468
rect 7984 2456 7990 2508
rect 10962 2496 10968 2508
rect 9232 2468 10968 2496
rect 1578 2428 1584 2440
rect 1539 2400 1584 2428
rect 1578 2388 1584 2400
rect 1636 2388 1642 2440
rect 2409 2431 2467 2437
rect 2409 2397 2421 2431
rect 2455 2428 2467 2431
rect 2590 2428 2596 2440
rect 2455 2400 2596 2428
rect 2455 2397 2467 2400
rect 2409 2391 2467 2397
rect 2590 2388 2596 2400
rect 2648 2388 2654 2440
rect 3234 2428 3240 2440
rect 3195 2400 3240 2428
rect 3234 2388 3240 2400
rect 3292 2388 3298 2440
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2428 4307 2431
rect 4798 2428 4804 2440
rect 4295 2400 4804 2428
rect 4295 2397 4307 2400
rect 4249 2391 4307 2397
rect 4798 2388 4804 2400
rect 4856 2388 4862 2440
rect 5442 2388 5448 2440
rect 5500 2428 5506 2440
rect 5537 2431 5595 2437
rect 5537 2428 5549 2431
rect 5500 2400 5549 2428
rect 5500 2388 5506 2400
rect 5537 2397 5549 2400
rect 5583 2397 5595 2431
rect 5537 2391 5595 2397
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2428 5871 2431
rect 6178 2428 6184 2440
rect 5859 2400 6184 2428
rect 5859 2397 5871 2400
rect 5813 2391 5871 2397
rect 6178 2388 6184 2400
rect 6236 2388 6242 2440
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 9232 2437 9260 2468
rect 10962 2456 10968 2468
rect 11020 2456 11026 2508
rect 13630 2496 13636 2508
rect 12406 2468 13636 2496
rect 7285 2431 7343 2437
rect 7285 2428 7297 2431
rect 7248 2400 7297 2428
rect 7248 2388 7254 2400
rect 7285 2397 7297 2400
rect 7331 2397 7343 2431
rect 7285 2391 7343 2397
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2397 9275 2431
rect 9217 2391 9275 2397
rect 9582 2388 9588 2440
rect 9640 2428 9646 2440
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 9640 2400 10149 2428
rect 9640 2388 9646 2400
rect 10137 2397 10149 2400
rect 10183 2397 10195 2431
rect 11514 2428 11520 2440
rect 11475 2400 11520 2428
rect 10137 2391 10195 2397
rect 11514 2388 11520 2400
rect 11572 2388 11578 2440
rect 12253 2431 12311 2437
rect 12253 2397 12265 2431
rect 12299 2428 12311 2431
rect 12406 2428 12434 2468
rect 13630 2456 13636 2468
rect 13688 2456 13694 2508
rect 22370 2496 22376 2508
rect 15488 2468 22376 2496
rect 12299 2400 12434 2428
rect 12299 2397 12311 2400
rect 12253 2391 12311 2397
rect 13170 2388 13176 2440
rect 13228 2428 13234 2440
rect 13265 2431 13323 2437
rect 13265 2428 13277 2431
rect 13228 2400 13277 2428
rect 13228 2388 13234 2400
rect 13265 2397 13277 2400
rect 13311 2397 13323 2431
rect 13265 2391 13323 2397
rect 13906 2388 13912 2440
rect 13964 2428 13970 2440
rect 14369 2431 14427 2437
rect 14369 2428 14381 2431
rect 13964 2400 14381 2428
rect 13964 2388 13970 2400
rect 14369 2397 14381 2400
rect 14415 2428 14427 2431
rect 14550 2428 14556 2440
rect 14415 2400 14556 2428
rect 14415 2397 14427 2400
rect 14369 2391 14427 2397
rect 14550 2388 14556 2400
rect 14608 2388 14614 2440
rect 15102 2428 15108 2440
rect 15063 2400 15108 2428
rect 15102 2388 15108 2400
rect 15160 2388 15166 2440
rect 6733 2363 6791 2369
rect 4448 2332 6684 2360
rect 4448 2301 4476 2332
rect 4433 2295 4491 2301
rect 4433 2261 4445 2295
rect 4479 2261 4491 2295
rect 6656 2292 6684 2332
rect 6733 2329 6745 2363
rect 6779 2360 6791 2363
rect 8110 2360 8116 2372
rect 6779 2332 8116 2360
rect 6779 2329 6791 2332
rect 6733 2323 6791 2329
rect 8110 2320 8116 2332
rect 8168 2320 8174 2372
rect 8478 2320 8484 2372
rect 8536 2360 8542 2372
rect 9600 2360 9628 2388
rect 8536 2332 9628 2360
rect 8536 2320 8542 2332
rect 10410 2320 10416 2372
rect 10468 2360 10474 2372
rect 15488 2360 15516 2468
rect 22370 2456 22376 2468
rect 22428 2456 22434 2508
rect 23032 2440 23060 2604
rect 26973 2601 26985 2604
rect 27019 2601 27031 2635
rect 26973 2595 27031 2601
rect 51994 2592 52000 2644
rect 52052 2632 52058 2644
rect 55309 2635 55367 2641
rect 55309 2632 55321 2635
rect 52052 2604 55321 2632
rect 52052 2592 52058 2604
rect 55309 2601 55321 2604
rect 55355 2601 55367 2635
rect 55309 2595 55367 2601
rect 25777 2567 25835 2573
rect 25777 2533 25789 2567
rect 25823 2564 25835 2567
rect 26418 2564 26424 2576
rect 25823 2536 26424 2564
rect 25823 2533 25835 2536
rect 25777 2527 25835 2533
rect 26418 2524 26424 2536
rect 26476 2524 26482 2576
rect 27709 2567 27767 2573
rect 27709 2533 27721 2567
rect 27755 2564 27767 2567
rect 28350 2564 28356 2576
rect 27755 2536 28356 2564
rect 27755 2533 27767 2536
rect 27709 2527 27767 2533
rect 28350 2524 28356 2536
rect 28408 2524 28414 2576
rect 34146 2524 34152 2576
rect 34204 2564 34210 2576
rect 35989 2567 36047 2573
rect 35989 2564 36001 2567
rect 34204 2536 36001 2564
rect 34204 2524 34210 2536
rect 35989 2533 36001 2536
rect 36035 2533 36047 2567
rect 35989 2527 36047 2533
rect 38010 2524 38016 2576
rect 38068 2564 38074 2576
rect 39853 2567 39911 2573
rect 39853 2564 39865 2567
rect 38068 2536 39865 2564
rect 38068 2524 38074 2536
rect 39853 2533 39865 2536
rect 39899 2533 39911 2567
rect 39853 2527 39911 2533
rect 41874 2524 41880 2576
rect 41932 2564 41938 2576
rect 43717 2567 43775 2573
rect 43717 2564 43729 2567
rect 41932 2536 43729 2564
rect 41932 2524 41938 2536
rect 43717 2533 43729 2536
rect 43763 2533 43775 2567
rect 43717 2527 43775 2533
rect 45738 2524 45744 2576
rect 45796 2564 45802 2576
rect 47581 2567 47639 2573
rect 47581 2564 47593 2567
rect 45796 2536 47593 2564
rect 45796 2524 45802 2536
rect 47581 2533 47593 2536
rect 47627 2533 47639 2567
rect 47581 2527 47639 2533
rect 49602 2524 49608 2576
rect 49660 2564 49666 2576
rect 51445 2567 51503 2573
rect 51445 2564 51457 2567
rect 49660 2536 51457 2564
rect 49660 2524 49666 2536
rect 51445 2533 51457 2536
rect 51491 2533 51503 2567
rect 51445 2527 51503 2533
rect 54021 2567 54079 2573
rect 54021 2533 54033 2567
rect 54067 2533 54079 2567
rect 54021 2527 54079 2533
rect 31938 2456 31944 2508
rect 31996 2496 32002 2508
rect 32769 2499 32827 2505
rect 32769 2496 32781 2499
rect 31996 2468 32781 2496
rect 31996 2456 32002 2468
rect 32769 2465 32781 2468
rect 32815 2465 32827 2499
rect 32769 2459 32827 2465
rect 33042 2456 33048 2508
rect 33100 2496 33106 2508
rect 34701 2499 34759 2505
rect 34701 2496 34713 2499
rect 33100 2468 34713 2496
rect 33100 2456 33106 2468
rect 34701 2465 34713 2468
rect 34747 2465 34759 2499
rect 34701 2459 34759 2465
rect 35526 2456 35532 2508
rect 35584 2496 35590 2508
rect 37277 2499 37335 2505
rect 37277 2496 37289 2499
rect 35584 2468 37289 2496
rect 35584 2456 35590 2468
rect 37277 2465 37289 2468
rect 37323 2465 37335 2499
rect 37277 2459 37335 2465
rect 38838 2456 38844 2508
rect 38896 2496 38902 2508
rect 40497 2499 40555 2505
rect 40497 2496 40509 2499
rect 38896 2468 40509 2496
rect 38896 2456 38902 2468
rect 40497 2465 40509 2468
rect 40543 2465 40555 2499
rect 40497 2459 40555 2465
rect 40770 2456 40776 2508
rect 40828 2496 40834 2508
rect 42429 2499 42487 2505
rect 42429 2496 42441 2499
rect 40828 2468 42441 2496
rect 40828 2456 40834 2468
rect 42429 2465 42441 2468
rect 42475 2465 42487 2499
rect 42429 2459 42487 2465
rect 43254 2456 43260 2508
rect 43312 2496 43318 2508
rect 45005 2499 45063 2505
rect 45005 2496 45017 2499
rect 43312 2468 45017 2496
rect 43312 2456 43318 2468
rect 45005 2465 45017 2468
rect 45051 2465 45063 2499
rect 45005 2459 45063 2465
rect 46566 2456 46572 2508
rect 46624 2496 46630 2508
rect 48225 2499 48283 2505
rect 48225 2496 48237 2499
rect 46624 2468 48237 2496
rect 46624 2456 46630 2468
rect 48225 2465 48237 2468
rect 48271 2465 48283 2499
rect 48225 2459 48283 2465
rect 48498 2456 48504 2508
rect 48556 2496 48562 2508
rect 50157 2499 50215 2505
rect 50157 2496 50169 2499
rect 48556 2468 50169 2496
rect 48556 2456 48562 2468
rect 50157 2465 50169 2468
rect 50203 2465 50215 2499
rect 52733 2499 52791 2505
rect 52733 2496 52745 2499
rect 50157 2459 50215 2465
rect 51046 2468 52745 2496
rect 16669 2431 16727 2437
rect 16669 2397 16681 2431
rect 16715 2428 16727 2431
rect 16850 2428 16856 2440
rect 16715 2400 16856 2428
rect 16715 2397 16727 2400
rect 16669 2391 16727 2397
rect 16850 2388 16856 2400
rect 16908 2428 16914 2440
rect 17494 2428 17500 2440
rect 16908 2400 17500 2428
rect 16908 2388 16914 2400
rect 17494 2388 17500 2400
rect 17552 2388 17558 2440
rect 17865 2431 17923 2437
rect 17865 2397 17877 2431
rect 17911 2428 17923 2431
rect 19058 2428 19064 2440
rect 17911 2400 19064 2428
rect 17911 2397 17923 2400
rect 17865 2391 17923 2397
rect 19058 2388 19064 2400
rect 19116 2388 19122 2440
rect 19426 2388 19432 2440
rect 19484 2428 19490 2440
rect 19521 2431 19579 2437
rect 19521 2428 19533 2431
rect 19484 2400 19533 2428
rect 19484 2388 19490 2400
rect 19521 2397 19533 2400
rect 19567 2397 19579 2431
rect 22094 2428 22100 2440
rect 19521 2391 19579 2397
rect 20364 2400 22100 2428
rect 20364 2372 20392 2400
rect 22094 2388 22100 2400
rect 22152 2388 22158 2440
rect 22189 2431 22247 2437
rect 22189 2397 22201 2431
rect 22235 2428 22247 2431
rect 22646 2428 22652 2440
rect 22235 2400 22652 2428
rect 22235 2397 22247 2400
rect 22189 2391 22247 2397
rect 22646 2388 22652 2400
rect 22704 2388 22710 2440
rect 22925 2431 22983 2437
rect 22925 2397 22937 2431
rect 22971 2428 22983 2431
rect 23014 2428 23020 2440
rect 22971 2400 23020 2428
rect 22971 2397 22983 2400
rect 22925 2391 22983 2397
rect 23014 2388 23020 2400
rect 23072 2388 23078 2440
rect 23290 2388 23296 2440
rect 23348 2428 23354 2440
rect 23385 2431 23443 2437
rect 23385 2428 23397 2431
rect 23348 2400 23397 2428
rect 23348 2388 23354 2400
rect 23385 2397 23397 2400
rect 23431 2428 23443 2431
rect 24397 2431 24455 2437
rect 24397 2428 24409 2431
rect 23431 2400 24409 2428
rect 23431 2397 23443 2400
rect 23385 2391 23443 2397
rect 24397 2397 24409 2400
rect 24443 2397 24455 2431
rect 24397 2391 24455 2397
rect 25133 2431 25191 2437
rect 25133 2397 25145 2431
rect 25179 2428 25191 2431
rect 25866 2428 25872 2440
rect 25179 2400 25872 2428
rect 25179 2397 25191 2400
rect 25133 2391 25191 2397
rect 25866 2388 25872 2400
rect 25924 2388 25930 2440
rect 26421 2431 26479 2437
rect 26421 2397 26433 2431
rect 26467 2428 26479 2431
rect 27246 2428 27252 2440
rect 26467 2400 27252 2428
rect 26467 2397 26479 2400
rect 26421 2391 26479 2397
rect 27246 2388 27252 2400
rect 27304 2388 27310 2440
rect 28353 2431 28411 2437
rect 27356 2400 27752 2428
rect 10468 2332 15516 2360
rect 15933 2363 15991 2369
rect 10468 2320 10474 2332
rect 15933 2329 15945 2363
rect 15979 2360 15991 2363
rect 17954 2360 17960 2372
rect 15979 2332 17960 2360
rect 15979 2329 15991 2332
rect 15933 2323 15991 2329
rect 17954 2320 17960 2332
rect 18012 2320 18018 2372
rect 18509 2363 18567 2369
rect 18509 2329 18521 2363
rect 18555 2360 18567 2363
rect 20346 2360 20352 2372
rect 18555 2332 20352 2360
rect 18555 2329 18567 2332
rect 18509 2323 18567 2329
rect 20346 2320 20352 2332
rect 20404 2320 20410 2372
rect 20441 2363 20499 2369
rect 20441 2329 20453 2363
rect 20487 2360 20499 2363
rect 20714 2360 20720 2372
rect 20487 2332 20720 2360
rect 20487 2329 20499 2332
rect 20441 2323 20499 2329
rect 20714 2320 20720 2332
rect 20772 2320 20778 2372
rect 21085 2363 21143 2369
rect 21085 2329 21097 2363
rect 21131 2360 21143 2363
rect 21910 2360 21916 2372
rect 21131 2332 21916 2360
rect 21131 2329 21143 2332
rect 21085 2323 21143 2329
rect 21910 2320 21916 2332
rect 21968 2320 21974 2372
rect 27356 2360 27384 2400
rect 22020 2332 27384 2360
rect 27724 2360 27752 2400
rect 28353 2397 28365 2431
rect 28399 2428 28411 2431
rect 28902 2428 28908 2440
rect 28399 2400 28908 2428
rect 28399 2397 28411 2400
rect 28353 2391 28411 2397
rect 28902 2388 28908 2400
rect 28960 2388 28966 2440
rect 28997 2431 29055 2437
rect 28997 2397 29009 2431
rect 29043 2428 29055 2431
rect 29454 2428 29460 2440
rect 29043 2400 29460 2428
rect 29043 2397 29055 2400
rect 28997 2391 29055 2397
rect 29454 2388 29460 2400
rect 29512 2388 29518 2440
rect 30101 2431 30159 2437
rect 30101 2397 30113 2431
rect 30147 2428 30159 2431
rect 30282 2428 30288 2440
rect 30147 2400 30288 2428
rect 30147 2397 30159 2400
rect 30101 2391 30159 2397
rect 30282 2388 30288 2400
rect 30340 2388 30346 2440
rect 30745 2431 30803 2437
rect 30745 2397 30757 2431
rect 30791 2428 30803 2431
rect 30834 2428 30840 2440
rect 30791 2400 30840 2428
rect 30791 2397 30803 2400
rect 30745 2391 30803 2397
rect 30834 2388 30840 2400
rect 30892 2388 30898 2440
rect 31110 2388 31116 2440
rect 31168 2428 31174 2440
rect 31205 2431 31263 2437
rect 31205 2428 31217 2431
rect 31168 2400 31217 2428
rect 31168 2388 31174 2400
rect 31205 2397 31217 2400
rect 31251 2397 31263 2431
rect 31205 2391 31263 2397
rect 31386 2388 31392 2440
rect 31444 2428 31450 2440
rect 32125 2431 32183 2437
rect 32125 2428 32137 2431
rect 31444 2400 32137 2428
rect 31444 2388 31450 2400
rect 32125 2397 32137 2400
rect 32171 2397 32183 2431
rect 32125 2391 32183 2397
rect 32490 2388 32496 2440
rect 32548 2428 32554 2440
rect 33413 2431 33471 2437
rect 33413 2428 33425 2431
rect 32548 2400 33425 2428
rect 32548 2388 32554 2400
rect 33413 2397 33425 2400
rect 33459 2397 33471 2431
rect 33413 2391 33471 2397
rect 33594 2388 33600 2440
rect 33652 2428 33658 2440
rect 35345 2431 35403 2437
rect 35345 2428 35357 2431
rect 33652 2400 35357 2428
rect 33652 2388 33658 2400
rect 35345 2397 35357 2400
rect 35391 2397 35403 2431
rect 35345 2391 35403 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 37921 2431 37979 2437
rect 37921 2428 37933 2431
rect 36136 2400 37933 2428
rect 36136 2388 36142 2400
rect 37921 2397 37933 2400
rect 37967 2397 37979 2431
rect 37921 2391 37979 2397
rect 38565 2431 38623 2437
rect 38565 2397 38577 2431
rect 38611 2397 38623 2431
rect 38565 2391 38623 2397
rect 27724 2332 35894 2360
rect 7742 2292 7748 2304
rect 6656 2264 7748 2292
rect 4433 2255 4491 2261
rect 7742 2252 7748 2264
rect 7800 2252 7806 2304
rect 8846 2252 8852 2304
rect 8904 2292 8910 2304
rect 9033 2295 9091 2301
rect 9033 2292 9045 2295
rect 8904 2264 9045 2292
rect 8904 2252 8910 2264
rect 9033 2261 9045 2264
rect 9079 2261 9091 2295
rect 15286 2292 15292 2304
rect 15247 2264 15292 2292
rect 9033 2255 9091 2261
rect 15286 2252 15292 2264
rect 15344 2252 15350 2304
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 22020 2301 22048 2332
rect 19337 2295 19395 2301
rect 19337 2292 19349 2295
rect 17460 2264 19349 2292
rect 17460 2252 17466 2264
rect 19337 2261 19349 2264
rect 19383 2261 19395 2295
rect 19337 2255 19395 2261
rect 22005 2295 22063 2301
rect 22005 2261 22017 2295
rect 22051 2261 22063 2295
rect 22005 2255 22063 2261
rect 23569 2295 23627 2301
rect 23569 2261 23581 2295
rect 23615 2292 23627 2295
rect 35710 2292 35716 2304
rect 23615 2264 35716 2292
rect 23615 2261 23627 2264
rect 23569 2255 23627 2261
rect 35710 2252 35716 2264
rect 35768 2252 35774 2304
rect 35866 2292 35894 2332
rect 36906 2320 36912 2372
rect 36964 2360 36970 2372
rect 38580 2360 38608 2391
rect 39390 2388 39396 2440
rect 39448 2428 39454 2440
rect 41141 2431 41199 2437
rect 41141 2428 41153 2431
rect 39448 2400 41153 2428
rect 39448 2388 39454 2400
rect 41141 2397 41153 2400
rect 41187 2397 41199 2431
rect 41141 2391 41199 2397
rect 41322 2388 41328 2440
rect 41380 2428 41386 2440
rect 43073 2431 43131 2437
rect 43073 2428 43085 2431
rect 41380 2400 43085 2428
rect 41380 2388 41386 2400
rect 43073 2397 43085 2400
rect 43119 2397 43131 2431
rect 43073 2391 43131 2397
rect 43806 2388 43812 2440
rect 43864 2428 43870 2440
rect 45649 2431 45707 2437
rect 45649 2428 45661 2431
rect 43864 2400 45661 2428
rect 43864 2388 43870 2400
rect 45649 2397 45661 2400
rect 45695 2397 45707 2431
rect 45649 2391 45707 2397
rect 46293 2431 46351 2437
rect 46293 2397 46305 2431
rect 46339 2397 46351 2431
rect 46293 2391 46351 2397
rect 36964 2332 38608 2360
rect 36964 2320 36970 2332
rect 44634 2320 44640 2372
rect 44692 2360 44698 2372
rect 46308 2360 46336 2391
rect 47118 2388 47124 2440
rect 47176 2428 47182 2440
rect 48869 2431 48927 2437
rect 48869 2428 48881 2431
rect 47176 2400 48881 2428
rect 47176 2388 47182 2400
rect 48869 2397 48881 2400
rect 48915 2397 48927 2431
rect 48869 2391 48927 2397
rect 49050 2388 49056 2440
rect 49108 2428 49114 2440
rect 50801 2431 50859 2437
rect 50801 2428 50813 2431
rect 49108 2400 50813 2428
rect 49108 2388 49114 2400
rect 50801 2397 50813 2400
rect 50847 2397 50859 2431
rect 50801 2391 50859 2397
rect 50890 2388 50896 2440
rect 50948 2428 50954 2440
rect 51046 2428 51074 2468
rect 52733 2465 52745 2468
rect 52779 2465 52791 2499
rect 54036 2496 54064 2527
rect 57882 2496 57888 2508
rect 54036 2468 54156 2496
rect 57843 2468 57888 2496
rect 52733 2459 52791 2465
rect 50948 2400 51074 2428
rect 50948 2388 50954 2400
rect 52546 2388 52552 2440
rect 52604 2428 52610 2440
rect 53377 2431 53435 2437
rect 53377 2428 53389 2431
rect 52604 2400 53389 2428
rect 52604 2388 52610 2400
rect 53377 2397 53389 2400
rect 53423 2397 53435 2431
rect 53377 2391 53435 2397
rect 44692 2332 46336 2360
rect 44692 2320 44698 2332
rect 46750 2292 46756 2304
rect 35866 2264 46756 2292
rect 46750 2252 46756 2264
rect 46808 2252 46814 2304
rect 51258 2252 51264 2304
rect 51316 2292 51322 2304
rect 54128 2292 54156 2468
rect 57882 2456 57888 2468
rect 57940 2456 57946 2508
rect 55950 2428 55956 2440
rect 55911 2400 55956 2428
rect 55950 2388 55956 2400
rect 56008 2388 56014 2440
rect 56594 2428 56600 2440
rect 56555 2400 56600 2428
rect 56594 2388 56600 2400
rect 56652 2388 56658 2440
rect 51316 2264 54156 2292
rect 51316 2252 51322 2264
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 14550 2048 14556 2100
rect 14608 2088 14614 2100
rect 16114 2088 16120 2100
rect 14608 2060 16120 2088
rect 14608 2048 14614 2060
rect 16114 2048 16120 2060
rect 16172 2048 16178 2100
rect 18874 2048 18880 2100
rect 18932 2088 18938 2100
rect 19610 2088 19616 2100
rect 18932 2060 19616 2088
rect 18932 2048 18938 2060
rect 19610 2048 19616 2060
rect 19668 2048 19674 2100
rect 25130 2088 25136 2100
rect 22066 2060 25136 2088
rect 5442 1980 5448 2032
rect 5500 2020 5506 2032
rect 10042 2020 10048 2032
rect 5500 1992 10048 2020
rect 5500 1980 5506 1992
rect 10042 1980 10048 1992
rect 10100 1980 10106 2032
rect 15286 1980 15292 2032
rect 15344 2020 15350 2032
rect 22066 2020 22094 2060
rect 25130 2048 25136 2060
rect 25188 2048 25194 2100
rect 52362 2048 52368 2100
rect 52420 2088 52426 2100
rect 55950 2088 55956 2100
rect 52420 2060 55956 2088
rect 52420 2048 52426 2060
rect 55950 2048 55956 2060
rect 56008 2048 56014 2100
rect 15344 1992 22094 2020
rect 15344 1980 15350 1992
rect 22462 1980 22468 2032
rect 22520 2020 22526 2032
rect 22646 2020 22652 2032
rect 22520 1992 22652 2020
rect 22520 1980 22526 1992
rect 22646 1980 22652 1992
rect 22704 1980 22710 2032
rect 53558 1980 53564 2032
rect 53616 2020 53622 2032
rect 57882 2020 57888 2032
rect 53616 1992 57888 2020
rect 53616 1980 53622 1992
rect 57882 1980 57888 1992
rect 57940 1980 57946 2032
rect 4062 1912 4068 1964
rect 4120 1952 4126 1964
rect 11514 1952 11520 1964
rect 4120 1924 11520 1952
rect 4120 1912 4126 1924
rect 11514 1912 11520 1924
rect 11572 1912 11578 1964
rect 22370 1912 22376 1964
rect 22428 1952 22434 1964
rect 29546 1952 29552 1964
rect 22428 1924 29552 1952
rect 22428 1912 22434 1924
rect 29546 1912 29552 1924
rect 29604 1912 29610 1964
rect 7926 1844 7932 1896
rect 7984 1884 7990 1896
rect 8110 1884 8116 1896
rect 7984 1856 8116 1884
rect 7984 1844 7990 1856
rect 8110 1844 8116 1856
rect 8168 1844 8174 1896
rect 13170 1844 13176 1896
rect 13228 1884 13234 1896
rect 15286 1884 15292 1896
rect 13228 1856 15292 1884
rect 13228 1844 13234 1856
rect 15286 1844 15292 1856
rect 15344 1844 15350 1896
rect 18874 1708 18880 1760
rect 18932 1748 18938 1760
rect 19058 1748 19064 1760
rect 18932 1720 19064 1748
rect 18932 1708 18938 1720
rect 19058 1708 19064 1720
rect 19116 1708 19122 1760
rect 20714 1708 20720 1760
rect 20772 1748 20778 1760
rect 21082 1748 21088 1760
rect 20772 1720 21088 1748
rect 20772 1708 20778 1720
rect 21082 1708 21088 1720
rect 21140 1708 21146 1760
rect 20254 1504 20260 1556
rect 20312 1504 20318 1556
rect 1578 1436 1584 1488
rect 1636 1476 1642 1488
rect 8110 1476 8116 1488
rect 1636 1448 8116 1476
rect 1636 1436 1642 1448
rect 8110 1436 8116 1448
rect 8168 1436 8174 1488
rect 15562 1300 15568 1352
rect 15620 1340 15626 1352
rect 16022 1340 16028 1352
rect 15620 1312 16028 1340
rect 15620 1300 15626 1312
rect 16022 1300 16028 1312
rect 16080 1300 16086 1352
rect 19518 1300 19524 1352
rect 19576 1340 19582 1352
rect 19794 1340 19800 1352
rect 19576 1312 19800 1340
rect 19576 1300 19582 1312
rect 19794 1300 19800 1312
rect 19852 1300 19858 1352
rect 19978 1300 19984 1352
rect 20036 1340 20042 1352
rect 20272 1340 20300 1504
rect 52730 1368 52736 1420
rect 52788 1408 52794 1420
rect 53006 1408 53012 1420
rect 52788 1380 53012 1408
rect 52788 1368 52794 1380
rect 53006 1368 53012 1380
rect 53064 1368 53070 1420
rect 56594 1408 56600 1420
rect 53116 1380 56600 1408
rect 20036 1312 20300 1340
rect 20036 1300 20042 1312
rect 19426 1164 19432 1216
rect 19484 1164 19490 1216
rect 19444 944 19472 1164
rect 52546 1136 52552 1148
rect 51000 1108 52552 1136
rect 20162 1028 20168 1080
rect 20220 1068 20226 1080
rect 20346 1068 20352 1080
rect 20220 1040 20352 1068
rect 20220 1028 20226 1040
rect 20346 1028 20352 1040
rect 20404 1028 20410 1080
rect 51000 944 51028 1108
rect 52546 1096 52552 1108
rect 52604 1096 52610 1148
rect 6178 892 6184 944
rect 6236 932 6242 944
rect 6730 932 6736 944
rect 6236 904 6736 932
rect 6236 892 6242 904
rect 6730 892 6736 904
rect 6788 892 6794 944
rect 19426 892 19432 944
rect 19484 892 19490 944
rect 50982 892 50988 944
rect 51040 892 51046 944
rect 52546 892 52552 944
rect 52604 892 52610 944
rect 52914 892 52920 944
rect 52972 932 52978 944
rect 53116 932 53144 1380
rect 56594 1368 56600 1380
rect 56652 1368 56658 1420
rect 52972 904 53144 932
rect 52972 892 52978 904
rect 52564 864 52592 892
rect 54754 864 54760 876
rect 52564 836 54760 864
rect 54754 824 54760 836
rect 54812 824 54818 876
<< via1 >>
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 1768 57536 1820 57588
rect 3332 57536 3384 57588
rect 4896 57536 4948 57588
rect 6460 57536 6512 57588
rect 8024 57536 8076 57588
rect 9680 57536 9732 57588
rect 11152 57536 11204 57588
rect 12716 57536 12768 57588
rect 14280 57536 14332 57588
rect 15844 57536 15896 57588
rect 17408 57536 17460 57588
rect 19340 57536 19392 57588
rect 20720 57536 20772 57588
rect 22100 57536 22152 57588
rect 23664 57536 23716 57588
rect 25228 57536 25280 57588
rect 26792 57536 26844 57588
rect 28356 57536 28408 57588
rect 29920 57536 29972 57588
rect 31484 57536 31536 57588
rect 33140 57536 33192 57588
rect 34612 57536 34664 57588
rect 36176 57536 36228 57588
rect 37740 57536 37792 57588
rect 39304 57536 39356 57588
rect 40868 57536 40920 57588
rect 42432 57536 42484 57588
rect 44180 57536 44232 57588
rect 45560 57536 45612 57588
rect 47124 57536 47176 57588
rect 26332 57468 26384 57520
rect 2688 57400 2740 57452
rect 4068 57443 4120 57452
rect 4068 57409 4077 57443
rect 4077 57409 4111 57443
rect 4111 57409 4120 57443
rect 4068 57400 4120 57409
rect 5264 57443 5316 57452
rect 5264 57409 5273 57443
rect 5273 57409 5307 57443
rect 5307 57409 5316 57443
rect 5264 57400 5316 57409
rect 6828 57443 6880 57452
rect 6828 57409 6837 57443
rect 6837 57409 6871 57443
rect 6871 57409 6880 57443
rect 6828 57400 6880 57409
rect 11796 57443 11848 57452
rect 11796 57409 11805 57443
rect 11805 57409 11839 57443
rect 11839 57409 11848 57443
rect 11796 57400 11848 57409
rect 13084 57443 13136 57452
rect 13084 57409 13093 57443
rect 13093 57409 13127 57443
rect 13127 57409 13136 57443
rect 13084 57400 13136 57409
rect 15752 57400 15804 57452
rect 16948 57443 17000 57452
rect 16948 57409 16957 57443
rect 16957 57409 16991 57443
rect 16991 57409 17000 57443
rect 16948 57400 17000 57409
rect 17500 57443 17552 57452
rect 17500 57409 17509 57443
rect 17509 57409 17543 57443
rect 17543 57409 17552 57443
rect 17500 57400 17552 57409
rect 18696 57400 18748 57452
rect 19524 57400 19576 57452
rect 22192 57443 22244 57452
rect 22192 57409 22201 57443
rect 22201 57409 22235 57443
rect 22235 57409 22244 57443
rect 22192 57400 22244 57409
rect 24400 57443 24452 57452
rect 24400 57409 24409 57443
rect 24409 57409 24443 57443
rect 24443 57409 24452 57443
rect 24400 57400 24452 57409
rect 25320 57443 25372 57452
rect 25320 57409 25329 57443
rect 25329 57409 25363 57443
rect 25363 57409 25372 57443
rect 25320 57400 25372 57409
rect 26976 57443 27028 57452
rect 26976 57409 26985 57443
rect 26985 57409 27019 57443
rect 27019 57409 27028 57443
rect 26976 57400 27028 57409
rect 28448 57443 28500 57452
rect 28448 57409 28457 57443
rect 28457 57409 28491 57443
rect 28491 57409 28500 57443
rect 28448 57400 28500 57409
rect 30380 57468 30432 57520
rect 30104 57400 30156 57452
rect 32220 57400 32272 57452
rect 33232 57400 33284 57452
rect 19984 57332 20036 57384
rect 18512 57264 18564 57316
rect 24676 57264 24728 57316
rect 37188 57264 37240 57316
rect 40776 57400 40828 57452
rect 42524 57443 42576 57452
rect 42524 57409 42533 57443
rect 42533 57409 42567 57443
rect 42567 57409 42576 57443
rect 42524 57400 42576 57409
rect 44088 57443 44140 57452
rect 44088 57409 44097 57443
rect 44097 57409 44131 57443
rect 44131 57409 44140 57443
rect 44088 57400 44140 57409
rect 44180 57400 44232 57452
rect 47584 57443 47636 57452
rect 47584 57409 47593 57443
rect 47593 57409 47627 57443
rect 47627 57409 47636 57443
rect 47584 57400 47636 57409
rect 48688 57400 48740 57452
rect 50160 57400 50212 57452
rect 51816 57400 51868 57452
rect 53380 57400 53432 57452
rect 56600 57443 56652 57452
rect 56600 57409 56609 57443
rect 56609 57409 56643 57443
rect 56643 57409 56652 57443
rect 56600 57400 56652 57409
rect 58072 57400 58124 57452
rect 54944 57332 54996 57384
rect 2688 57239 2740 57248
rect 2688 57205 2697 57239
rect 2697 57205 2731 57239
rect 2731 57205 2740 57239
rect 2688 57196 2740 57205
rect 18972 57196 19024 57248
rect 20168 57196 20220 57248
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 18696 57035 18748 57044
rect 18696 57001 18705 57035
rect 18705 57001 18739 57035
rect 18739 57001 18748 57035
rect 18696 56992 18748 57001
rect 19524 57035 19576 57044
rect 19524 57001 19533 57035
rect 19533 57001 19567 57035
rect 19567 57001 19576 57035
rect 19524 56992 19576 57001
rect 19984 57035 20036 57044
rect 19984 57001 19993 57035
rect 19993 57001 20027 57035
rect 20027 57001 20036 57035
rect 19984 56992 20036 57001
rect 57520 57035 57572 57044
rect 57520 57001 57529 57035
rect 57529 57001 57563 57035
rect 57563 57001 57572 57035
rect 57520 56992 57572 57001
rect 6828 56924 6880 56976
rect 18788 56924 18840 56976
rect 19340 56924 19392 56976
rect 11796 56856 11848 56908
rect 1400 56831 1452 56840
rect 1400 56797 1409 56831
rect 1409 56797 1443 56831
rect 1443 56797 1452 56831
rect 1400 56788 1452 56797
rect 18144 56788 18196 56840
rect 20168 56831 20220 56840
rect 19064 56720 19116 56772
rect 20168 56797 20177 56831
rect 20177 56797 20211 56831
rect 20211 56797 20220 56831
rect 20168 56788 20220 56797
rect 57888 56788 57940 56840
rect 20720 56695 20772 56704
rect 20720 56661 20729 56695
rect 20729 56661 20763 56695
rect 20763 56661 20772 56695
rect 20720 56652 20772 56661
rect 23388 56652 23440 56704
rect 42524 56720 42576 56772
rect 40776 56695 40828 56704
rect 40776 56661 40785 56695
rect 40785 56661 40819 56695
rect 40819 56661 40828 56695
rect 40776 56652 40828 56661
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 13084 56448 13136 56500
rect 15752 56491 15804 56500
rect 15752 56457 15761 56491
rect 15761 56457 15795 56491
rect 15795 56457 15804 56491
rect 15752 56448 15804 56457
rect 17500 56491 17552 56500
rect 17500 56457 17509 56491
rect 17509 56457 17543 56491
rect 17543 56457 17552 56491
rect 17500 56448 17552 56457
rect 18788 56491 18840 56500
rect 18788 56457 18797 56491
rect 18797 56457 18831 56491
rect 18831 56457 18840 56491
rect 18788 56448 18840 56457
rect 22192 56448 22244 56500
rect 24400 56448 24452 56500
rect 24676 56491 24728 56500
rect 24676 56457 24685 56491
rect 24685 56457 24719 56491
rect 24719 56457 24728 56491
rect 24676 56448 24728 56457
rect 26332 56448 26384 56500
rect 26976 56448 27028 56500
rect 28448 56448 28500 56500
rect 30104 56448 30156 56500
rect 32220 56448 32272 56500
rect 33232 56448 33284 56500
rect 37188 56448 37240 56500
rect 44180 56448 44232 56500
rect 47584 56448 47636 56500
rect 14188 56312 14240 56364
rect 15936 56355 15988 56364
rect 15936 56321 15945 56355
rect 15945 56321 15979 56355
rect 15979 56321 15988 56355
rect 15936 56312 15988 56321
rect 17684 56355 17736 56364
rect 17684 56321 17693 56355
rect 17693 56321 17727 56355
rect 17727 56321 17736 56355
rect 17684 56312 17736 56321
rect 19432 56380 19484 56432
rect 18880 56312 18932 56364
rect 18972 56355 19024 56364
rect 18972 56321 18981 56355
rect 18981 56321 19015 56355
rect 19015 56321 19024 56355
rect 18972 56312 19024 56321
rect 19984 56312 20036 56364
rect 20720 56380 20772 56432
rect 20904 56312 20956 56364
rect 21732 56312 21784 56364
rect 22560 56355 22612 56364
rect 22560 56321 22569 56355
rect 22569 56321 22603 56355
rect 22603 56321 22612 56355
rect 22560 56312 22612 56321
rect 23020 56312 23072 56364
rect 23756 56312 23808 56364
rect 24400 56312 24452 56364
rect 25136 56355 25188 56364
rect 25136 56321 25145 56355
rect 25145 56321 25179 56355
rect 25179 56321 25188 56355
rect 25136 56312 25188 56321
rect 26056 56312 26108 56364
rect 26792 56312 26844 56364
rect 27988 56312 28040 56364
rect 29184 56355 29236 56364
rect 29184 56321 29193 56355
rect 29193 56321 29227 56355
rect 29227 56321 29236 56355
rect 29184 56312 29236 56321
rect 29920 56312 29972 56364
rect 30932 56312 30984 56364
rect 32128 56355 32180 56364
rect 32128 56321 32137 56355
rect 32137 56321 32171 56355
rect 32171 56321 32180 56355
rect 32128 56312 32180 56321
rect 35716 56312 35768 56364
rect 43812 56355 43864 56364
rect 43812 56321 43821 56355
rect 43821 56321 43855 56355
rect 43855 56321 43864 56355
rect 43812 56312 43864 56321
rect 46756 56312 46808 56364
rect 58440 56312 58492 56364
rect 5264 56244 5316 56296
rect 4068 56176 4120 56228
rect 20168 56244 20220 56296
rect 14188 56151 14240 56160
rect 14188 56117 14197 56151
rect 14197 56117 14231 56151
rect 14231 56117 14240 56151
rect 14188 56108 14240 56117
rect 40776 56244 40828 56296
rect 29920 56219 29972 56228
rect 29920 56185 29929 56219
rect 29929 56185 29963 56219
rect 29963 56185 29972 56219
rect 29920 56176 29972 56185
rect 44088 56176 44140 56228
rect 20076 56151 20128 56160
rect 20076 56117 20085 56151
rect 20085 56117 20119 56151
rect 20119 56117 20128 56151
rect 20076 56108 20128 56117
rect 23388 56151 23440 56160
rect 23388 56117 23397 56151
rect 23397 56117 23431 56151
rect 23431 56117 23440 56151
rect 23388 56108 23440 56117
rect 25320 56108 25372 56160
rect 27988 56151 28040 56160
rect 27988 56117 27997 56151
rect 27997 56117 28031 56151
rect 28031 56117 28040 56151
rect 27988 56108 28040 56117
rect 30380 56108 30432 56160
rect 46756 56151 46808 56160
rect 46756 56117 46765 56151
rect 46765 56117 46799 56151
rect 46799 56117 46808 56151
rect 46756 56108 46808 56117
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 2688 55904 2740 55956
rect 20076 55904 20128 55956
rect 16948 55836 17000 55888
rect 18512 55879 18564 55888
rect 18512 55845 18521 55879
rect 18521 55845 18555 55879
rect 18555 55845 18564 55879
rect 18512 55836 18564 55845
rect 19340 55836 19392 55888
rect 20076 55768 20128 55820
rect 22560 55768 22612 55820
rect 1400 55743 1452 55752
rect 1400 55709 1409 55743
rect 1409 55709 1443 55743
rect 1443 55709 1452 55743
rect 1400 55700 1452 55709
rect 17776 55700 17828 55752
rect 18788 55700 18840 55752
rect 15936 55564 15988 55616
rect 16488 55564 16540 55616
rect 17040 55607 17092 55616
rect 17040 55573 17049 55607
rect 17049 55573 17083 55607
rect 17083 55573 17092 55607
rect 17040 55564 17092 55573
rect 20260 55607 20312 55616
rect 20260 55573 20269 55607
rect 20269 55573 20303 55607
rect 20303 55573 20312 55607
rect 20260 55564 20312 55573
rect 20904 55607 20956 55616
rect 20904 55573 20913 55607
rect 20913 55573 20947 55607
rect 20947 55573 20956 55607
rect 20904 55564 20956 55573
rect 21732 55607 21784 55616
rect 21732 55573 21741 55607
rect 21741 55573 21775 55607
rect 21775 55573 21784 55607
rect 21732 55564 21784 55573
rect 23020 55607 23072 55616
rect 23020 55573 23029 55607
rect 23029 55573 23063 55607
rect 23063 55573 23072 55607
rect 23020 55564 23072 55573
rect 23756 55607 23808 55616
rect 23756 55573 23765 55607
rect 23765 55573 23799 55607
rect 23799 55573 23808 55607
rect 23756 55564 23808 55573
rect 24400 55607 24452 55616
rect 24400 55573 24409 55607
rect 24409 55573 24443 55607
rect 24443 55573 24452 55607
rect 24400 55564 24452 55573
rect 25136 55564 25188 55616
rect 26056 55607 26108 55616
rect 26056 55573 26065 55607
rect 26065 55573 26099 55607
rect 26099 55573 26108 55607
rect 26056 55564 26108 55573
rect 26792 55607 26844 55616
rect 26792 55573 26801 55607
rect 26801 55573 26835 55607
rect 26835 55573 26844 55607
rect 26792 55564 26844 55573
rect 29184 55564 29236 55616
rect 30932 55607 30984 55616
rect 30932 55573 30941 55607
rect 30941 55573 30975 55607
rect 30975 55573 30984 55607
rect 30932 55564 30984 55573
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 17776 55335 17828 55344
rect 17776 55301 17785 55335
rect 17785 55301 17819 55335
rect 17819 55301 17828 55335
rect 17776 55292 17828 55301
rect 18788 55335 18840 55344
rect 18788 55301 18797 55335
rect 18797 55301 18831 55335
rect 18831 55301 18840 55335
rect 18788 55292 18840 55301
rect 19800 55335 19852 55344
rect 19800 55301 19809 55335
rect 19809 55301 19843 55335
rect 19843 55301 19852 55335
rect 19800 55292 19852 55301
rect 19984 55292 20036 55344
rect 58164 55131 58216 55140
rect 58164 55097 58173 55131
rect 58173 55097 58207 55131
rect 58207 55097 58216 55131
rect 58164 55088 58216 55097
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 1400 54655 1452 54664
rect 1400 54621 1409 54655
rect 1409 54621 1443 54655
rect 1443 54621 1452 54655
rect 1400 54612 1452 54621
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 57888 53932 57940 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 1400 53567 1452 53576
rect 1400 53533 1409 53567
rect 1409 53533 1443 53567
rect 1443 53533 1452 53567
rect 1400 53524 1452 53533
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 1400 52479 1452 52488
rect 1400 52445 1409 52479
rect 1409 52445 1443 52479
rect 1443 52445 1452 52479
rect 1400 52436 1452 52445
rect 57888 52436 57940 52488
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 1400 51391 1452 51400
rect 1400 51357 1409 51391
rect 1409 51357 1443 51391
rect 1443 51357 1452 51391
rect 1400 51348 1452 51357
rect 58164 51391 58216 51400
rect 58164 51357 58173 51391
rect 58173 51357 58207 51391
rect 58207 51357 58216 51391
rect 58164 51348 58216 51357
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 16212 50328 16264 50380
rect 20904 50328 20956 50380
rect 1400 50303 1452 50312
rect 1400 50269 1409 50303
rect 1409 50269 1443 50303
rect 1443 50269 1452 50303
rect 1400 50260 1452 50269
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 58164 49759 58216 49768
rect 58164 49725 58173 49759
rect 58173 49725 58207 49759
rect 58207 49725 58216 49759
rect 58164 49716 58216 49725
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 1400 49215 1452 49224
rect 1400 49181 1409 49215
rect 1409 49181 1443 49215
rect 1443 49181 1452 49215
rect 1400 49172 1452 49181
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 58164 48535 58216 48544
rect 58164 48501 58173 48535
rect 58173 48501 58207 48535
rect 58207 48501 58216 48535
rect 58164 48492 58216 48501
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 1400 48127 1452 48136
rect 1400 48093 1409 48127
rect 1409 48093 1443 48127
rect 1443 48093 1452 48127
rect 1400 48084 1452 48093
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 58164 47039 58216 47048
rect 58164 47005 58173 47039
rect 58173 47005 58207 47039
rect 58207 47005 58216 47039
rect 58164 46996 58216 47005
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 58164 45951 58216 45960
rect 58164 45917 58173 45951
rect 58173 45917 58207 45951
rect 58207 45917 58216 45951
rect 58164 45908 58216 45917
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 13636 44820 13688 44872
rect 24400 44820 24452 44872
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 58164 44251 58216 44260
rect 58164 44217 58173 44251
rect 58173 44217 58207 44251
rect 58207 44217 58216 44251
rect 58164 44208 58216 44217
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 58164 43095 58216 43104
rect 58164 43061 58173 43095
rect 58173 43061 58207 43095
rect 58207 43061 58216 43095
rect 58164 43052 58216 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 16580 42551 16632 42560
rect 16580 42517 16589 42551
rect 16589 42517 16623 42551
rect 16623 42517 16632 42551
rect 16580 42508 16632 42517
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 16672 42211 16724 42220
rect 16672 42177 16681 42211
rect 16681 42177 16715 42211
rect 16715 42177 16724 42211
rect 16672 42168 16724 42177
rect 16948 42168 17000 42220
rect 16028 41964 16080 42016
rect 17316 41964 17368 42016
rect 18604 41964 18656 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 14740 41692 14792 41744
rect 18604 41735 18656 41744
rect 13912 41624 13964 41676
rect 18604 41701 18613 41735
rect 18613 41701 18647 41735
rect 18647 41701 18656 41735
rect 18604 41692 18656 41701
rect 24308 41692 24360 41744
rect 12440 41488 12492 41540
rect 12992 41531 13044 41540
rect 12992 41497 13001 41531
rect 13001 41497 13035 41531
rect 13035 41497 13044 41531
rect 12992 41488 13044 41497
rect 14556 41599 14608 41608
rect 14556 41565 14565 41599
rect 14565 41565 14599 41599
rect 14599 41565 14608 41599
rect 14556 41556 14608 41565
rect 14740 41599 14792 41608
rect 14740 41565 14749 41599
rect 14749 41565 14783 41599
rect 14783 41565 14792 41599
rect 14740 41556 14792 41565
rect 16028 41599 16080 41608
rect 16028 41565 16037 41599
rect 16037 41565 16071 41599
rect 16071 41565 16080 41599
rect 16028 41556 16080 41565
rect 16580 41556 16632 41608
rect 18696 41624 18748 41676
rect 26056 41624 26108 41676
rect 17132 41599 17184 41608
rect 17132 41565 17141 41599
rect 17141 41565 17175 41599
rect 17175 41565 17184 41599
rect 17132 41556 17184 41565
rect 17316 41599 17368 41608
rect 17316 41565 17325 41599
rect 17325 41565 17359 41599
rect 17359 41565 17368 41599
rect 17316 41556 17368 41565
rect 19984 41556 20036 41608
rect 58164 41599 58216 41608
rect 58164 41565 58173 41599
rect 58173 41565 58207 41599
rect 58207 41565 58216 41599
rect 58164 41556 58216 41565
rect 17960 41488 18012 41540
rect 20260 41488 20312 41540
rect 9864 41420 9916 41472
rect 13084 41420 13136 41472
rect 13544 41463 13596 41472
rect 13544 41429 13553 41463
rect 13553 41429 13587 41463
rect 13587 41429 13596 41463
rect 13544 41420 13596 41429
rect 14096 41463 14148 41472
rect 14096 41429 14105 41463
rect 14105 41429 14139 41463
rect 14139 41429 14148 41463
rect 14096 41420 14148 41429
rect 15292 41463 15344 41472
rect 15292 41429 15301 41463
rect 15301 41429 15335 41463
rect 15335 41429 15344 41463
rect 15292 41420 15344 41429
rect 16396 41420 16448 41472
rect 17776 41420 17828 41472
rect 19432 41420 19484 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 12992 41216 13044 41268
rect 6552 41148 6604 41200
rect 11060 41148 11112 41200
rect 16580 41216 16632 41268
rect 7656 41080 7708 41132
rect 10600 41080 10652 41132
rect 7104 41012 7156 41064
rect 13084 41123 13136 41132
rect 13084 41089 13093 41123
rect 13093 41089 13127 41123
rect 13127 41089 13136 41123
rect 16672 41191 16724 41200
rect 16672 41157 16681 41191
rect 16681 41157 16715 41191
rect 16715 41157 16724 41191
rect 16672 41148 16724 41157
rect 17132 41216 17184 41268
rect 13084 41080 13136 41089
rect 13912 41012 13964 41064
rect 13544 40944 13596 40996
rect 6368 40919 6420 40928
rect 6368 40885 6377 40919
rect 6377 40885 6411 40919
rect 6411 40885 6420 40919
rect 6368 40876 6420 40885
rect 7564 40919 7616 40928
rect 7564 40885 7573 40919
rect 7573 40885 7607 40919
rect 7607 40885 7616 40919
rect 7564 40876 7616 40885
rect 10416 40876 10468 40928
rect 12624 40919 12676 40928
rect 12624 40885 12633 40919
rect 12633 40885 12667 40919
rect 12667 40885 12676 40919
rect 12624 40876 12676 40885
rect 13728 40919 13780 40928
rect 13728 40885 13737 40919
rect 13737 40885 13771 40919
rect 13771 40885 13780 40919
rect 13728 40876 13780 40885
rect 14372 41123 14424 41132
rect 14372 41089 14381 41123
rect 14381 41089 14415 41123
rect 14415 41089 14424 41123
rect 14372 41080 14424 41089
rect 14740 41080 14792 41132
rect 15016 41123 15068 41132
rect 15016 41089 15025 41123
rect 15025 41089 15059 41123
rect 15059 41089 15068 41123
rect 15016 41080 15068 41089
rect 17040 41080 17092 41132
rect 17960 41123 18012 41132
rect 14188 40944 14240 40996
rect 17960 41089 17969 41123
rect 17969 41089 18003 41123
rect 18003 41089 18012 41123
rect 17960 41080 18012 41089
rect 18604 41080 18656 41132
rect 18696 41012 18748 41064
rect 18604 40944 18656 40996
rect 17684 40876 17736 40928
rect 18420 40919 18472 40928
rect 18420 40885 18429 40919
rect 18429 40885 18463 40919
rect 18463 40885 18472 40919
rect 18420 40876 18472 40885
rect 24124 41216 24176 41268
rect 20628 41148 20680 41200
rect 20076 41080 20128 41132
rect 20260 41080 20312 41132
rect 19524 40919 19576 40928
rect 19524 40885 19533 40919
rect 19533 40885 19567 40919
rect 19567 40885 19576 40919
rect 19524 40876 19576 40885
rect 22100 40876 22152 40928
rect 23756 40944 23808 40996
rect 23020 40876 23072 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 9864 40672 9916 40724
rect 14556 40672 14608 40724
rect 18604 40715 18656 40724
rect 18604 40681 18613 40715
rect 18613 40681 18647 40715
rect 18647 40681 18656 40715
rect 18604 40672 18656 40681
rect 15200 40604 15252 40656
rect 9220 40536 9272 40588
rect 13912 40536 13964 40588
rect 14188 40536 14240 40588
rect 14372 40579 14424 40588
rect 14372 40545 14381 40579
rect 14381 40545 14415 40579
rect 14415 40545 14424 40579
rect 14372 40536 14424 40545
rect 6092 40511 6144 40520
rect 3976 40443 4028 40452
rect 3976 40409 3985 40443
rect 3985 40409 4019 40443
rect 4019 40409 4028 40443
rect 3976 40400 4028 40409
rect 6092 40477 6101 40511
rect 6101 40477 6135 40511
rect 6135 40477 6144 40511
rect 6092 40468 6144 40477
rect 6368 40511 6420 40520
rect 6368 40477 6402 40511
rect 6402 40477 6420 40511
rect 6368 40468 6420 40477
rect 9864 40511 9916 40520
rect 9864 40477 9873 40511
rect 9873 40477 9907 40511
rect 9907 40477 9916 40511
rect 9864 40468 9916 40477
rect 10048 40511 10100 40520
rect 10048 40477 10057 40511
rect 10057 40477 10091 40511
rect 10091 40477 10100 40511
rect 10048 40468 10100 40477
rect 10508 40468 10560 40520
rect 12624 40468 12676 40520
rect 12808 40468 12860 40520
rect 13820 40468 13872 40520
rect 15384 40468 15436 40520
rect 16396 40511 16448 40520
rect 16396 40477 16430 40511
rect 16430 40477 16448 40511
rect 16396 40468 16448 40477
rect 18328 40468 18380 40520
rect 19524 40511 19576 40520
rect 19524 40477 19558 40511
rect 19558 40477 19576 40511
rect 19524 40468 19576 40477
rect 22100 40511 22152 40520
rect 22100 40477 22109 40511
rect 22109 40477 22143 40511
rect 22143 40477 22152 40511
rect 22100 40468 22152 40477
rect 10140 40400 10192 40452
rect 13084 40400 13136 40452
rect 22284 40511 22336 40520
rect 22284 40477 22293 40511
rect 22293 40477 22327 40511
rect 22327 40477 22336 40511
rect 22284 40468 22336 40477
rect 22468 40511 22520 40520
rect 22468 40477 22477 40511
rect 22477 40477 22511 40511
rect 22511 40477 22520 40511
rect 22468 40468 22520 40477
rect 23388 40468 23440 40520
rect 27344 40511 27396 40520
rect 27344 40477 27353 40511
rect 27353 40477 27387 40511
rect 27387 40477 27396 40511
rect 27344 40468 27396 40477
rect 31208 40511 31260 40520
rect 31208 40477 31217 40511
rect 31217 40477 31251 40511
rect 31251 40477 31260 40511
rect 31208 40468 31260 40477
rect 58164 40511 58216 40520
rect 58164 40477 58173 40511
rect 58173 40477 58207 40511
rect 58207 40477 58216 40511
rect 58164 40468 58216 40477
rect 4620 40332 4672 40384
rect 6368 40332 6420 40384
rect 7748 40332 7800 40384
rect 9588 40375 9640 40384
rect 9588 40341 9597 40375
rect 9597 40341 9631 40375
rect 9631 40341 9640 40375
rect 9588 40332 9640 40341
rect 12440 40332 12492 40384
rect 12624 40375 12676 40384
rect 12624 40341 12633 40375
rect 12633 40341 12667 40375
rect 12667 40341 12676 40375
rect 12624 40332 12676 40341
rect 15108 40332 15160 40384
rect 22744 40400 22796 40452
rect 23112 40400 23164 40452
rect 27620 40443 27672 40452
rect 27620 40409 27654 40443
rect 27654 40409 27672 40443
rect 27620 40400 27672 40409
rect 31484 40443 31536 40452
rect 31484 40409 31518 40443
rect 31518 40409 31536 40443
rect 31484 40400 31536 40409
rect 16948 40332 17000 40384
rect 17500 40375 17552 40384
rect 17500 40341 17509 40375
rect 17509 40341 17543 40375
rect 17543 40341 17552 40375
rect 17500 40332 17552 40341
rect 18604 40332 18656 40384
rect 19432 40332 19484 40384
rect 20352 40332 20404 40384
rect 20628 40375 20680 40384
rect 20628 40341 20637 40375
rect 20637 40341 20671 40375
rect 20671 40341 20680 40375
rect 20628 40332 20680 40341
rect 22100 40332 22152 40384
rect 23296 40332 23348 40384
rect 28724 40375 28776 40384
rect 28724 40341 28733 40375
rect 28733 40341 28767 40375
rect 28767 40341 28776 40375
rect 28724 40332 28776 40341
rect 32036 40332 32088 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 3516 40128 3568 40180
rect 3976 40171 4028 40180
rect 3976 40137 3985 40171
rect 3985 40137 4019 40171
rect 4019 40137 4028 40171
rect 3976 40128 4028 40137
rect 6092 40060 6144 40112
rect 3792 39992 3844 40044
rect 6368 39992 6420 40044
rect 2596 39967 2648 39976
rect 2596 39933 2605 39967
rect 2605 39933 2639 39967
rect 2639 39933 2648 39967
rect 2596 39924 2648 39933
rect 7748 40128 7800 40180
rect 11244 40128 11296 40180
rect 7104 40060 7156 40112
rect 9220 40060 9272 40112
rect 9588 40060 9640 40112
rect 12808 40171 12860 40180
rect 12808 40137 12817 40171
rect 12817 40137 12851 40171
rect 12851 40137 12860 40171
rect 12808 40128 12860 40137
rect 17040 40128 17092 40180
rect 19984 40128 20036 40180
rect 27620 40171 27672 40180
rect 27620 40137 27629 40171
rect 27629 40137 27663 40171
rect 27663 40137 27672 40171
rect 27620 40128 27672 40137
rect 10508 39992 10560 40044
rect 10692 39992 10744 40044
rect 11704 40035 11756 40044
rect 11704 40001 11713 40035
rect 11713 40001 11747 40035
rect 11747 40001 11756 40035
rect 11704 39992 11756 40001
rect 12624 40060 12676 40112
rect 18420 40060 18472 40112
rect 21456 40060 21508 40112
rect 28724 40060 28776 40112
rect 29092 40103 29144 40112
rect 29092 40069 29101 40103
rect 29101 40069 29135 40103
rect 29135 40069 29144 40103
rect 29092 40060 29144 40069
rect 9220 39967 9272 39976
rect 9220 39933 9229 39967
rect 9229 39933 9263 39967
rect 9263 39933 9272 39967
rect 9220 39924 9272 39933
rect 14096 39992 14148 40044
rect 17776 40035 17828 40044
rect 17776 40001 17794 40035
rect 17794 40001 17828 40035
rect 17776 39992 17828 40001
rect 20996 39992 21048 40044
rect 22284 39992 22336 40044
rect 22468 40035 22520 40044
rect 22468 40001 22477 40035
rect 22477 40001 22511 40035
rect 22511 40001 22520 40035
rect 22468 39992 22520 40001
rect 22652 40035 22704 40044
rect 22652 40001 22661 40035
rect 22661 40001 22695 40035
rect 22695 40001 22704 40035
rect 22652 39992 22704 40001
rect 22744 40035 22796 40044
rect 22744 40001 22753 40035
rect 22753 40001 22787 40035
rect 22787 40001 22796 40035
rect 22744 39992 22796 40001
rect 23020 39992 23072 40044
rect 15384 39924 15436 39976
rect 10140 39788 10192 39840
rect 10508 39788 10560 39840
rect 13820 39788 13872 39840
rect 15384 39788 15436 39840
rect 18328 39924 18380 39976
rect 27068 39992 27120 40044
rect 27988 40035 28040 40044
rect 27988 40001 27997 40035
rect 27997 40001 28031 40035
rect 28031 40001 28040 40035
rect 27988 39992 28040 40001
rect 28264 40035 28316 40044
rect 28264 40001 28273 40035
rect 28273 40001 28307 40035
rect 28307 40001 28316 40035
rect 28264 39992 28316 40001
rect 23572 39831 23624 39840
rect 23572 39797 23581 39831
rect 23581 39797 23615 39831
rect 23615 39797 23624 39831
rect 23572 39788 23624 39797
rect 24768 39788 24820 39840
rect 27068 39831 27120 39840
rect 27068 39797 27077 39831
rect 27077 39797 27111 39831
rect 27111 39797 27120 39831
rect 27068 39788 27120 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 3792 39627 3844 39636
rect 3792 39593 3801 39627
rect 3801 39593 3835 39627
rect 3835 39593 3844 39627
rect 3792 39584 3844 39593
rect 2596 39448 2648 39500
rect 5264 39516 5316 39568
rect 4620 39448 4672 39500
rect 11704 39584 11756 39636
rect 14096 39584 14148 39636
rect 15016 39584 15068 39636
rect 15200 39584 15252 39636
rect 16304 39584 16356 39636
rect 23020 39584 23072 39636
rect 23480 39584 23532 39636
rect 31484 39627 31536 39636
rect 31484 39593 31493 39627
rect 31493 39593 31527 39627
rect 31527 39593 31536 39627
rect 31484 39584 31536 39593
rect 15384 39448 15436 39500
rect 4896 39380 4948 39432
rect 7288 39380 7340 39432
rect 7656 39423 7708 39432
rect 7656 39389 7665 39423
rect 7665 39389 7699 39423
rect 7699 39389 7708 39423
rect 7656 39380 7708 39389
rect 9220 39423 9272 39432
rect 9220 39389 9229 39423
rect 9229 39389 9263 39423
rect 9263 39389 9272 39423
rect 9220 39380 9272 39389
rect 11060 39423 11112 39432
rect 11060 39389 11069 39423
rect 11069 39389 11103 39423
rect 11103 39389 11112 39423
rect 11060 39380 11112 39389
rect 11244 39423 11296 39432
rect 11244 39389 11253 39423
rect 11253 39389 11287 39423
rect 11287 39389 11296 39423
rect 11244 39380 11296 39389
rect 4620 39312 4672 39364
rect 6092 39312 6144 39364
rect 9956 39312 10008 39364
rect 14188 39380 14240 39432
rect 22560 39380 22612 39432
rect 23204 39423 23256 39432
rect 23204 39389 23213 39423
rect 23213 39389 23247 39423
rect 23247 39389 23256 39423
rect 23204 39380 23256 39389
rect 6828 39244 6880 39296
rect 8208 39244 8260 39296
rect 13728 39312 13780 39364
rect 22008 39312 22060 39364
rect 22100 39355 22152 39364
rect 22100 39321 22118 39355
rect 22118 39321 22152 39355
rect 22100 39312 22152 39321
rect 22468 39312 22520 39364
rect 22744 39312 22796 39364
rect 23848 39380 23900 39432
rect 27344 39380 27396 39432
rect 28264 39380 28316 39432
rect 30288 39380 30340 39432
rect 31116 39423 31168 39432
rect 31116 39389 31125 39423
rect 31125 39389 31159 39423
rect 31159 39389 31168 39423
rect 31116 39380 31168 39389
rect 31300 39380 31352 39432
rect 24768 39312 24820 39364
rect 27528 39355 27580 39364
rect 27528 39321 27562 39355
rect 27562 39321 27580 39355
rect 27528 39312 27580 39321
rect 31760 39312 31812 39364
rect 32036 39312 32088 39364
rect 10600 39287 10652 39296
rect 10600 39253 10609 39287
rect 10609 39253 10643 39287
rect 10643 39253 10652 39287
rect 10600 39244 10652 39253
rect 16856 39287 16908 39296
rect 16856 39253 16865 39287
rect 16865 39253 16899 39287
rect 16899 39253 16908 39287
rect 16856 39244 16908 39253
rect 20996 39287 21048 39296
rect 20996 39253 21005 39287
rect 21005 39253 21039 39287
rect 21039 39253 21048 39287
rect 20996 39244 21048 39253
rect 23388 39244 23440 39296
rect 28632 39287 28684 39296
rect 28632 39253 28641 39287
rect 28641 39253 28675 39287
rect 28675 39253 28684 39287
rect 28632 39244 28684 39253
rect 30564 39244 30616 39296
rect 31300 39244 31352 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 9956 39083 10008 39092
rect 2504 38904 2556 38956
rect 9956 39049 9965 39083
rect 9965 39049 9999 39083
rect 9999 39049 10008 39083
rect 9956 39040 10008 39049
rect 13084 39083 13136 39092
rect 5080 38972 5132 39024
rect 4620 38947 4672 38956
rect 4620 38913 4629 38947
rect 4629 38913 4663 38947
rect 4663 38913 4672 38947
rect 4620 38904 4672 38913
rect 4896 38947 4948 38956
rect 4896 38913 4905 38947
rect 4905 38913 4939 38947
rect 4939 38913 4948 38947
rect 6368 38947 6420 38956
rect 4896 38904 4948 38913
rect 6368 38913 6377 38947
rect 6377 38913 6411 38947
rect 6411 38913 6420 38947
rect 6368 38904 6420 38913
rect 6828 38904 6880 38956
rect 13084 39049 13093 39083
rect 13093 39049 13127 39083
rect 13127 39049 13136 39083
rect 13084 39040 13136 39049
rect 18328 39083 18380 39092
rect 18328 39049 18337 39083
rect 18337 39049 18371 39083
rect 18371 39049 18380 39083
rect 18328 39040 18380 39049
rect 22652 39040 22704 39092
rect 27528 39083 27580 39092
rect 27528 39049 27537 39083
rect 27537 39049 27571 39083
rect 27571 39049 27580 39083
rect 27528 39040 27580 39049
rect 27988 39040 28040 39092
rect 4712 38768 4764 38820
rect 8208 38836 8260 38888
rect 10692 38904 10744 38956
rect 12900 38947 12952 38956
rect 12900 38913 12909 38947
rect 12909 38913 12943 38947
rect 12943 38913 12952 38947
rect 12900 38904 12952 38913
rect 16856 38904 16908 38956
rect 21456 38972 21508 39024
rect 23112 38972 23164 39024
rect 23572 38904 23624 38956
rect 26976 38947 27028 38956
rect 26976 38913 26985 38947
rect 26985 38913 27019 38947
rect 27019 38913 27028 38947
rect 31116 38972 31168 39024
rect 26976 38904 27028 38913
rect 28264 38904 28316 38956
rect 10140 38768 10192 38820
rect 10416 38768 10468 38820
rect 3976 38700 4028 38752
rect 4620 38700 4672 38752
rect 6552 38700 6604 38752
rect 6644 38700 6696 38752
rect 7288 38700 7340 38752
rect 13820 38700 13872 38752
rect 27068 38836 27120 38888
rect 28080 38836 28132 38888
rect 58164 38811 58216 38820
rect 58164 38777 58173 38811
rect 58173 38777 58207 38811
rect 58207 38777 58216 38811
rect 58164 38768 58216 38777
rect 18972 38700 19024 38752
rect 23848 38743 23900 38752
rect 23848 38709 23857 38743
rect 23857 38709 23891 38743
rect 23891 38709 23900 38743
rect 23848 38700 23900 38709
rect 26792 38700 26844 38752
rect 28816 38700 28868 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 4712 38496 4764 38548
rect 6092 38539 6144 38548
rect 6092 38505 6101 38539
rect 6101 38505 6135 38539
rect 6135 38505 6144 38539
rect 6092 38496 6144 38505
rect 2872 38335 2924 38344
rect 2872 38301 2881 38335
rect 2881 38301 2915 38335
rect 2915 38301 2924 38335
rect 2872 38292 2924 38301
rect 4620 38360 4672 38412
rect 3056 38335 3108 38344
rect 3056 38301 3065 38335
rect 3065 38301 3099 38335
rect 3099 38301 3108 38335
rect 3056 38292 3108 38301
rect 4896 38292 4948 38344
rect 6460 38428 6512 38480
rect 6644 38360 6696 38412
rect 3976 38267 4028 38276
rect 2136 38156 2188 38208
rect 3424 38156 3476 38208
rect 3976 38233 3985 38267
rect 3985 38233 4019 38267
rect 4019 38233 4028 38267
rect 3976 38224 4028 38233
rect 6736 38335 6788 38344
rect 6736 38301 6745 38335
rect 6745 38301 6779 38335
rect 6779 38301 6788 38335
rect 6736 38292 6788 38301
rect 7656 38292 7708 38344
rect 10600 38292 10652 38344
rect 17500 38496 17552 38548
rect 23480 38496 23532 38548
rect 25504 38496 25556 38548
rect 28080 38539 28132 38548
rect 28080 38505 28089 38539
rect 28089 38505 28123 38539
rect 28123 38505 28132 38539
rect 28080 38496 28132 38505
rect 16120 38335 16172 38344
rect 16120 38301 16129 38335
rect 16129 38301 16163 38335
rect 16163 38301 16172 38335
rect 16764 38335 16816 38344
rect 16120 38292 16172 38301
rect 16764 38301 16773 38335
rect 16773 38301 16807 38335
rect 16807 38301 16816 38335
rect 16764 38292 16816 38301
rect 17040 38335 17092 38344
rect 17040 38301 17049 38335
rect 17049 38301 17083 38335
rect 17083 38301 17092 38335
rect 17040 38292 17092 38301
rect 17132 38335 17184 38344
rect 17132 38301 17141 38335
rect 17141 38301 17175 38335
rect 17175 38301 17184 38335
rect 31208 38360 31260 38412
rect 31668 38360 31720 38412
rect 17132 38292 17184 38301
rect 19432 38335 19484 38344
rect 19432 38301 19442 38335
rect 19442 38301 19476 38335
rect 19476 38301 19484 38335
rect 19432 38292 19484 38301
rect 20260 38292 20312 38344
rect 24676 38292 24728 38344
rect 28632 38292 28684 38344
rect 30196 38292 30248 38344
rect 6644 38224 6696 38276
rect 9312 38267 9364 38276
rect 9312 38233 9321 38267
rect 9321 38233 9355 38267
rect 9355 38233 9364 38267
rect 9312 38224 9364 38233
rect 15936 38267 15988 38276
rect 15936 38233 15945 38267
rect 15945 38233 15979 38267
rect 15979 38233 15988 38267
rect 15936 38224 15988 38233
rect 6368 38156 6420 38208
rect 6460 38156 6512 38208
rect 8024 38156 8076 38208
rect 9220 38156 9272 38208
rect 10232 38156 10284 38208
rect 19248 38224 19300 38276
rect 20628 38224 20680 38276
rect 24400 38224 24452 38276
rect 29092 38224 29144 38276
rect 30380 38224 30432 38276
rect 31944 38292 31996 38344
rect 31760 38267 31812 38276
rect 31760 38233 31769 38267
rect 31769 38233 31803 38267
rect 31803 38233 31812 38267
rect 31760 38224 31812 38233
rect 17316 38199 17368 38208
rect 17316 38165 17325 38199
rect 17325 38165 17359 38199
rect 17359 38165 17368 38199
rect 17316 38156 17368 38165
rect 21088 38156 21140 38208
rect 25964 38199 26016 38208
rect 25964 38165 25973 38199
rect 25973 38165 26007 38199
rect 26007 38165 26016 38199
rect 25964 38156 26016 38165
rect 29552 38199 29604 38208
rect 29552 38165 29561 38199
rect 29561 38165 29595 38199
rect 29595 38165 29604 38199
rect 29552 38156 29604 38165
rect 30472 38156 30524 38208
rect 32312 38199 32364 38208
rect 32312 38165 32321 38199
rect 32321 38165 32355 38199
rect 32355 38165 32364 38199
rect 32312 38156 32364 38165
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 3056 37995 3108 38004
rect 3056 37961 3065 37995
rect 3065 37961 3099 37995
rect 3099 37961 3108 37995
rect 3056 37952 3108 37961
rect 6368 37952 6420 38004
rect 10048 37952 10100 38004
rect 3424 37927 3476 37936
rect 3424 37893 3433 37927
rect 3433 37893 3467 37927
rect 3467 37893 3476 37927
rect 3424 37884 3476 37893
rect 10416 37927 10468 37936
rect 10416 37893 10425 37927
rect 10425 37893 10459 37927
rect 10459 37893 10468 37927
rect 10416 37884 10468 37893
rect 11060 37884 11112 37936
rect 12532 37952 12584 38004
rect 15936 37952 15988 38004
rect 12440 37884 12492 37936
rect 19248 37952 19300 38004
rect 19616 37952 19668 38004
rect 24400 37995 24452 38004
rect 24400 37961 24409 37995
rect 24409 37961 24443 37995
rect 24443 37961 24452 37995
rect 24400 37952 24452 37961
rect 19984 37884 20036 37936
rect 23480 37884 23532 37936
rect 3240 37859 3292 37868
rect 3240 37825 3249 37859
rect 3249 37825 3283 37859
rect 3283 37825 3292 37859
rect 3240 37816 3292 37825
rect 11244 37816 11296 37868
rect 11888 37859 11940 37868
rect 11888 37825 11897 37859
rect 11897 37825 11931 37859
rect 11931 37825 11940 37859
rect 11888 37816 11940 37825
rect 16120 37816 16172 37868
rect 17132 37816 17184 37868
rect 17316 37859 17368 37868
rect 17316 37825 17325 37859
rect 17325 37825 17359 37859
rect 17359 37825 17368 37859
rect 17316 37816 17368 37825
rect 17408 37859 17460 37868
rect 17408 37825 17418 37859
rect 17418 37825 17452 37859
rect 17452 37825 17460 37859
rect 17408 37816 17460 37825
rect 12900 37748 12952 37800
rect 17868 37680 17920 37732
rect 2872 37612 2924 37664
rect 5632 37612 5684 37664
rect 8300 37612 8352 37664
rect 9312 37612 9364 37664
rect 17960 37655 18012 37664
rect 17960 37621 17969 37655
rect 17969 37621 18003 37655
rect 18003 37621 18012 37655
rect 17960 37612 18012 37621
rect 18328 37816 18380 37868
rect 18512 37816 18564 37868
rect 20076 37816 20128 37868
rect 20444 37859 20496 37868
rect 20444 37825 20453 37859
rect 20453 37825 20487 37859
rect 20487 37825 20496 37859
rect 20444 37816 20496 37825
rect 24124 37816 24176 37868
rect 20260 37680 20312 37732
rect 24676 37680 24728 37732
rect 24952 37816 25004 37868
rect 19432 37612 19484 37664
rect 19984 37612 20036 37664
rect 23020 37612 23072 37664
rect 24124 37612 24176 37664
rect 24584 37612 24636 37664
rect 25964 37884 26016 37936
rect 28816 37816 28868 37868
rect 30288 37859 30340 37868
rect 30288 37825 30297 37859
rect 30297 37825 30331 37859
rect 30331 37825 30340 37859
rect 30288 37816 30340 37825
rect 30472 37859 30524 37868
rect 30472 37825 30481 37859
rect 30481 37825 30515 37859
rect 30515 37825 30524 37859
rect 30472 37816 30524 37825
rect 30656 37859 30708 37868
rect 30656 37825 30665 37859
rect 30665 37825 30699 37859
rect 30699 37825 30708 37859
rect 30656 37816 30708 37825
rect 32588 37859 32640 37868
rect 32588 37825 32622 37859
rect 32622 37825 32640 37859
rect 32588 37816 32640 37825
rect 31116 37748 31168 37800
rect 31668 37748 31720 37800
rect 27436 37612 27488 37664
rect 28908 37612 28960 37664
rect 30932 37655 30984 37664
rect 30932 37621 30941 37655
rect 30941 37621 30975 37655
rect 30975 37621 30984 37655
rect 30932 37612 30984 37621
rect 33784 37612 33836 37664
rect 35532 37612 35584 37664
rect 58164 37655 58216 37664
rect 58164 37621 58173 37655
rect 58173 37621 58207 37655
rect 58207 37621 58216 37655
rect 58164 37612 58216 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 16764 37451 16816 37460
rect 16764 37417 16773 37451
rect 16773 37417 16807 37451
rect 16807 37417 16816 37451
rect 16764 37408 16816 37417
rect 17408 37408 17460 37460
rect 18512 37408 18564 37460
rect 20444 37451 20496 37460
rect 20444 37417 20453 37451
rect 20453 37417 20487 37451
rect 20487 37417 20496 37451
rect 20444 37408 20496 37417
rect 17868 37340 17920 37392
rect 2596 37204 2648 37256
rect 2136 37179 2188 37188
rect 2136 37145 2170 37179
rect 2170 37145 2188 37179
rect 2136 37136 2188 37145
rect 7012 37136 7064 37188
rect 3240 37111 3292 37120
rect 3240 37077 3249 37111
rect 3249 37077 3283 37111
rect 3283 37077 3292 37111
rect 3240 37068 3292 37077
rect 7472 37247 7524 37256
rect 7472 37213 7481 37247
rect 7481 37213 7515 37247
rect 7515 37213 7524 37247
rect 7748 37247 7800 37256
rect 7472 37204 7524 37213
rect 7748 37213 7757 37247
rect 7757 37213 7791 37247
rect 7791 37213 7800 37247
rect 7748 37204 7800 37213
rect 7840 37247 7892 37256
rect 7840 37213 7849 37247
rect 7849 37213 7883 37247
rect 7883 37213 7892 37247
rect 7840 37204 7892 37213
rect 11888 37204 11940 37256
rect 13176 37204 13228 37256
rect 15384 37247 15436 37256
rect 15384 37213 15393 37247
rect 15393 37213 15427 37247
rect 15427 37213 15436 37247
rect 15384 37204 15436 37213
rect 17040 37204 17092 37256
rect 17592 37247 17644 37256
rect 17592 37213 17607 37247
rect 17607 37213 17641 37247
rect 17641 37213 17644 37247
rect 17776 37247 17828 37256
rect 17592 37204 17644 37213
rect 17776 37213 17785 37247
rect 17785 37213 17819 37247
rect 17819 37213 17828 37247
rect 17776 37204 17828 37213
rect 18972 37272 19024 37324
rect 23020 37340 23072 37392
rect 31668 37340 31720 37392
rect 34888 37340 34940 37392
rect 7656 37179 7708 37188
rect 7656 37145 7665 37179
rect 7665 37145 7699 37179
rect 7699 37145 7708 37179
rect 7656 37136 7708 37145
rect 10232 37136 10284 37188
rect 14648 37136 14700 37188
rect 8392 37068 8444 37120
rect 14556 37068 14608 37120
rect 15476 37136 15528 37188
rect 17316 37136 17368 37188
rect 20260 37204 20312 37256
rect 22008 37204 22060 37256
rect 19616 37179 19668 37188
rect 19616 37145 19625 37179
rect 19625 37145 19659 37179
rect 19659 37145 19668 37179
rect 19616 37136 19668 37145
rect 20444 37136 20496 37188
rect 20536 37136 20588 37188
rect 23388 37247 23440 37256
rect 23388 37213 23397 37247
rect 23397 37213 23431 37247
rect 23431 37213 23440 37247
rect 23388 37204 23440 37213
rect 24768 37204 24820 37256
rect 31668 37204 31720 37256
rect 32312 37204 32364 37256
rect 33508 37204 33560 37256
rect 20628 37068 20680 37120
rect 22284 37111 22336 37120
rect 22284 37077 22293 37111
rect 22293 37077 22327 37111
rect 22327 37077 22336 37111
rect 22284 37068 22336 37077
rect 22928 37068 22980 37120
rect 23020 37068 23072 37120
rect 24584 37136 24636 37188
rect 25044 37136 25096 37188
rect 30932 37136 30984 37188
rect 34152 37136 34204 37188
rect 24492 37068 24544 37120
rect 28172 37068 28224 37120
rect 29276 37068 29328 37120
rect 29644 37111 29696 37120
rect 29644 37077 29653 37111
rect 29653 37077 29687 37111
rect 29687 37077 29696 37111
rect 29644 37068 29696 37077
rect 31944 37111 31996 37120
rect 31944 37077 31953 37111
rect 31953 37077 31987 37111
rect 31987 37077 31996 37111
rect 31944 37068 31996 37077
rect 33876 37068 33928 37120
rect 35624 37204 35676 37256
rect 35348 37111 35400 37120
rect 35348 37077 35357 37111
rect 35357 37077 35391 37111
rect 35391 37077 35400 37111
rect 35348 37068 35400 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 2596 36796 2648 36848
rect 5172 36796 5224 36848
rect 7656 36864 7708 36916
rect 12532 36864 12584 36916
rect 14648 36864 14700 36916
rect 15476 36907 15528 36916
rect 15476 36873 15485 36907
rect 15485 36873 15519 36907
rect 15519 36873 15528 36907
rect 15476 36864 15528 36873
rect 17776 36864 17828 36916
rect 18972 36864 19024 36916
rect 20536 36864 20588 36916
rect 24768 36864 24820 36916
rect 30380 36864 30432 36916
rect 32588 36907 32640 36916
rect 32588 36873 32597 36907
rect 32597 36873 32631 36907
rect 32631 36873 32640 36907
rect 32588 36864 32640 36873
rect 6828 36839 6880 36848
rect 6828 36805 6837 36839
rect 6837 36805 6871 36839
rect 6871 36805 6880 36839
rect 6828 36796 6880 36805
rect 7472 36796 7524 36848
rect 7840 36728 7892 36780
rect 7932 36771 7984 36780
rect 7932 36737 7941 36771
rect 7941 36737 7975 36771
rect 7975 36737 7984 36771
rect 7932 36728 7984 36737
rect 9772 36728 9824 36780
rect 14004 36728 14056 36780
rect 16764 36796 16816 36848
rect 19432 36796 19484 36848
rect 15384 36728 15436 36780
rect 15732 36771 15784 36780
rect 15732 36737 15741 36771
rect 15741 36737 15775 36771
rect 15775 36737 15784 36771
rect 15732 36728 15784 36737
rect 16120 36771 16172 36780
rect 16120 36737 16129 36771
rect 16129 36737 16163 36771
rect 16163 36737 16172 36771
rect 17040 36771 17092 36780
rect 16120 36728 16172 36737
rect 17040 36737 17049 36771
rect 17049 36737 17083 36771
rect 17083 36737 17092 36771
rect 17040 36728 17092 36737
rect 17868 36728 17920 36780
rect 19800 36771 19852 36780
rect 19800 36737 19809 36771
rect 19809 36737 19843 36771
rect 19843 36737 19852 36771
rect 19984 36771 20036 36780
rect 19800 36728 19852 36737
rect 19984 36737 19993 36771
rect 19993 36737 20027 36771
rect 20027 36737 20036 36771
rect 19984 36728 20036 36737
rect 28816 36796 28868 36848
rect 33416 36864 33468 36916
rect 35440 36864 35492 36916
rect 8300 36592 8352 36644
rect 15844 36592 15896 36644
rect 18696 36660 18748 36712
rect 19248 36660 19300 36712
rect 19984 36592 20036 36644
rect 20260 36592 20312 36644
rect 22284 36728 22336 36780
rect 23020 36771 23072 36780
rect 23020 36737 23029 36771
rect 23029 36737 23063 36771
rect 23063 36737 23072 36771
rect 23020 36728 23072 36737
rect 23572 36728 23624 36780
rect 27436 36771 27488 36780
rect 27436 36737 27445 36771
rect 27445 36737 27479 36771
rect 27479 36737 27488 36771
rect 27436 36728 27488 36737
rect 27528 36728 27580 36780
rect 27988 36728 28040 36780
rect 29276 36771 29328 36780
rect 29276 36737 29285 36771
rect 29285 36737 29319 36771
rect 29319 36737 29328 36771
rect 29276 36728 29328 36737
rect 29460 36771 29512 36780
rect 29460 36737 29469 36771
rect 29469 36737 29503 36771
rect 29503 36737 29512 36771
rect 29460 36728 29512 36737
rect 24492 36660 24544 36712
rect 29000 36660 29052 36712
rect 29644 36771 29696 36780
rect 29644 36737 29653 36771
rect 29653 36737 29687 36771
rect 29687 36737 29696 36771
rect 29644 36728 29696 36737
rect 30288 36728 30340 36780
rect 33876 36796 33928 36848
rect 31392 36703 31444 36712
rect 31392 36669 31401 36703
rect 31401 36669 31435 36703
rect 31435 36669 31444 36703
rect 31392 36660 31444 36669
rect 33140 36728 33192 36780
rect 33508 36728 33560 36780
rect 34244 36728 34296 36780
rect 34888 36771 34940 36780
rect 34888 36737 34897 36771
rect 34897 36737 34931 36771
rect 34931 36737 34940 36771
rect 34888 36728 34940 36737
rect 34704 36660 34756 36712
rect 25228 36592 25280 36644
rect 7104 36567 7156 36576
rect 7104 36533 7113 36567
rect 7113 36533 7147 36567
rect 7147 36533 7156 36567
rect 7104 36524 7156 36533
rect 7472 36524 7524 36576
rect 15476 36524 15528 36576
rect 16120 36524 16172 36576
rect 17592 36524 17644 36576
rect 19432 36524 19484 36576
rect 19800 36524 19852 36576
rect 20352 36524 20404 36576
rect 22284 36524 22336 36576
rect 22652 36567 22704 36576
rect 22652 36533 22661 36567
rect 22661 36533 22695 36567
rect 22695 36533 22704 36567
rect 22652 36524 22704 36533
rect 28448 36524 28500 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 5172 36363 5224 36372
rect 5172 36329 5181 36363
rect 5181 36329 5215 36363
rect 5215 36329 5224 36363
rect 5172 36320 5224 36329
rect 7012 36363 7064 36372
rect 7012 36329 7021 36363
rect 7021 36329 7055 36363
rect 7055 36329 7064 36363
rect 7012 36320 7064 36329
rect 11060 36320 11112 36372
rect 12532 36363 12584 36372
rect 12532 36329 12541 36363
rect 12541 36329 12575 36363
rect 12575 36329 12584 36363
rect 12532 36320 12584 36329
rect 14004 36320 14056 36372
rect 14372 36320 14424 36372
rect 15108 36320 15160 36372
rect 15752 36320 15804 36372
rect 16304 36363 16356 36372
rect 16304 36329 16313 36363
rect 16313 36329 16347 36363
rect 16347 36329 16356 36363
rect 16304 36320 16356 36329
rect 27068 36363 27120 36372
rect 27068 36329 27077 36363
rect 27077 36329 27111 36363
rect 27111 36329 27120 36363
rect 27068 36320 27120 36329
rect 27528 36363 27580 36372
rect 27528 36329 27537 36363
rect 27537 36329 27571 36363
rect 27571 36329 27580 36363
rect 27528 36320 27580 36329
rect 29460 36320 29512 36372
rect 34152 36363 34204 36372
rect 34152 36329 34161 36363
rect 34161 36329 34195 36363
rect 34195 36329 34204 36363
rect 34152 36320 34204 36329
rect 34704 36320 34756 36372
rect 23664 36252 23716 36304
rect 28816 36252 28868 36304
rect 32312 36252 32364 36304
rect 2596 36184 2648 36236
rect 5356 36184 5408 36236
rect 20996 36184 21048 36236
rect 4620 36048 4672 36100
rect 6644 35980 6696 36032
rect 7472 36159 7524 36168
rect 7472 36125 7481 36159
rect 7481 36125 7515 36159
rect 7515 36125 7524 36159
rect 7472 36116 7524 36125
rect 9312 36116 9364 36168
rect 10232 36116 10284 36168
rect 14372 36159 14424 36168
rect 14372 36125 14381 36159
rect 14381 36125 14415 36159
rect 14415 36125 14424 36159
rect 14372 36116 14424 36125
rect 10416 36091 10468 36100
rect 10416 36057 10450 36091
rect 10450 36057 10468 36091
rect 10416 36048 10468 36057
rect 13084 36048 13136 36100
rect 13360 36091 13412 36100
rect 13360 36057 13369 36091
rect 13369 36057 13403 36091
rect 13403 36057 13412 36091
rect 13360 36048 13412 36057
rect 13820 36048 13872 36100
rect 14280 36048 14332 36100
rect 14556 36159 14608 36168
rect 14556 36125 14565 36159
rect 14565 36125 14599 36159
rect 14599 36125 14608 36159
rect 14556 36116 14608 36125
rect 14740 36159 14792 36168
rect 14740 36125 14749 36159
rect 14749 36125 14783 36159
rect 14783 36125 14792 36159
rect 22284 36159 22336 36168
rect 14740 36116 14792 36125
rect 22284 36125 22293 36159
rect 22293 36125 22327 36159
rect 22327 36125 22336 36159
rect 22284 36116 22336 36125
rect 27436 36184 27488 36236
rect 23480 36159 23532 36168
rect 23480 36125 23489 36159
rect 23489 36125 23523 36159
rect 23523 36125 23532 36159
rect 23480 36116 23532 36125
rect 24492 36116 24544 36168
rect 27068 36116 27120 36168
rect 34796 36184 34848 36236
rect 28172 36159 28224 36168
rect 15844 36048 15896 36100
rect 17316 36048 17368 36100
rect 9496 35980 9548 36032
rect 10140 35980 10192 36032
rect 11704 35980 11756 36032
rect 14004 35980 14056 36032
rect 22100 36023 22152 36032
rect 22100 35989 22109 36023
rect 22109 35989 22143 36023
rect 22143 35989 22152 36023
rect 23020 36048 23072 36100
rect 23848 36091 23900 36100
rect 23848 36057 23857 36091
rect 23857 36057 23891 36091
rect 23891 36057 23900 36091
rect 23848 36048 23900 36057
rect 26240 36091 26292 36100
rect 26240 36057 26258 36091
rect 26258 36057 26292 36091
rect 26240 36048 26292 36057
rect 22100 35980 22152 35989
rect 23664 35980 23716 36032
rect 24400 36023 24452 36032
rect 24400 35989 24409 36023
rect 24409 35989 24443 36023
rect 24443 35989 24452 36023
rect 24400 35980 24452 35989
rect 28172 36125 28181 36159
rect 28181 36125 28215 36159
rect 28215 36125 28224 36159
rect 28172 36116 28224 36125
rect 28448 36048 28500 36100
rect 29460 36048 29512 36100
rect 31392 36116 31444 36168
rect 33508 36116 33560 36168
rect 30472 36048 30524 36100
rect 29000 35980 29052 36032
rect 30380 36023 30432 36032
rect 30380 35989 30389 36023
rect 30389 35989 30423 36023
rect 30423 35989 30432 36023
rect 33692 36048 33744 36100
rect 35348 36116 35400 36168
rect 58164 36159 58216 36168
rect 58164 36125 58173 36159
rect 58173 36125 58207 36159
rect 58207 36125 58216 36159
rect 58164 36116 58216 36125
rect 30380 35980 30432 35989
rect 33416 35980 33468 36032
rect 35440 36048 35492 36100
rect 34704 35980 34756 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 13360 35776 13412 35828
rect 24676 35776 24728 35828
rect 5172 35708 5224 35760
rect 2872 35640 2924 35692
rect 7196 35640 7248 35692
rect 11060 35708 11112 35760
rect 11520 35751 11572 35760
rect 11520 35717 11529 35751
rect 11529 35717 11563 35751
rect 11563 35717 11572 35751
rect 11520 35708 11572 35717
rect 13176 35751 13228 35760
rect 13176 35717 13185 35751
rect 13185 35717 13219 35751
rect 13219 35717 13228 35751
rect 13176 35708 13228 35717
rect 23480 35751 23532 35760
rect 23480 35717 23489 35751
rect 23489 35717 23523 35751
rect 23523 35717 23532 35751
rect 23480 35708 23532 35717
rect 26240 35776 26292 35828
rect 28264 35776 28316 35828
rect 30656 35776 30708 35828
rect 33140 35776 33192 35828
rect 10232 35640 10284 35692
rect 11980 35640 12032 35692
rect 13452 35640 13504 35692
rect 16488 35640 16540 35692
rect 17040 35640 17092 35692
rect 18512 35640 18564 35692
rect 23664 35683 23716 35692
rect 23664 35649 23673 35683
rect 23673 35649 23707 35683
rect 23707 35649 23716 35683
rect 23664 35640 23716 35649
rect 24400 35640 24452 35692
rect 7932 35572 7984 35624
rect 9312 35615 9364 35624
rect 9312 35581 9321 35615
rect 9321 35581 9355 35615
rect 9355 35581 9364 35615
rect 9312 35572 9364 35581
rect 9772 35615 9824 35624
rect 9772 35581 9781 35615
rect 9781 35581 9815 35615
rect 9815 35581 9824 35615
rect 9772 35572 9824 35581
rect 10140 35572 10192 35624
rect 10692 35572 10744 35624
rect 25228 35640 25280 35692
rect 27988 35708 28040 35760
rect 33784 35708 33836 35760
rect 31760 35640 31812 35692
rect 33692 35683 33744 35692
rect 33692 35649 33701 35683
rect 33701 35649 33735 35683
rect 33735 35649 33744 35683
rect 33692 35640 33744 35649
rect 14004 35504 14056 35556
rect 28172 35504 28224 35556
rect 4712 35479 4764 35488
rect 4712 35445 4721 35479
rect 4721 35445 4755 35479
rect 4755 35445 4764 35479
rect 4712 35436 4764 35445
rect 6092 35436 6144 35488
rect 6552 35436 6604 35488
rect 10600 35436 10652 35488
rect 13912 35479 13964 35488
rect 13912 35445 13921 35479
rect 13921 35445 13955 35479
rect 13955 35445 13964 35479
rect 13912 35436 13964 35445
rect 14740 35436 14792 35488
rect 17776 35479 17828 35488
rect 17776 35445 17785 35479
rect 17785 35445 17819 35479
rect 17819 35445 17828 35479
rect 17776 35436 17828 35445
rect 22376 35479 22428 35488
rect 22376 35445 22385 35479
rect 22385 35445 22419 35479
rect 22419 35445 22428 35479
rect 22376 35436 22428 35445
rect 23020 35479 23072 35488
rect 23020 35445 23029 35479
rect 23029 35445 23063 35479
rect 23063 35445 23072 35479
rect 23020 35436 23072 35445
rect 25872 35436 25924 35488
rect 34244 35504 34296 35556
rect 36452 35504 36504 35556
rect 33692 35436 33744 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 4620 35232 4672 35284
rect 6092 35232 6144 35284
rect 7196 35275 7248 35284
rect 7196 35241 7205 35275
rect 7205 35241 7239 35275
rect 7239 35241 7248 35275
rect 7196 35232 7248 35241
rect 2688 34960 2740 35012
rect 4712 35071 4764 35080
rect 4712 35037 4721 35071
rect 4721 35037 4755 35071
rect 4755 35037 4764 35071
rect 4988 35164 5040 35216
rect 7564 35164 7616 35216
rect 11980 35275 12032 35284
rect 4712 35028 4764 35037
rect 11980 35241 11989 35275
rect 11989 35241 12023 35275
rect 12023 35241 12032 35275
rect 11980 35232 12032 35241
rect 19156 35232 19208 35284
rect 19432 35275 19484 35284
rect 19432 35241 19441 35275
rect 19441 35241 19475 35275
rect 19475 35241 19484 35275
rect 19432 35232 19484 35241
rect 25044 35275 25096 35284
rect 25044 35241 25053 35275
rect 25053 35241 25087 35275
rect 25087 35241 25096 35275
rect 25044 35232 25096 35241
rect 10048 35096 10100 35148
rect 10232 35096 10284 35148
rect 15384 35096 15436 35148
rect 18604 35096 18656 35148
rect 5356 34960 5408 35012
rect 6368 35003 6420 35012
rect 6368 34969 6377 35003
rect 6377 34969 6411 35003
rect 6411 34969 6420 35003
rect 6368 34960 6420 34969
rect 6552 35003 6604 35012
rect 6552 34969 6561 35003
rect 6561 34969 6595 35003
rect 6595 34969 6604 35003
rect 6552 34960 6604 34969
rect 6736 34960 6788 35012
rect 9956 35028 10008 35080
rect 11980 35028 12032 35080
rect 13452 35028 13504 35080
rect 17684 35028 17736 35080
rect 20536 35028 20588 35080
rect 22008 35096 22060 35148
rect 23848 35096 23900 35148
rect 22744 35028 22796 35080
rect 24400 35071 24452 35080
rect 11060 34960 11112 35012
rect 13176 35003 13228 35012
rect 13176 34969 13185 35003
rect 13185 34969 13219 35003
rect 13219 34969 13228 35003
rect 13176 34960 13228 34969
rect 14096 34960 14148 35012
rect 17132 34960 17184 35012
rect 20352 34960 20404 35012
rect 24400 35037 24409 35071
rect 24409 35037 24443 35071
rect 24443 35037 24452 35071
rect 24400 35028 24452 35037
rect 24676 35071 24728 35080
rect 24676 35037 24685 35071
rect 24685 35037 24719 35071
rect 24719 35037 24728 35071
rect 24676 35028 24728 35037
rect 5632 34892 5684 34944
rect 15108 34892 15160 34944
rect 18512 34935 18564 34944
rect 18512 34901 18521 34935
rect 18521 34901 18555 34935
rect 18555 34901 18564 34935
rect 18512 34892 18564 34901
rect 20260 34935 20312 34944
rect 20260 34901 20269 34935
rect 20269 34901 20303 34935
rect 20303 34901 20312 34935
rect 20260 34892 20312 34901
rect 22192 34892 22244 34944
rect 22560 34892 22612 34944
rect 23940 34892 23992 34944
rect 24308 34892 24360 34944
rect 25964 35164 26016 35216
rect 33324 35164 33376 35216
rect 29276 35028 29328 35080
rect 30196 35028 30248 35080
rect 31760 35071 31812 35080
rect 31760 35037 31769 35071
rect 31769 35037 31803 35071
rect 31803 35037 31812 35071
rect 58164 35071 58216 35080
rect 31760 35028 31812 35037
rect 58164 35037 58173 35071
rect 58173 35037 58207 35071
rect 58207 35037 58216 35071
rect 58164 35028 58216 35037
rect 28908 34960 28960 35012
rect 29828 34960 29880 35012
rect 29552 34892 29604 34944
rect 30472 35003 30524 35012
rect 30472 34969 30481 35003
rect 30481 34969 30515 35003
rect 30515 34969 30524 35003
rect 30472 34960 30524 34969
rect 31208 34960 31260 35012
rect 31576 34892 31628 34944
rect 34244 34892 34296 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 4620 34688 4672 34740
rect 5632 34688 5684 34740
rect 9128 34688 9180 34740
rect 10416 34688 10468 34740
rect 2596 34595 2648 34604
rect 2596 34561 2605 34595
rect 2605 34561 2639 34595
rect 2639 34561 2648 34595
rect 2596 34552 2648 34561
rect 4712 34416 4764 34468
rect 6552 34620 6604 34672
rect 9496 34663 9548 34672
rect 9496 34629 9505 34663
rect 9505 34629 9539 34663
rect 9539 34629 9548 34663
rect 9496 34620 9548 34629
rect 5448 34552 5500 34604
rect 7564 34552 7616 34604
rect 8392 34595 8444 34604
rect 8392 34561 8401 34595
rect 8401 34561 8435 34595
rect 8435 34561 8444 34595
rect 8392 34552 8444 34561
rect 8668 34595 8720 34604
rect 8024 34484 8076 34536
rect 8668 34561 8677 34595
rect 8677 34561 8711 34595
rect 8711 34561 8720 34595
rect 8668 34552 8720 34561
rect 9588 34552 9640 34604
rect 9956 34552 10008 34604
rect 12808 34620 12860 34672
rect 16120 34688 16172 34740
rect 17132 34731 17184 34740
rect 17132 34697 17141 34731
rect 17141 34697 17175 34731
rect 17175 34697 17184 34731
rect 17132 34688 17184 34697
rect 17592 34688 17644 34740
rect 16304 34620 16356 34672
rect 17316 34620 17368 34672
rect 10968 34595 11020 34604
rect 10048 34484 10100 34536
rect 10968 34561 10977 34595
rect 10977 34561 11011 34595
rect 11011 34561 11020 34595
rect 10968 34552 11020 34561
rect 11520 34595 11572 34604
rect 11520 34561 11529 34595
rect 11529 34561 11563 34595
rect 11563 34561 11572 34595
rect 11520 34552 11572 34561
rect 11704 34595 11756 34604
rect 11704 34561 11713 34595
rect 11713 34561 11747 34595
rect 11747 34561 11756 34595
rect 11704 34552 11756 34561
rect 13268 34595 13320 34604
rect 13268 34561 13277 34595
rect 13277 34561 13311 34595
rect 13311 34561 13320 34595
rect 13268 34552 13320 34561
rect 13452 34595 13504 34604
rect 13452 34561 13461 34595
rect 13461 34561 13495 34595
rect 13495 34561 13504 34595
rect 13452 34552 13504 34561
rect 13176 34484 13228 34536
rect 11520 34416 11572 34468
rect 16764 34552 16816 34604
rect 17684 34552 17736 34604
rect 17868 34552 17920 34604
rect 18696 34552 18748 34604
rect 20076 34688 20128 34740
rect 20352 34688 20404 34740
rect 20536 34620 20588 34672
rect 25872 34688 25924 34740
rect 21824 34620 21876 34672
rect 19432 34552 19484 34604
rect 18052 34484 18104 34536
rect 16304 34416 16356 34468
rect 17500 34416 17552 34468
rect 18604 34416 18656 34468
rect 19248 34416 19300 34468
rect 20260 34552 20312 34604
rect 20628 34552 20680 34604
rect 21732 34552 21784 34604
rect 22192 34595 22244 34604
rect 22192 34561 22201 34595
rect 22201 34561 22235 34595
rect 22235 34561 22244 34595
rect 22192 34552 22244 34561
rect 28356 34620 28408 34672
rect 30564 34688 30616 34740
rect 31576 34731 31628 34740
rect 31576 34697 31585 34731
rect 31585 34697 31619 34731
rect 31619 34697 31628 34731
rect 31576 34688 31628 34697
rect 33968 34688 34020 34740
rect 21548 34484 21600 34536
rect 22100 34484 22152 34536
rect 22744 34552 22796 34604
rect 28264 34484 28316 34536
rect 22468 34416 22520 34468
rect 29000 34416 29052 34468
rect 29552 34595 29604 34604
rect 29552 34561 29561 34595
rect 29561 34561 29595 34595
rect 29595 34561 29604 34595
rect 29552 34552 29604 34561
rect 29736 34595 29788 34604
rect 29736 34561 29745 34595
rect 29745 34561 29779 34595
rect 29779 34561 29788 34595
rect 29736 34552 29788 34561
rect 33508 34552 33560 34604
rect 29828 34484 29880 34536
rect 34244 34552 34296 34604
rect 35808 34484 35860 34536
rect 34796 34416 34848 34468
rect 4896 34348 4948 34400
rect 5448 34348 5500 34400
rect 7564 34348 7616 34400
rect 11796 34348 11848 34400
rect 14556 34348 14608 34400
rect 19800 34348 19852 34400
rect 22836 34391 22888 34400
rect 22836 34357 22845 34391
rect 22845 34357 22879 34391
rect 22879 34357 22888 34391
rect 22836 34348 22888 34357
rect 24768 34391 24820 34400
rect 24768 34357 24777 34391
rect 24777 34357 24811 34391
rect 24811 34357 24820 34391
rect 24768 34348 24820 34357
rect 27712 34391 27764 34400
rect 27712 34357 27721 34391
rect 27721 34357 27755 34391
rect 27755 34357 27764 34391
rect 27712 34348 27764 34357
rect 30196 34348 30248 34400
rect 33324 34391 33376 34400
rect 33324 34357 33333 34391
rect 33333 34357 33367 34391
rect 33367 34357 33376 34391
rect 33324 34348 33376 34357
rect 33876 34348 33928 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 5448 34144 5500 34196
rect 11060 34187 11112 34196
rect 11060 34153 11069 34187
rect 11069 34153 11103 34187
rect 11103 34153 11112 34187
rect 11060 34144 11112 34153
rect 14556 34187 14608 34196
rect 14556 34153 14565 34187
rect 14565 34153 14599 34187
rect 14599 34153 14608 34187
rect 14556 34144 14608 34153
rect 15108 34144 15160 34196
rect 5080 34076 5132 34128
rect 14280 34076 14332 34128
rect 17316 34076 17368 34128
rect 4896 34008 4948 34060
rect 6736 34008 6788 34060
rect 10048 34008 10100 34060
rect 5448 33940 5500 33992
rect 10140 33940 10192 33992
rect 10600 33983 10652 33992
rect 10600 33949 10622 33983
rect 10622 33949 10652 33983
rect 10600 33940 10652 33949
rect 11520 33983 11572 33992
rect 11520 33949 11529 33983
rect 11529 33949 11563 33983
rect 11563 33949 11572 33983
rect 11520 33940 11572 33949
rect 5080 33915 5132 33924
rect 5080 33881 5089 33915
rect 5089 33881 5123 33915
rect 5123 33881 5132 33915
rect 5080 33872 5132 33881
rect 5540 33872 5592 33924
rect 6368 33872 6420 33924
rect 3792 33847 3844 33856
rect 3792 33813 3801 33847
rect 3801 33813 3835 33847
rect 3835 33813 3844 33847
rect 3792 33804 3844 33813
rect 7380 33804 7432 33856
rect 8116 33804 8168 33856
rect 8392 33804 8444 33856
rect 14924 33940 14976 33992
rect 17040 33940 17092 33992
rect 14648 33915 14700 33924
rect 14648 33881 14657 33915
rect 14657 33881 14691 33915
rect 14691 33881 14700 33915
rect 14648 33872 14700 33881
rect 17500 33940 17552 33992
rect 17868 34008 17920 34060
rect 17776 33983 17828 33992
rect 17776 33949 17785 33983
rect 17785 33949 17819 33983
rect 17819 33949 17828 33983
rect 17776 33940 17828 33949
rect 18604 34144 18656 34196
rect 21824 34187 21876 34196
rect 21824 34153 21833 34187
rect 21833 34153 21867 34187
rect 21867 34153 21876 34187
rect 21824 34144 21876 34153
rect 25872 34187 25924 34196
rect 25872 34153 25881 34187
rect 25881 34153 25915 34187
rect 25915 34153 25924 34187
rect 25872 34144 25924 34153
rect 34796 34144 34848 34196
rect 18512 34008 18564 34060
rect 17868 33872 17920 33924
rect 20444 34008 20496 34060
rect 22008 34008 22060 34060
rect 29736 34008 29788 34060
rect 30748 34008 30800 34060
rect 19800 33983 19852 33992
rect 19800 33949 19814 33983
rect 19814 33949 19848 33983
rect 19848 33949 19852 33983
rect 19800 33940 19852 33949
rect 22836 33940 22888 33992
rect 23480 33940 23532 33992
rect 27068 33940 27120 33992
rect 29920 33983 29972 33992
rect 29920 33949 29929 33983
rect 29929 33949 29963 33983
rect 29963 33949 29972 33983
rect 29920 33940 29972 33949
rect 30380 33940 30432 33992
rect 33692 34076 33744 34128
rect 33508 33983 33560 33992
rect 33508 33949 33517 33983
rect 33517 33949 33551 33983
rect 33551 33949 33560 33983
rect 33508 33940 33560 33949
rect 33968 34008 34020 34060
rect 33876 33983 33928 33992
rect 33876 33949 33885 33983
rect 33885 33949 33919 33983
rect 33919 33949 33928 33983
rect 33876 33940 33928 33949
rect 15936 33804 15988 33856
rect 16948 33804 17000 33856
rect 20260 33872 20312 33924
rect 21456 33915 21508 33924
rect 21456 33881 21465 33915
rect 21465 33881 21499 33915
rect 21499 33881 21508 33915
rect 21456 33872 21508 33881
rect 25044 33915 25096 33924
rect 19984 33847 20036 33856
rect 19984 33813 19993 33847
rect 19993 33813 20027 33847
rect 20027 33813 20036 33847
rect 19984 33804 20036 33813
rect 25044 33881 25053 33915
rect 25053 33881 25087 33915
rect 25087 33881 25096 33915
rect 25044 33872 25096 33881
rect 27252 33915 27304 33924
rect 27252 33881 27286 33915
rect 27286 33881 27304 33915
rect 31208 33915 31260 33924
rect 27252 33872 27304 33881
rect 31208 33881 31217 33915
rect 31217 33881 31251 33915
rect 31251 33881 31260 33915
rect 31208 33872 31260 33881
rect 31392 33915 31444 33924
rect 31392 33881 31401 33915
rect 31401 33881 31435 33915
rect 31435 33881 31444 33915
rect 31392 33872 31444 33881
rect 34428 33872 34480 33924
rect 34612 33940 34664 33992
rect 24492 33804 24544 33856
rect 25228 33847 25280 33856
rect 25228 33813 25237 33847
rect 25237 33813 25271 33847
rect 25271 33813 25280 33847
rect 25228 33804 25280 33813
rect 28356 33847 28408 33856
rect 28356 33813 28365 33847
rect 28365 33813 28399 33847
rect 28399 33813 28408 33847
rect 28356 33804 28408 33813
rect 30564 33804 30616 33856
rect 34152 33847 34204 33856
rect 34152 33813 34161 33847
rect 34161 33813 34195 33847
rect 34195 33813 34204 33847
rect 34152 33804 34204 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 4712 33600 4764 33652
rect 5172 33600 5224 33652
rect 6460 33600 6512 33652
rect 7104 33600 7156 33652
rect 8024 33643 8076 33652
rect 8024 33609 8033 33643
rect 8033 33609 8067 33643
rect 8067 33609 8076 33643
rect 8024 33600 8076 33609
rect 8116 33600 8168 33652
rect 3792 33532 3844 33584
rect 4620 33575 4672 33584
rect 4620 33541 4629 33575
rect 4629 33541 4663 33575
rect 4663 33541 4672 33575
rect 4620 33532 4672 33541
rect 5356 33532 5408 33584
rect 17776 33600 17828 33652
rect 27252 33643 27304 33652
rect 27252 33609 27261 33643
rect 27261 33609 27295 33643
rect 27295 33609 27304 33643
rect 27252 33600 27304 33609
rect 13912 33532 13964 33584
rect 14924 33532 14976 33584
rect 2596 33507 2648 33516
rect 2596 33473 2605 33507
rect 2605 33473 2639 33507
rect 2639 33473 2648 33507
rect 2596 33464 2648 33473
rect 5540 33464 5592 33516
rect 6920 33507 6972 33516
rect 6920 33473 6954 33507
rect 6954 33473 6972 33507
rect 6920 33464 6972 33473
rect 11704 33464 11756 33516
rect 15016 33464 15068 33516
rect 15936 33532 15988 33584
rect 16304 33532 16356 33584
rect 19156 33575 19208 33584
rect 19156 33541 19165 33575
rect 19165 33541 19199 33575
rect 19199 33541 19208 33575
rect 19156 33532 19208 33541
rect 15292 33507 15344 33516
rect 15292 33473 15301 33507
rect 15301 33473 15335 33507
rect 15335 33473 15344 33507
rect 15292 33464 15344 33473
rect 15476 33507 15528 33516
rect 15476 33473 15485 33507
rect 15485 33473 15519 33507
rect 15519 33473 15528 33507
rect 15476 33464 15528 33473
rect 16488 33464 16540 33516
rect 5080 33260 5132 33312
rect 17040 33396 17092 33448
rect 8668 33328 8720 33380
rect 18328 33371 18380 33380
rect 7012 33260 7064 33312
rect 10968 33260 11020 33312
rect 12992 33303 13044 33312
rect 12992 33269 13001 33303
rect 13001 33269 13035 33303
rect 13035 33269 13044 33303
rect 12992 33260 13044 33269
rect 18328 33337 18337 33371
rect 18337 33337 18371 33371
rect 18371 33337 18380 33371
rect 18328 33328 18380 33337
rect 16948 33260 17000 33312
rect 21916 33464 21968 33516
rect 24676 33532 24728 33584
rect 24400 33507 24452 33516
rect 24400 33473 24409 33507
rect 24409 33473 24443 33507
rect 24443 33473 24452 33507
rect 24400 33464 24452 33473
rect 24952 33464 25004 33516
rect 25228 33507 25280 33516
rect 25228 33473 25237 33507
rect 25237 33473 25271 33507
rect 25271 33473 25280 33507
rect 25228 33464 25280 33473
rect 25872 33464 25924 33516
rect 24768 33396 24820 33448
rect 23848 33328 23900 33380
rect 24308 33328 24360 33380
rect 26884 33328 26936 33380
rect 23664 33260 23716 33312
rect 26240 33260 26292 33312
rect 26976 33260 27028 33312
rect 27712 33507 27764 33516
rect 27712 33473 27721 33507
rect 27721 33473 27755 33507
rect 27755 33473 27764 33507
rect 27712 33464 27764 33473
rect 28172 33464 28224 33516
rect 29552 33464 29604 33516
rect 30656 33600 30708 33652
rect 34428 33600 34480 33652
rect 32312 33532 32364 33584
rect 34152 33532 34204 33584
rect 30288 33396 30340 33448
rect 30564 33507 30616 33516
rect 30564 33473 30573 33507
rect 30573 33473 30607 33507
rect 30607 33473 30616 33507
rect 30564 33464 30616 33473
rect 30748 33507 30800 33516
rect 30748 33473 30757 33507
rect 30757 33473 30791 33507
rect 30791 33473 30800 33507
rect 30748 33464 30800 33473
rect 31668 33464 31720 33516
rect 32956 33507 33008 33516
rect 32956 33473 32990 33507
rect 32990 33473 33008 33507
rect 32956 33464 33008 33473
rect 36084 33396 36136 33448
rect 31116 33328 31168 33380
rect 58164 33371 58216 33380
rect 58164 33337 58173 33371
rect 58173 33337 58207 33371
rect 58207 33337 58216 33371
rect 58164 33328 58216 33337
rect 29552 33303 29604 33312
rect 29552 33269 29561 33303
rect 29561 33269 29595 33303
rect 29595 33269 29604 33303
rect 29552 33260 29604 33269
rect 30104 33303 30156 33312
rect 30104 33269 30113 33303
rect 30113 33269 30147 33303
rect 30147 33269 30156 33303
rect 30104 33260 30156 33269
rect 34152 33260 34204 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 5264 33056 5316 33108
rect 6920 33056 6972 33108
rect 15292 33056 15344 33108
rect 17960 33056 18012 33108
rect 20352 33056 20404 33108
rect 24400 33056 24452 33108
rect 26240 33056 26292 33108
rect 28172 33056 28224 33108
rect 4988 32988 5040 33040
rect 17224 32988 17276 33040
rect 5724 32716 5776 32768
rect 6644 32852 6696 32904
rect 9864 32920 9916 32972
rect 16488 32920 16540 32972
rect 24308 32920 24360 32972
rect 24952 32920 25004 32972
rect 32312 32963 32364 32972
rect 32312 32929 32321 32963
rect 32321 32929 32355 32963
rect 32355 32929 32364 32963
rect 32312 32920 32364 32929
rect 33968 32920 34020 32972
rect 7380 32895 7432 32904
rect 7380 32861 7389 32895
rect 7389 32861 7423 32895
rect 7423 32861 7432 32895
rect 7380 32852 7432 32861
rect 8024 32895 8076 32904
rect 8024 32861 8033 32895
rect 8033 32861 8067 32895
rect 8067 32861 8076 32895
rect 8024 32852 8076 32861
rect 9312 32852 9364 32904
rect 11060 32852 11112 32904
rect 7564 32784 7616 32836
rect 7748 32784 7800 32836
rect 9772 32784 9824 32836
rect 10140 32827 10192 32836
rect 10140 32793 10149 32827
rect 10149 32793 10183 32827
rect 10183 32793 10192 32827
rect 10140 32784 10192 32793
rect 10692 32784 10744 32836
rect 16120 32852 16172 32904
rect 16304 32895 16356 32904
rect 16304 32861 16314 32895
rect 16314 32861 16348 32895
rect 16348 32861 16356 32895
rect 16304 32852 16356 32861
rect 16948 32852 17000 32904
rect 17684 32895 17736 32904
rect 17684 32861 17693 32895
rect 17693 32861 17727 32895
rect 17727 32861 17736 32895
rect 17684 32852 17736 32861
rect 17776 32852 17828 32904
rect 23480 32895 23532 32904
rect 23480 32861 23489 32895
rect 23489 32861 23523 32895
rect 23523 32861 23532 32895
rect 23480 32852 23532 32861
rect 26884 32895 26936 32904
rect 26884 32861 26902 32895
rect 26902 32861 26936 32895
rect 26884 32852 26936 32861
rect 27068 32852 27120 32904
rect 27252 32852 27304 32904
rect 12992 32784 13044 32836
rect 13544 32784 13596 32836
rect 16028 32784 16080 32836
rect 18420 32827 18472 32836
rect 18420 32793 18429 32827
rect 18429 32793 18463 32827
rect 18463 32793 18472 32827
rect 18420 32784 18472 32793
rect 18696 32784 18748 32836
rect 19984 32784 20036 32836
rect 21364 32784 21416 32836
rect 23664 32827 23716 32836
rect 23664 32793 23673 32827
rect 23673 32793 23707 32827
rect 23707 32793 23716 32827
rect 23664 32784 23716 32793
rect 24216 32784 24268 32836
rect 29920 32852 29972 32904
rect 31760 32852 31812 32904
rect 32128 32852 32180 32904
rect 35808 32895 35860 32904
rect 35808 32861 35826 32895
rect 35826 32861 35860 32895
rect 36084 32895 36136 32904
rect 35808 32852 35860 32861
rect 36084 32861 36093 32895
rect 36093 32861 36127 32895
rect 36127 32861 36136 32895
rect 36084 32852 36136 32861
rect 38936 32852 38988 32904
rect 34152 32784 34204 32836
rect 10784 32716 10836 32768
rect 10968 32716 11020 32768
rect 15016 32716 15068 32768
rect 16120 32716 16172 32768
rect 17592 32716 17644 32768
rect 22100 32759 22152 32768
rect 22100 32725 22109 32759
rect 22109 32725 22143 32759
rect 22143 32725 22152 32759
rect 22100 32716 22152 32725
rect 25044 32716 25096 32768
rect 29736 32759 29788 32768
rect 29736 32725 29745 32759
rect 29745 32725 29779 32759
rect 29779 32725 29788 32759
rect 29736 32716 29788 32725
rect 30380 32716 30432 32768
rect 32404 32716 32456 32768
rect 34612 32716 34664 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 5448 32512 5500 32564
rect 5540 32512 5592 32564
rect 12808 32512 12860 32564
rect 14004 32555 14056 32564
rect 14004 32521 14013 32555
rect 14013 32521 14047 32555
rect 14047 32521 14056 32555
rect 14004 32512 14056 32521
rect 14740 32512 14792 32564
rect 17684 32512 17736 32564
rect 17960 32512 18012 32564
rect 18420 32512 18472 32564
rect 24308 32512 24360 32564
rect 9404 32444 9456 32496
rect 9956 32444 10008 32496
rect 2136 32376 2188 32428
rect 1860 32308 1912 32360
rect 7104 32376 7156 32428
rect 7748 32376 7800 32428
rect 6552 32308 6604 32360
rect 8576 32351 8628 32360
rect 8576 32317 8585 32351
rect 8585 32317 8619 32351
rect 8619 32317 8628 32351
rect 8576 32308 8628 32317
rect 10416 32308 10468 32360
rect 10784 32419 10836 32428
rect 10784 32385 10793 32419
rect 10793 32385 10827 32419
rect 10827 32385 10836 32419
rect 10784 32376 10836 32385
rect 10968 32419 11020 32428
rect 10968 32385 10977 32419
rect 10977 32385 11011 32419
rect 11011 32385 11020 32419
rect 10968 32376 11020 32385
rect 14924 32376 14976 32428
rect 15016 32376 15068 32428
rect 17776 32419 17828 32428
rect 17776 32385 17785 32419
rect 17785 32385 17819 32419
rect 17819 32385 17828 32419
rect 17776 32376 17828 32385
rect 15384 32308 15436 32360
rect 17684 32308 17736 32360
rect 17960 32419 18012 32428
rect 17960 32385 17969 32419
rect 17969 32385 18003 32419
rect 18003 32385 18012 32419
rect 20536 32444 20588 32496
rect 29552 32512 29604 32564
rect 31208 32512 31260 32564
rect 32956 32512 33008 32564
rect 28448 32487 28500 32496
rect 28448 32453 28457 32487
rect 28457 32453 28491 32487
rect 28491 32453 28500 32487
rect 28448 32444 28500 32453
rect 32312 32444 32364 32496
rect 17960 32376 18012 32385
rect 18328 32376 18380 32428
rect 22100 32376 22152 32428
rect 24032 32376 24084 32428
rect 24308 32419 24360 32428
rect 24308 32385 24317 32419
rect 24317 32385 24351 32419
rect 24351 32385 24360 32419
rect 24308 32376 24360 32385
rect 28540 32419 28592 32428
rect 3608 32215 3660 32224
rect 3608 32181 3617 32215
rect 3617 32181 3651 32215
rect 3651 32181 3660 32215
rect 3608 32172 3660 32181
rect 6828 32172 6880 32224
rect 10324 32215 10376 32224
rect 10324 32181 10333 32215
rect 10333 32181 10367 32215
rect 10367 32181 10376 32215
rect 10324 32172 10376 32181
rect 10416 32172 10468 32224
rect 10692 32172 10744 32224
rect 10968 32172 11020 32224
rect 17960 32240 18012 32292
rect 13820 32172 13872 32224
rect 17868 32172 17920 32224
rect 28172 32308 28224 32360
rect 28540 32385 28549 32419
rect 28549 32385 28583 32419
rect 28583 32385 28592 32419
rect 28540 32376 28592 32385
rect 28724 32419 28776 32428
rect 28724 32385 28733 32419
rect 28733 32385 28767 32419
rect 28767 32385 28776 32419
rect 28724 32376 28776 32385
rect 30840 32376 30892 32428
rect 32404 32419 32456 32428
rect 29368 32308 29420 32360
rect 32404 32385 32413 32419
rect 32413 32385 32447 32419
rect 32447 32385 32456 32419
rect 32404 32376 32456 32385
rect 32588 32419 32640 32428
rect 32588 32385 32597 32419
rect 32597 32385 32631 32419
rect 32631 32385 32640 32419
rect 32588 32376 32640 32385
rect 36636 32376 36688 32428
rect 33508 32308 33560 32360
rect 38936 32308 38988 32360
rect 23480 32240 23532 32292
rect 28724 32240 28776 32292
rect 29644 32240 29696 32292
rect 23756 32172 23808 32224
rect 24400 32172 24452 32224
rect 26700 32172 26752 32224
rect 37280 32215 37332 32224
rect 37280 32181 37289 32215
rect 37289 32181 37323 32215
rect 37323 32181 37332 32215
rect 37280 32172 37332 32181
rect 58164 32215 58216 32224
rect 58164 32181 58173 32215
rect 58173 32181 58207 32215
rect 58207 32181 58216 32215
rect 58164 32172 58216 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2136 32011 2188 32020
rect 2136 31977 2145 32011
rect 2145 31977 2179 32011
rect 2179 31977 2188 32011
rect 2136 31968 2188 31977
rect 6184 31968 6236 32020
rect 7012 31968 7064 32020
rect 8208 31968 8260 32020
rect 11060 31968 11112 32020
rect 14556 31968 14608 32020
rect 23756 31968 23808 32020
rect 24124 31968 24176 32020
rect 27252 31968 27304 32020
rect 5264 31900 5316 31952
rect 5448 31900 5500 31952
rect 2320 31764 2372 31816
rect 2596 31807 2648 31816
rect 2596 31773 2605 31807
rect 2605 31773 2639 31807
rect 2639 31773 2648 31807
rect 2596 31764 2648 31773
rect 2780 31807 2832 31816
rect 2780 31773 2789 31807
rect 2789 31773 2823 31807
rect 2823 31773 2832 31807
rect 2780 31764 2832 31773
rect 4988 31764 5040 31816
rect 2688 31696 2740 31748
rect 4896 31696 4948 31748
rect 5264 31807 5316 31816
rect 5264 31773 5273 31807
rect 5273 31773 5307 31807
rect 5307 31773 5316 31807
rect 5264 31764 5316 31773
rect 8300 31900 8352 31952
rect 11336 31900 11388 31952
rect 17224 31900 17276 31952
rect 27896 31900 27948 31952
rect 8208 31832 8260 31884
rect 12900 31832 12952 31884
rect 10324 31764 10376 31816
rect 13452 31832 13504 31884
rect 17960 31832 18012 31884
rect 4804 31671 4856 31680
rect 4804 31637 4813 31671
rect 4813 31637 4847 31671
rect 4847 31637 4856 31671
rect 4804 31628 4856 31637
rect 7380 31696 7432 31748
rect 13084 31696 13136 31748
rect 14556 31804 14608 31816
rect 14556 31770 14565 31804
rect 14565 31770 14599 31804
rect 14599 31770 14608 31804
rect 14740 31807 14792 31816
rect 14556 31764 14608 31770
rect 14740 31773 14749 31807
rect 14749 31773 14783 31807
rect 14783 31773 14792 31807
rect 14740 31764 14792 31773
rect 16856 31764 16908 31816
rect 20444 31764 20496 31816
rect 24676 31832 24728 31884
rect 28448 31968 28500 32020
rect 30748 31968 30800 32020
rect 31024 31968 31076 32020
rect 31392 31968 31444 32020
rect 32588 31968 32640 32020
rect 36636 32011 36688 32020
rect 36636 31977 36645 32011
rect 36645 31977 36679 32011
rect 36679 31977 36688 32011
rect 36636 31968 36688 31977
rect 33416 31900 33468 31952
rect 22560 31807 22612 31816
rect 22560 31773 22569 31807
rect 22569 31773 22603 31807
rect 22603 31773 22612 31807
rect 22560 31764 22612 31773
rect 24860 31764 24912 31816
rect 28172 31764 28224 31816
rect 28356 31807 28408 31816
rect 28356 31773 28365 31807
rect 28365 31773 28399 31807
rect 28399 31773 28408 31807
rect 28632 31807 28684 31816
rect 28356 31764 28408 31773
rect 28632 31773 28641 31807
rect 28641 31773 28675 31807
rect 28675 31773 28684 31807
rect 28632 31764 28684 31773
rect 30104 31764 30156 31816
rect 30932 31764 30984 31816
rect 35992 31807 36044 31816
rect 35992 31773 36001 31807
rect 36001 31773 36035 31807
rect 36035 31773 36044 31807
rect 35992 31764 36044 31773
rect 36176 31807 36228 31816
rect 36176 31773 36185 31807
rect 36185 31773 36219 31807
rect 36219 31773 36228 31807
rect 36176 31764 36228 31773
rect 6552 31628 6604 31680
rect 14096 31671 14148 31680
rect 14096 31637 14105 31671
rect 14105 31637 14139 31671
rect 14139 31637 14148 31671
rect 14096 31628 14148 31637
rect 15568 31696 15620 31748
rect 28448 31739 28500 31748
rect 28448 31705 28457 31739
rect 28457 31705 28491 31739
rect 28491 31705 28500 31739
rect 28448 31696 28500 31705
rect 15844 31628 15896 31680
rect 17868 31628 17920 31680
rect 26056 31671 26108 31680
rect 26056 31637 26065 31671
rect 26065 31637 26099 31671
rect 26099 31637 26108 31671
rect 26056 31628 26108 31637
rect 32404 31628 32456 31680
rect 36268 31628 36320 31680
rect 37648 31628 37700 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 2596 31424 2648 31476
rect 5264 31424 5316 31476
rect 8300 31467 8352 31476
rect 8300 31433 8309 31467
rect 8309 31433 8343 31467
rect 8343 31433 8352 31467
rect 8300 31424 8352 31433
rect 13084 31424 13136 31476
rect 13544 31424 13596 31476
rect 5540 31356 5592 31408
rect 6552 31356 6604 31408
rect 14096 31356 14148 31408
rect 2872 31288 2924 31340
rect 3332 31288 3384 31340
rect 5632 31331 5684 31340
rect 5632 31297 5641 31331
rect 5641 31297 5675 31331
rect 5675 31297 5684 31331
rect 5632 31288 5684 31297
rect 3608 31220 3660 31272
rect 6828 31331 6880 31340
rect 6828 31297 6842 31331
rect 6842 31297 6876 31331
rect 6876 31297 6880 31331
rect 6828 31288 6880 31297
rect 7380 31288 7432 31340
rect 10140 31288 10192 31340
rect 14924 31331 14976 31340
rect 14924 31297 14933 31331
rect 14933 31297 14967 31331
rect 14967 31297 14976 31331
rect 14924 31288 14976 31297
rect 15384 31424 15436 31476
rect 16028 31424 16080 31476
rect 16856 31424 16908 31476
rect 25320 31424 25372 31476
rect 25964 31424 26016 31476
rect 32128 31467 32180 31476
rect 32128 31433 32137 31467
rect 32137 31433 32171 31467
rect 32171 31433 32180 31467
rect 36176 31467 36228 31476
rect 32128 31424 32180 31433
rect 15476 31356 15528 31408
rect 7932 31220 7984 31272
rect 15200 31220 15252 31272
rect 16948 31288 17000 31340
rect 13912 31152 13964 31204
rect 14648 31152 14700 31204
rect 16580 31220 16632 31272
rect 16672 31220 16724 31272
rect 28540 31356 28592 31408
rect 31576 31356 31628 31408
rect 36176 31433 36185 31467
rect 36185 31433 36219 31467
rect 36219 31433 36228 31467
rect 36176 31424 36228 31433
rect 18696 31288 18748 31340
rect 19984 31288 20036 31340
rect 20996 31288 21048 31340
rect 21456 31288 21508 31340
rect 23388 31288 23440 31340
rect 23848 31288 23900 31340
rect 24032 31288 24084 31340
rect 17868 31220 17920 31272
rect 25504 31288 25556 31340
rect 26056 31288 26108 31340
rect 28080 31288 28132 31340
rect 30932 31288 30984 31340
rect 31208 31331 31260 31340
rect 31208 31297 31217 31331
rect 31217 31297 31251 31331
rect 31251 31297 31260 31331
rect 31208 31288 31260 31297
rect 31944 31288 31996 31340
rect 28540 31220 28592 31272
rect 30748 31220 30800 31272
rect 32404 31331 32456 31340
rect 32404 31297 32413 31331
rect 32413 31297 32447 31331
rect 32447 31297 32456 31331
rect 32404 31288 32456 31297
rect 33232 31288 33284 31340
rect 35808 31331 35860 31340
rect 35808 31297 35817 31331
rect 35817 31297 35851 31331
rect 35851 31297 35860 31331
rect 35808 31288 35860 31297
rect 33508 31220 33560 31272
rect 37280 31288 37332 31340
rect 37648 31331 37700 31340
rect 37648 31297 37657 31331
rect 37657 31297 37691 31331
rect 37691 31297 37700 31331
rect 37648 31288 37700 31297
rect 2320 31084 2372 31136
rect 4068 31084 4120 31136
rect 6644 31084 6696 31136
rect 10140 31127 10192 31136
rect 10140 31093 10149 31127
rect 10149 31093 10183 31127
rect 10183 31093 10192 31127
rect 10140 31084 10192 31093
rect 12348 31084 12400 31136
rect 16028 31084 16080 31136
rect 20720 31084 20772 31136
rect 22744 31084 22796 31136
rect 24032 31127 24084 31136
rect 24032 31093 24041 31127
rect 24041 31093 24075 31127
rect 24075 31093 24084 31127
rect 24032 31084 24084 31093
rect 28080 31127 28132 31136
rect 28080 31093 28089 31127
rect 28089 31093 28123 31127
rect 28123 31093 28132 31127
rect 28080 31084 28132 31093
rect 28908 31084 28960 31136
rect 30564 31084 30616 31136
rect 32220 31084 32272 31136
rect 38936 31127 38988 31136
rect 38936 31093 38945 31127
rect 38945 31093 38979 31127
rect 38979 31093 38988 31127
rect 38936 31084 38988 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 7932 30880 7984 30932
rect 12348 30880 12400 30932
rect 14924 30880 14976 30932
rect 1860 30787 1912 30796
rect 1860 30753 1869 30787
rect 1869 30753 1903 30787
rect 1903 30753 1912 30787
rect 1860 30744 1912 30753
rect 8208 30676 8260 30728
rect 11060 30676 11112 30728
rect 13084 30719 13136 30728
rect 13084 30685 13093 30719
rect 13093 30685 13127 30719
rect 13127 30685 13136 30719
rect 13084 30676 13136 30685
rect 13176 30719 13228 30728
rect 13176 30685 13185 30719
rect 13185 30685 13219 30719
rect 13219 30685 13228 30719
rect 13176 30676 13228 30685
rect 13820 30676 13872 30728
rect 14280 30719 14332 30728
rect 14280 30685 14289 30719
rect 14289 30685 14323 30719
rect 14323 30685 14332 30719
rect 14280 30676 14332 30685
rect 15476 30880 15528 30932
rect 16764 30880 16816 30932
rect 20076 30812 20128 30864
rect 15200 30676 15252 30728
rect 15752 30676 15804 30728
rect 17868 30676 17920 30728
rect 22560 30812 22612 30864
rect 22468 30744 22520 30796
rect 2136 30651 2188 30660
rect 2136 30617 2170 30651
rect 2170 30617 2188 30651
rect 4804 30651 4856 30660
rect 2136 30608 2188 30617
rect 4804 30617 4838 30651
rect 4838 30617 4856 30651
rect 4804 30608 4856 30617
rect 6644 30651 6696 30660
rect 6644 30617 6678 30651
rect 6678 30617 6696 30651
rect 6644 30608 6696 30617
rect 13268 30608 13320 30660
rect 15660 30608 15712 30660
rect 18052 30608 18104 30660
rect 22744 30719 22796 30728
rect 22744 30685 22753 30719
rect 22753 30685 22787 30719
rect 22787 30685 22796 30719
rect 27252 30744 27304 30796
rect 32312 30812 32364 30864
rect 34060 30812 34112 30864
rect 30288 30744 30340 30796
rect 22744 30676 22796 30685
rect 24308 30676 24360 30728
rect 24584 30676 24636 30728
rect 30104 30719 30156 30728
rect 30104 30685 30113 30719
rect 30113 30685 30147 30719
rect 30147 30685 30156 30719
rect 30104 30676 30156 30685
rect 30196 30676 30248 30728
rect 30472 30676 30524 30728
rect 32220 30719 32272 30728
rect 32220 30685 32229 30719
rect 32229 30685 32263 30719
rect 32263 30685 32272 30719
rect 32220 30676 32272 30685
rect 33324 30744 33376 30796
rect 36268 30812 36320 30864
rect 33416 30719 33468 30728
rect 33416 30685 33425 30719
rect 33425 30685 33459 30719
rect 33459 30685 33468 30719
rect 33416 30676 33468 30685
rect 33508 30719 33560 30728
rect 33508 30685 33517 30719
rect 33517 30685 33551 30719
rect 33551 30685 33560 30719
rect 33784 30719 33836 30728
rect 33508 30676 33560 30685
rect 33784 30685 33793 30719
rect 33793 30685 33827 30719
rect 33827 30685 33836 30719
rect 33784 30676 33836 30685
rect 35348 30719 35400 30728
rect 35348 30685 35357 30719
rect 35357 30685 35391 30719
rect 35391 30685 35400 30719
rect 35348 30676 35400 30685
rect 35992 30719 36044 30728
rect 35992 30685 36001 30719
rect 36001 30685 36035 30719
rect 36035 30685 36044 30719
rect 35992 30676 36044 30685
rect 37924 30719 37976 30728
rect 24124 30608 24176 30660
rect 24676 30651 24728 30660
rect 24676 30617 24685 30651
rect 24685 30617 24719 30651
rect 24719 30617 24728 30651
rect 24676 30608 24728 30617
rect 3424 30540 3476 30592
rect 5632 30540 5684 30592
rect 6736 30540 6788 30592
rect 7012 30540 7064 30592
rect 10048 30540 10100 30592
rect 15200 30540 15252 30592
rect 19340 30583 19392 30592
rect 19340 30549 19349 30583
rect 19349 30549 19383 30583
rect 19383 30549 19392 30583
rect 19340 30540 19392 30549
rect 20260 30583 20312 30592
rect 20260 30549 20269 30583
rect 20269 30549 20303 30583
rect 20303 30549 20312 30583
rect 20260 30540 20312 30549
rect 22376 30540 22428 30592
rect 25320 30540 25372 30592
rect 26240 30608 26292 30660
rect 31208 30608 31260 30660
rect 33600 30651 33652 30660
rect 33600 30617 33609 30651
rect 33609 30617 33643 30651
rect 33643 30617 33652 30651
rect 33600 30608 33652 30617
rect 35164 30651 35216 30660
rect 35164 30617 35173 30651
rect 35173 30617 35207 30651
rect 35207 30617 35216 30651
rect 35164 30608 35216 30617
rect 28908 30540 28960 30592
rect 30380 30540 30432 30592
rect 33140 30540 33192 30592
rect 33876 30540 33928 30592
rect 37924 30685 37933 30719
rect 37933 30685 37967 30719
rect 37967 30685 37976 30719
rect 37924 30676 37976 30685
rect 38568 30676 38620 30728
rect 38936 30676 38988 30728
rect 58164 30719 58216 30728
rect 58164 30685 58173 30719
rect 58173 30685 58207 30719
rect 58207 30685 58216 30719
rect 58164 30676 58216 30685
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 2136 30379 2188 30388
rect 2136 30345 2145 30379
rect 2145 30345 2179 30379
rect 2179 30345 2188 30379
rect 2136 30336 2188 30345
rect 7380 30379 7432 30388
rect 7380 30345 7389 30379
rect 7389 30345 7423 30379
rect 7423 30345 7432 30379
rect 7380 30336 7432 30345
rect 30196 30336 30248 30388
rect 30380 30336 30432 30388
rect 37648 30336 37700 30388
rect 2872 30268 2924 30320
rect 3332 30268 3384 30320
rect 7564 30268 7616 30320
rect 8392 30268 8444 30320
rect 2780 30243 2832 30252
rect 2780 30209 2789 30243
rect 2789 30209 2823 30243
rect 2823 30209 2832 30243
rect 2780 30200 2832 30209
rect 3148 30200 3200 30252
rect 3424 30243 3476 30252
rect 3424 30209 3433 30243
rect 3433 30209 3467 30243
rect 3467 30209 3476 30243
rect 3424 30200 3476 30209
rect 10968 30268 11020 30320
rect 15660 30311 15712 30320
rect 15660 30277 15669 30311
rect 15669 30277 15703 30311
rect 15703 30277 15712 30311
rect 15660 30268 15712 30277
rect 16120 30268 16172 30320
rect 18052 30311 18104 30320
rect 18052 30277 18061 30311
rect 18061 30277 18095 30311
rect 18095 30277 18104 30311
rect 18052 30268 18104 30277
rect 9864 30200 9916 30252
rect 11060 30200 11112 30252
rect 11704 30200 11756 30252
rect 14556 30200 14608 30252
rect 15016 30243 15068 30252
rect 15016 30209 15025 30243
rect 15025 30209 15059 30243
rect 15059 30209 15068 30243
rect 15016 30200 15068 30209
rect 15200 30243 15252 30252
rect 15200 30209 15209 30243
rect 15209 30209 15243 30243
rect 15243 30209 15252 30243
rect 15200 30200 15252 30209
rect 10048 30132 10100 30184
rect 11888 30132 11940 30184
rect 2688 30064 2740 30116
rect 9220 29996 9272 30048
rect 14280 30064 14332 30116
rect 15844 30200 15896 30252
rect 16580 30200 16632 30252
rect 17408 30200 17460 30252
rect 19248 30268 19300 30320
rect 16764 30132 16816 30184
rect 18512 30243 18564 30252
rect 18512 30209 18521 30243
rect 18521 30209 18555 30243
rect 18555 30209 18564 30243
rect 18512 30200 18564 30209
rect 19340 30243 19392 30252
rect 14740 29996 14792 30048
rect 15568 30064 15620 30116
rect 18604 30132 18656 30184
rect 19340 30209 19349 30243
rect 19349 30209 19383 30243
rect 19383 30209 19392 30243
rect 19340 30200 19392 30209
rect 19708 30268 19760 30320
rect 19984 30268 20036 30320
rect 17960 30064 18012 30116
rect 19616 30132 19668 30184
rect 20444 30268 20496 30320
rect 22560 30268 22612 30320
rect 24216 30311 24268 30320
rect 20996 30243 21048 30252
rect 20996 30209 21005 30243
rect 21005 30209 21039 30243
rect 21039 30209 21048 30243
rect 20996 30200 21048 30209
rect 22376 30243 22428 30252
rect 22376 30209 22410 30243
rect 22410 30209 22428 30243
rect 22376 30200 22428 30209
rect 24216 30277 24225 30311
rect 24225 30277 24259 30311
rect 24259 30277 24268 30311
rect 24216 30268 24268 30277
rect 26240 30268 26292 30320
rect 29276 30311 29328 30320
rect 29276 30277 29285 30311
rect 29285 30277 29319 30311
rect 29319 30277 29328 30311
rect 29276 30268 29328 30277
rect 31024 30311 31076 30320
rect 31024 30277 31033 30311
rect 31033 30277 31067 30311
rect 31067 30277 31076 30311
rect 31024 30268 31076 30277
rect 31208 30268 31260 30320
rect 33140 30268 33192 30320
rect 24492 30243 24544 30252
rect 20260 30132 20312 30184
rect 22100 30175 22152 30184
rect 22100 30141 22109 30175
rect 22109 30141 22143 30175
rect 22143 30141 22152 30175
rect 22100 30132 22152 30141
rect 23204 30132 23256 30184
rect 24492 30209 24501 30243
rect 24501 30209 24535 30243
rect 24535 30209 24544 30243
rect 24492 30200 24544 30209
rect 24952 30200 25004 30252
rect 25320 30243 25372 30252
rect 25320 30209 25329 30243
rect 25329 30209 25363 30243
rect 25363 30209 25372 30243
rect 25320 30200 25372 30209
rect 24860 30132 24912 30184
rect 25504 30243 25556 30252
rect 25504 30209 25513 30243
rect 25513 30209 25547 30243
rect 25547 30209 25556 30243
rect 25504 30200 25556 30209
rect 19708 30064 19760 30116
rect 20628 30064 20680 30116
rect 23388 30064 23440 30116
rect 16672 30039 16724 30048
rect 16672 30005 16681 30039
rect 16681 30005 16715 30039
rect 16715 30005 16724 30039
rect 16672 29996 16724 30005
rect 17500 30039 17552 30048
rect 17500 30005 17509 30039
rect 17509 30005 17543 30039
rect 17543 30005 17552 30039
rect 17500 29996 17552 30005
rect 20168 29996 20220 30048
rect 20444 29996 20496 30048
rect 20812 29996 20864 30048
rect 23848 29996 23900 30048
rect 25320 30064 25372 30116
rect 29552 30200 29604 30252
rect 30932 30243 30984 30252
rect 30932 30209 30941 30243
rect 30941 30209 30975 30243
rect 30975 30209 30984 30243
rect 30932 30200 30984 30209
rect 32036 30200 32088 30252
rect 33416 30200 33468 30252
rect 35532 30200 35584 30252
rect 35900 30243 35952 30252
rect 35900 30209 35909 30243
rect 35909 30209 35943 30243
rect 35943 30209 35952 30243
rect 35900 30200 35952 30209
rect 36360 30268 36412 30320
rect 31208 30064 31260 30116
rect 27804 29996 27856 30048
rect 28816 29996 28868 30048
rect 31392 29996 31444 30048
rect 33232 29996 33284 30048
rect 35164 30132 35216 30184
rect 35808 30132 35860 30184
rect 34244 30064 34296 30116
rect 37924 30064 37976 30116
rect 36544 30039 36596 30048
rect 36544 30005 36553 30039
rect 36553 30005 36587 30039
rect 36587 30005 36596 30039
rect 36544 29996 36596 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2872 29835 2924 29844
rect 2872 29801 2881 29835
rect 2881 29801 2915 29835
rect 2915 29801 2924 29835
rect 2872 29792 2924 29801
rect 7932 29792 7984 29844
rect 8116 29792 8168 29844
rect 10232 29792 10284 29844
rect 10968 29835 11020 29844
rect 10968 29801 10977 29835
rect 10977 29801 11011 29835
rect 11011 29801 11020 29835
rect 10968 29792 11020 29801
rect 11888 29835 11940 29844
rect 11888 29801 11897 29835
rect 11897 29801 11931 29835
rect 11931 29801 11940 29835
rect 11888 29792 11940 29801
rect 18512 29792 18564 29844
rect 19340 29792 19392 29844
rect 13452 29724 13504 29776
rect 15844 29767 15896 29776
rect 15844 29733 15853 29767
rect 15853 29733 15887 29767
rect 15887 29733 15896 29767
rect 15844 29724 15896 29733
rect 17132 29724 17184 29776
rect 25504 29792 25556 29844
rect 27804 29835 27856 29844
rect 27804 29801 27813 29835
rect 27813 29801 27847 29835
rect 27847 29801 27856 29835
rect 27804 29792 27856 29801
rect 29552 29835 29604 29844
rect 29552 29801 29561 29835
rect 29561 29801 29595 29835
rect 29595 29801 29604 29835
rect 29552 29792 29604 29801
rect 22468 29724 22520 29776
rect 3240 29656 3292 29708
rect 3608 29588 3660 29640
rect 8208 29656 8260 29708
rect 11888 29656 11940 29708
rect 4712 29631 4764 29640
rect 4712 29597 4721 29631
rect 4721 29597 4755 29631
rect 4755 29597 4764 29631
rect 4712 29588 4764 29597
rect 9220 29588 9272 29640
rect 10784 29588 10836 29640
rect 12256 29588 12308 29640
rect 17500 29588 17552 29640
rect 17868 29588 17920 29640
rect 19616 29656 19668 29708
rect 20076 29588 20128 29640
rect 20720 29656 20772 29708
rect 22376 29656 22428 29708
rect 22560 29631 22612 29640
rect 22560 29597 22569 29631
rect 22569 29597 22603 29631
rect 22603 29597 22612 29631
rect 22560 29588 22612 29597
rect 25044 29724 25096 29776
rect 31116 29792 31168 29844
rect 35532 29792 35584 29844
rect 23388 29588 23440 29640
rect 23480 29588 23532 29640
rect 24952 29656 25004 29708
rect 25044 29631 25096 29640
rect 25044 29597 25053 29631
rect 25053 29597 25087 29631
rect 25087 29597 25096 29631
rect 25044 29588 25096 29597
rect 25320 29656 25372 29708
rect 4804 29520 4856 29572
rect 10048 29520 10100 29572
rect 4988 29452 5040 29504
rect 9956 29452 10008 29504
rect 11060 29452 11112 29504
rect 17960 29520 18012 29572
rect 18604 29520 18656 29572
rect 19340 29520 19392 29572
rect 20260 29520 20312 29572
rect 16764 29452 16816 29504
rect 17040 29452 17092 29504
rect 17408 29495 17460 29504
rect 17408 29461 17417 29495
rect 17417 29461 17451 29495
rect 17451 29461 17460 29495
rect 17408 29452 17460 29461
rect 20628 29520 20680 29572
rect 20904 29520 20956 29572
rect 23204 29520 23256 29572
rect 24400 29520 24452 29572
rect 27252 29588 27304 29640
rect 27804 29588 27856 29640
rect 28632 29631 28684 29640
rect 28632 29597 28641 29631
rect 28641 29597 28675 29631
rect 28675 29597 28684 29631
rect 28632 29588 28684 29597
rect 28816 29631 28868 29640
rect 28816 29597 28825 29631
rect 28825 29597 28859 29631
rect 28859 29597 28868 29631
rect 28816 29588 28868 29597
rect 29828 29588 29880 29640
rect 30932 29631 30984 29640
rect 30932 29597 30941 29631
rect 30941 29597 30975 29631
rect 30975 29597 30984 29631
rect 30932 29588 30984 29597
rect 33416 29588 33468 29640
rect 35348 29656 35400 29708
rect 37924 29699 37976 29708
rect 37924 29665 37940 29699
rect 37940 29665 37974 29699
rect 37974 29665 37976 29699
rect 37924 29656 37976 29665
rect 34428 29588 34480 29640
rect 36544 29588 36596 29640
rect 58164 29631 58216 29640
rect 58164 29597 58173 29631
rect 58173 29597 58207 29631
rect 58207 29597 58216 29631
rect 58164 29588 58216 29597
rect 22468 29452 22520 29504
rect 23664 29495 23716 29504
rect 23664 29461 23673 29495
rect 23673 29461 23707 29495
rect 23707 29461 23716 29495
rect 23664 29452 23716 29461
rect 24492 29452 24544 29504
rect 33600 29520 33652 29572
rect 33876 29563 33928 29572
rect 33876 29529 33885 29563
rect 33885 29529 33919 29563
rect 33919 29529 33928 29563
rect 33876 29520 33928 29529
rect 35808 29563 35860 29572
rect 35808 29529 35817 29563
rect 35817 29529 35851 29563
rect 35851 29529 35860 29563
rect 35808 29520 35860 29529
rect 35900 29520 35952 29572
rect 36636 29520 36688 29572
rect 33324 29452 33376 29504
rect 34336 29452 34388 29504
rect 36084 29452 36136 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 4620 29248 4672 29300
rect 3976 29180 4028 29232
rect 2688 29044 2740 29096
rect 2964 29155 3016 29164
rect 2964 29121 2973 29155
rect 2973 29121 3007 29155
rect 3007 29121 3016 29155
rect 2964 29112 3016 29121
rect 3148 29155 3200 29164
rect 3148 29121 3157 29155
rect 3157 29121 3191 29155
rect 3191 29121 3200 29155
rect 3148 29112 3200 29121
rect 3424 29112 3476 29164
rect 4712 29180 4764 29232
rect 4804 29112 4856 29164
rect 5172 29112 5224 29164
rect 11612 29248 11664 29300
rect 12808 29291 12860 29300
rect 12808 29257 12817 29291
rect 12817 29257 12851 29291
rect 12851 29257 12860 29291
rect 12808 29248 12860 29257
rect 15844 29248 15896 29300
rect 19892 29248 19944 29300
rect 7932 29223 7984 29232
rect 7932 29189 7941 29223
rect 7941 29189 7975 29223
rect 7975 29189 7984 29223
rect 7932 29180 7984 29189
rect 9404 29180 9456 29232
rect 10600 29180 10652 29232
rect 10968 29223 11020 29232
rect 10968 29189 10977 29223
rect 10977 29189 11011 29223
rect 11011 29189 11020 29223
rect 10968 29180 11020 29189
rect 11060 29180 11112 29232
rect 8208 29112 8260 29164
rect 10876 29112 10928 29164
rect 13360 29155 13412 29164
rect 3516 28976 3568 29028
rect 4712 28976 4764 29028
rect 4896 28976 4948 29028
rect 13360 29121 13369 29155
rect 13369 29121 13403 29155
rect 13403 29121 13412 29155
rect 13360 29112 13412 29121
rect 14372 29180 14424 29232
rect 17868 29223 17920 29232
rect 17868 29189 17877 29223
rect 17877 29189 17911 29223
rect 17911 29189 17920 29223
rect 17868 29180 17920 29189
rect 17960 29180 18012 29232
rect 20076 29223 20128 29232
rect 20076 29189 20085 29223
rect 20085 29189 20119 29223
rect 20119 29189 20128 29223
rect 20076 29180 20128 29189
rect 11704 29044 11756 29096
rect 13820 29155 13872 29164
rect 13820 29121 13834 29155
rect 13834 29121 13868 29155
rect 13868 29121 13872 29155
rect 13820 29112 13872 29121
rect 14280 29112 14332 29164
rect 19984 29112 20036 29164
rect 20260 29248 20312 29300
rect 23756 29248 23808 29300
rect 24400 29248 24452 29300
rect 25044 29248 25096 29300
rect 25228 29291 25280 29300
rect 25228 29257 25237 29291
rect 25237 29257 25271 29291
rect 25271 29257 25280 29291
rect 25228 29248 25280 29257
rect 25596 29248 25648 29300
rect 25872 29248 25924 29300
rect 29552 29248 29604 29300
rect 32312 29248 32364 29300
rect 21916 29180 21968 29232
rect 22192 29223 22244 29232
rect 22192 29189 22201 29223
rect 22201 29189 22235 29223
rect 22235 29189 22244 29223
rect 24492 29223 24544 29232
rect 22192 29180 22244 29189
rect 22376 29155 22428 29164
rect 15384 29044 15436 29096
rect 22376 29121 22385 29155
rect 22385 29121 22419 29155
rect 22419 29121 22428 29155
rect 22376 29112 22428 29121
rect 24492 29189 24501 29223
rect 24501 29189 24535 29223
rect 24535 29189 24544 29223
rect 24492 29180 24544 29189
rect 29460 29223 29512 29232
rect 29460 29189 29469 29223
rect 29469 29189 29503 29223
rect 29503 29189 29512 29223
rect 29460 29180 29512 29189
rect 23204 29112 23256 29164
rect 24308 29155 24360 29164
rect 24308 29121 24317 29155
rect 24317 29121 24351 29155
rect 24351 29121 24360 29155
rect 24308 29112 24360 29121
rect 24584 29112 24636 29164
rect 25412 29155 25464 29164
rect 25412 29121 25421 29155
rect 25421 29121 25455 29155
rect 25455 29121 25464 29155
rect 25412 29112 25464 29121
rect 26148 29155 26200 29164
rect 26148 29121 26157 29155
rect 26157 29121 26191 29155
rect 26191 29121 26200 29155
rect 26148 29112 26200 29121
rect 27344 29112 27396 29164
rect 29368 29155 29420 29164
rect 29368 29121 29377 29155
rect 29377 29121 29411 29155
rect 29411 29121 29420 29155
rect 29368 29112 29420 29121
rect 30748 29180 30800 29232
rect 35532 29248 35584 29300
rect 36452 29291 36504 29300
rect 36452 29257 36461 29291
rect 36461 29257 36495 29291
rect 36495 29257 36504 29291
rect 36452 29248 36504 29257
rect 36636 29248 36688 29300
rect 33876 29223 33928 29232
rect 33876 29189 33885 29223
rect 33885 29189 33919 29223
rect 33919 29189 33928 29223
rect 33876 29180 33928 29189
rect 22560 29044 22612 29096
rect 23664 29044 23716 29096
rect 30472 29112 30524 29164
rect 33416 29112 33468 29164
rect 34612 29180 34664 29232
rect 38568 29180 38620 29232
rect 38752 29180 38804 29232
rect 34520 29155 34572 29164
rect 34520 29121 34529 29155
rect 34529 29121 34563 29155
rect 34563 29121 34572 29155
rect 34520 29112 34572 29121
rect 38016 29112 38068 29164
rect 9956 28976 10008 29028
rect 10968 28976 11020 29028
rect 14924 28976 14976 29028
rect 16120 28976 16172 29028
rect 19340 29019 19392 29028
rect 19340 28985 19349 29019
rect 19349 28985 19383 29019
rect 19383 28985 19392 29019
rect 19340 28976 19392 28985
rect 20260 28976 20312 29028
rect 20536 28976 20588 29028
rect 23112 29019 23164 29028
rect 23112 28985 23121 29019
rect 23121 28985 23155 29019
rect 23155 28985 23164 29019
rect 23112 28976 23164 28985
rect 29184 29019 29236 29028
rect 29184 28985 29193 29019
rect 29193 28985 29227 29019
rect 29227 28985 29236 29019
rect 29184 28976 29236 28985
rect 34244 29044 34296 29096
rect 2504 28951 2556 28960
rect 2504 28917 2513 28951
rect 2513 28917 2547 28951
rect 2547 28917 2556 28951
rect 2504 28908 2556 28917
rect 8208 28908 8260 28960
rect 9496 28951 9548 28960
rect 9496 28917 9505 28951
rect 9505 28917 9539 28951
rect 9539 28917 9548 28951
rect 9496 28908 9548 28917
rect 14832 28908 14884 28960
rect 20904 28951 20956 28960
rect 20904 28917 20913 28951
rect 20913 28917 20947 28951
rect 20947 28917 20956 28951
rect 20904 28908 20956 28917
rect 21824 28951 21876 28960
rect 21824 28917 21833 28951
rect 21833 28917 21867 28951
rect 21867 28917 21876 28951
rect 21824 28908 21876 28917
rect 30104 28908 30156 28960
rect 31208 28976 31260 29028
rect 32588 28976 32640 29028
rect 33508 29019 33560 29028
rect 33508 28985 33517 29019
rect 33517 28985 33551 29019
rect 33551 28985 33560 29019
rect 33508 28976 33560 28985
rect 36268 29044 36320 29096
rect 37924 29087 37976 29096
rect 37924 29053 37933 29087
rect 37933 29053 37967 29087
rect 37967 29053 37976 29087
rect 37924 29044 37976 29053
rect 34244 28908 34296 28960
rect 35808 28976 35860 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 2964 28747 3016 28756
rect 2964 28713 2973 28747
rect 2973 28713 3007 28747
rect 3007 28713 3016 28747
rect 2964 28704 3016 28713
rect 8576 28704 8628 28756
rect 12808 28636 12860 28688
rect 3332 28500 3384 28552
rect 3792 28432 3844 28484
rect 4712 28500 4764 28552
rect 5172 28500 5224 28552
rect 9312 28500 9364 28552
rect 9496 28543 9548 28552
rect 9496 28509 9530 28543
rect 9530 28509 9548 28543
rect 9496 28500 9548 28509
rect 12532 28500 12584 28552
rect 12992 28500 13044 28552
rect 4804 28475 4856 28484
rect 4804 28441 4813 28475
rect 4813 28441 4847 28475
rect 4847 28441 4856 28475
rect 4804 28432 4856 28441
rect 9772 28432 9824 28484
rect 12440 28432 12492 28484
rect 6368 28364 6420 28416
rect 9680 28364 9732 28416
rect 10048 28364 10100 28416
rect 10600 28407 10652 28416
rect 10600 28373 10609 28407
rect 10609 28373 10643 28407
rect 10643 28373 10652 28407
rect 10600 28364 10652 28373
rect 12900 28407 12952 28416
rect 12900 28373 12909 28407
rect 12909 28373 12943 28407
rect 12943 28373 12952 28407
rect 12900 28364 12952 28373
rect 14556 28500 14608 28552
rect 14832 28543 14884 28552
rect 14832 28509 14841 28543
rect 14841 28509 14875 28543
rect 14875 28509 14884 28543
rect 14832 28500 14884 28509
rect 15568 28704 15620 28756
rect 26792 28704 26844 28756
rect 30104 28704 30156 28756
rect 35808 28704 35860 28756
rect 16856 28636 16908 28688
rect 24768 28636 24820 28688
rect 35532 28636 35584 28688
rect 36268 28636 36320 28688
rect 38016 28704 38068 28756
rect 23756 28568 23808 28620
rect 30748 28611 30800 28620
rect 30748 28577 30757 28611
rect 30757 28577 30791 28611
rect 30791 28577 30800 28611
rect 30748 28568 30800 28577
rect 33416 28568 33468 28620
rect 15844 28543 15896 28552
rect 13452 28432 13504 28484
rect 13912 28432 13964 28484
rect 15844 28509 15853 28543
rect 15853 28509 15887 28543
rect 15887 28509 15896 28543
rect 15844 28500 15896 28509
rect 24860 28500 24912 28552
rect 15200 28432 15252 28484
rect 20720 28432 20772 28484
rect 23480 28475 23532 28484
rect 23480 28441 23489 28475
rect 23489 28441 23523 28475
rect 23523 28441 23532 28475
rect 28908 28500 28960 28552
rect 29368 28500 29420 28552
rect 23480 28432 23532 28441
rect 25412 28432 25464 28484
rect 27160 28432 27212 28484
rect 30472 28500 30524 28552
rect 33784 28543 33836 28552
rect 33784 28509 33793 28543
rect 33793 28509 33827 28543
rect 33827 28509 33836 28543
rect 35900 28568 35952 28620
rect 36084 28568 36136 28620
rect 33784 28500 33836 28509
rect 35440 28500 35492 28552
rect 35992 28543 36044 28552
rect 35992 28509 36001 28543
rect 36001 28509 36035 28543
rect 36035 28509 36044 28543
rect 35992 28500 36044 28509
rect 36452 28500 36504 28552
rect 34428 28432 34480 28484
rect 37280 28475 37332 28484
rect 37280 28441 37289 28475
rect 37289 28441 37323 28475
rect 37323 28441 37332 28475
rect 37280 28432 37332 28441
rect 15292 28407 15344 28416
rect 15292 28373 15301 28407
rect 15301 28373 15335 28407
rect 15335 28373 15344 28407
rect 15292 28364 15344 28373
rect 16948 28407 17000 28416
rect 16948 28373 16957 28407
rect 16957 28373 16991 28407
rect 16991 28373 17000 28407
rect 16948 28364 17000 28373
rect 17960 28364 18012 28416
rect 29000 28407 29052 28416
rect 29000 28373 29009 28407
rect 29009 28373 29043 28407
rect 29043 28373 29052 28407
rect 29000 28364 29052 28373
rect 31484 28407 31536 28416
rect 31484 28373 31493 28407
rect 31493 28373 31527 28407
rect 31527 28373 31536 28407
rect 31484 28364 31536 28373
rect 34704 28407 34756 28416
rect 34704 28373 34713 28407
rect 34713 28373 34747 28407
rect 34747 28373 34756 28407
rect 34704 28364 34756 28373
rect 37464 28407 37516 28416
rect 37464 28373 37473 28407
rect 37473 28373 37507 28407
rect 37507 28373 37516 28407
rect 37464 28364 37516 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 3792 28203 3844 28212
rect 3792 28169 3801 28203
rect 3801 28169 3835 28203
rect 3835 28169 3844 28203
rect 3792 28160 3844 28169
rect 8576 28203 8628 28212
rect 2504 28092 2556 28144
rect 5356 28135 5408 28144
rect 5356 28101 5365 28135
rect 5365 28101 5399 28135
rect 5399 28101 5408 28135
rect 5356 28092 5408 28101
rect 4988 28067 5040 28076
rect 4988 28033 4997 28067
rect 4997 28033 5031 28067
rect 5031 28033 5040 28067
rect 4988 28024 5040 28033
rect 2412 27999 2464 28008
rect 2412 27965 2421 27999
rect 2421 27965 2455 27999
rect 2455 27965 2464 27999
rect 2412 27956 2464 27965
rect 3608 27956 3660 28008
rect 5172 27956 5224 28008
rect 5448 28024 5500 28076
rect 6736 28135 6788 28144
rect 6736 28101 6745 28135
rect 6745 28101 6779 28135
rect 6779 28101 6788 28135
rect 6736 28092 6788 28101
rect 6368 28067 6420 28076
rect 6368 28033 6377 28067
rect 6377 28033 6411 28067
rect 6411 28033 6420 28067
rect 6368 28024 6420 28033
rect 6552 28067 6604 28076
rect 6552 28033 6559 28067
rect 6559 28033 6604 28067
rect 6552 28024 6604 28033
rect 8576 28169 8585 28203
rect 8585 28169 8619 28203
rect 8619 28169 8628 28203
rect 8576 28160 8628 28169
rect 9404 28203 9456 28212
rect 9404 28169 9413 28203
rect 9413 28169 9447 28203
rect 9447 28169 9456 28203
rect 9404 28160 9456 28169
rect 12532 28160 12584 28212
rect 13360 28160 13412 28212
rect 13912 28203 13964 28212
rect 13912 28169 13921 28203
rect 13921 28169 13955 28203
rect 13955 28169 13964 28203
rect 13912 28160 13964 28169
rect 14372 28203 14424 28212
rect 14372 28169 14381 28203
rect 14381 28169 14415 28203
rect 14415 28169 14424 28203
rect 14372 28160 14424 28169
rect 17960 28160 18012 28212
rect 29000 28160 29052 28212
rect 30840 28160 30892 28212
rect 34428 28160 34480 28212
rect 35532 28203 35584 28212
rect 35532 28169 35541 28203
rect 35541 28169 35575 28203
rect 35575 28169 35584 28203
rect 35532 28160 35584 28169
rect 7104 28024 7156 28076
rect 9680 28092 9732 28144
rect 10600 28092 10652 28144
rect 12716 28135 12768 28144
rect 8208 27956 8260 28008
rect 9496 28024 9548 28076
rect 11612 28024 11664 28076
rect 11796 28067 11848 28076
rect 11796 28033 11805 28067
rect 11805 28033 11839 28067
rect 11839 28033 11848 28067
rect 12716 28101 12725 28135
rect 12725 28101 12759 28135
rect 12759 28101 12768 28135
rect 12716 28092 12768 28101
rect 13268 28092 13320 28144
rect 15292 28092 15344 28144
rect 22560 28092 22612 28144
rect 30748 28092 30800 28144
rect 31484 28092 31536 28144
rect 11796 28024 11848 28033
rect 12624 28024 12676 28076
rect 13176 28024 13228 28076
rect 6828 27888 6880 27940
rect 9772 27956 9824 28008
rect 10876 27956 10928 28008
rect 15200 28024 15252 28076
rect 15752 28067 15804 28076
rect 15752 28033 15761 28067
rect 15761 28033 15795 28067
rect 15795 28033 15804 28067
rect 15752 28024 15804 28033
rect 16948 28024 17000 28076
rect 14740 27888 14792 27940
rect 20076 28024 20128 28076
rect 29368 28024 29420 28076
rect 30104 28067 30156 28076
rect 30104 28033 30113 28067
rect 30113 28033 30147 28067
rect 30147 28033 30156 28067
rect 30104 28024 30156 28033
rect 36176 28092 36228 28144
rect 18236 27999 18288 28008
rect 18236 27965 18245 27999
rect 18245 27965 18279 27999
rect 18279 27965 18288 27999
rect 18236 27956 18288 27965
rect 19340 27956 19392 28008
rect 20260 27956 20312 28008
rect 5816 27820 5868 27872
rect 7840 27820 7892 27872
rect 9496 27820 9548 27872
rect 17316 27820 17368 27872
rect 17684 27820 17736 27872
rect 22284 27820 22336 27872
rect 24860 27820 24912 27872
rect 25504 27820 25556 27872
rect 29276 27820 29328 27872
rect 33140 27956 33192 28008
rect 33784 28024 33836 28076
rect 33876 27956 33928 28008
rect 32404 27888 32456 27940
rect 34796 28024 34848 28076
rect 35992 28024 36044 28076
rect 38752 28067 38804 28076
rect 38752 28033 38761 28067
rect 38761 28033 38795 28067
rect 38795 28033 38804 28067
rect 38752 28024 38804 28033
rect 37464 27956 37516 28008
rect 37280 27888 37332 27940
rect 58164 27931 58216 27940
rect 58164 27897 58173 27931
rect 58173 27897 58207 27931
rect 58207 27897 58216 27931
rect 58164 27888 58216 27897
rect 32956 27820 33008 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 11796 27616 11848 27668
rect 12440 27616 12492 27668
rect 5080 27548 5132 27600
rect 4896 27455 4948 27464
rect 4896 27421 4905 27455
rect 4905 27421 4939 27455
rect 4939 27421 4948 27455
rect 4896 27412 4948 27421
rect 5172 27455 5224 27464
rect 3056 27344 3108 27396
rect 5172 27421 5181 27455
rect 5181 27421 5215 27455
rect 5215 27421 5224 27455
rect 5172 27412 5224 27421
rect 8484 27548 8536 27600
rect 6552 27480 6604 27532
rect 5448 27412 5500 27464
rect 6460 27412 6512 27464
rect 7012 27455 7064 27464
rect 5632 27344 5684 27396
rect 7012 27421 7021 27455
rect 7021 27421 7055 27455
rect 7055 27421 7064 27455
rect 7012 27412 7064 27421
rect 7104 27455 7156 27464
rect 8208 27480 8260 27532
rect 9312 27480 9364 27532
rect 7104 27421 7118 27455
rect 7118 27421 7152 27455
rect 7152 27421 7156 27455
rect 7104 27412 7156 27421
rect 6828 27344 6880 27396
rect 7748 27387 7800 27396
rect 7748 27353 7757 27387
rect 7757 27353 7791 27387
rect 7791 27353 7800 27387
rect 7748 27344 7800 27353
rect 9220 27455 9272 27464
rect 9220 27421 9229 27455
rect 9229 27421 9263 27455
rect 9263 27421 9272 27455
rect 9220 27412 9272 27421
rect 9496 27412 9548 27464
rect 10876 27455 10928 27464
rect 10876 27421 10885 27455
rect 10885 27421 10919 27455
rect 10919 27421 10928 27455
rect 10876 27412 10928 27421
rect 11152 27455 11204 27464
rect 11152 27421 11161 27455
rect 11161 27421 11195 27455
rect 11195 27421 11204 27455
rect 11152 27412 11204 27421
rect 12164 27455 12216 27464
rect 12164 27421 12173 27455
rect 12173 27421 12207 27455
rect 12207 27421 12216 27455
rect 12164 27412 12216 27421
rect 12900 27412 12952 27464
rect 14740 27412 14792 27464
rect 17960 27548 18012 27600
rect 22376 27548 22428 27600
rect 16672 27455 16724 27464
rect 16672 27421 16681 27455
rect 16681 27421 16715 27455
rect 16715 27421 16724 27455
rect 16672 27412 16724 27421
rect 16580 27387 16632 27396
rect 16580 27353 16589 27387
rect 16589 27353 16623 27387
rect 16623 27353 16632 27387
rect 25320 27480 25372 27532
rect 30104 27480 30156 27532
rect 20720 27412 20772 27464
rect 21272 27412 21324 27464
rect 27252 27412 27304 27464
rect 16580 27344 16632 27353
rect 20996 27344 21048 27396
rect 22560 27344 22612 27396
rect 25412 27344 25464 27396
rect 33324 27412 33376 27464
rect 30840 27344 30892 27396
rect 34612 27344 34664 27396
rect 7932 27276 7984 27328
rect 8116 27319 8168 27328
rect 8116 27285 8125 27319
rect 8125 27285 8159 27319
rect 8159 27285 8168 27319
rect 8116 27276 8168 27285
rect 8392 27276 8444 27328
rect 17684 27319 17736 27328
rect 17684 27285 17693 27319
rect 17693 27285 17727 27319
rect 17727 27285 17736 27319
rect 17684 27276 17736 27285
rect 21916 27276 21968 27328
rect 22744 27276 22796 27328
rect 24768 27276 24820 27328
rect 29000 27276 29052 27328
rect 29920 27319 29972 27328
rect 29920 27285 29929 27319
rect 29929 27285 29963 27319
rect 29963 27285 29972 27319
rect 29920 27276 29972 27285
rect 33692 27276 33744 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 6552 27072 6604 27124
rect 10508 27072 10560 27124
rect 20812 27072 20864 27124
rect 3608 27047 3660 27056
rect 3608 27013 3617 27047
rect 3617 27013 3651 27047
rect 3651 27013 3660 27047
rect 3608 27004 3660 27013
rect 3240 26936 3292 26988
rect 5448 26936 5500 26988
rect 7932 26979 7984 26988
rect 7932 26945 7950 26979
rect 7950 26945 7984 26979
rect 7932 26936 7984 26945
rect 8208 26979 8260 26988
rect 8208 26945 8217 26979
rect 8217 26945 8251 26979
rect 8251 26945 8260 26979
rect 8208 26936 8260 26945
rect 9220 26936 9272 26988
rect 12716 26936 12768 26988
rect 13176 26979 13228 26988
rect 13176 26945 13185 26979
rect 13185 26945 13219 26979
rect 13219 26945 13228 26979
rect 13176 26936 13228 26945
rect 18696 27004 18748 27056
rect 17500 26936 17552 26988
rect 22100 27004 22152 27056
rect 22928 27004 22980 27056
rect 19248 26936 19300 26988
rect 23480 26979 23532 26988
rect 25044 27072 25096 27124
rect 25412 27115 25464 27124
rect 25412 27081 25421 27115
rect 25421 27081 25455 27115
rect 25455 27081 25464 27115
rect 25412 27072 25464 27081
rect 29368 27072 29420 27124
rect 23480 26945 23498 26979
rect 23498 26945 23532 26979
rect 23480 26936 23532 26945
rect 24768 26979 24820 26988
rect 9956 26868 10008 26920
rect 11152 26868 11204 26920
rect 12440 26868 12492 26920
rect 8300 26800 8352 26852
rect 9312 26800 9364 26852
rect 24768 26945 24777 26979
rect 24777 26945 24811 26979
rect 24811 26945 24820 26979
rect 24768 26936 24820 26945
rect 24584 26868 24636 26920
rect 25320 26936 25372 26988
rect 27436 26936 27488 26988
rect 30932 27004 30984 27056
rect 27988 26936 28040 26988
rect 33784 27072 33836 27124
rect 33324 27004 33376 27056
rect 33048 26936 33100 26988
rect 33232 26936 33284 26988
rect 34520 27004 34572 27056
rect 34152 26979 34204 26988
rect 25596 26800 25648 26852
rect 3976 26732 4028 26784
rect 9220 26775 9272 26784
rect 9220 26741 9229 26775
rect 9229 26741 9263 26775
rect 9263 26741 9272 26775
rect 9220 26732 9272 26741
rect 9496 26732 9548 26784
rect 20076 26732 20128 26784
rect 20628 26732 20680 26784
rect 22560 26732 22612 26784
rect 24124 26732 24176 26784
rect 25320 26732 25372 26784
rect 25688 26732 25740 26784
rect 26792 26732 26844 26784
rect 29920 26800 29972 26852
rect 34152 26945 34161 26979
rect 34161 26945 34195 26979
rect 34195 26945 34204 26979
rect 34152 26936 34204 26945
rect 34612 26979 34664 26988
rect 34612 26945 34621 26979
rect 34621 26945 34655 26979
rect 34655 26945 34664 26979
rect 34612 26936 34664 26945
rect 40592 26936 40644 26988
rect 29368 26732 29420 26784
rect 30288 26732 30340 26784
rect 30472 26732 30524 26784
rect 33968 26732 34020 26784
rect 34796 26732 34848 26784
rect 36268 26732 36320 26784
rect 38752 26775 38804 26784
rect 38752 26741 38761 26775
rect 38761 26741 38795 26775
rect 38795 26741 38804 26775
rect 38752 26732 38804 26741
rect 39948 26732 40000 26784
rect 58164 26775 58216 26784
rect 58164 26741 58173 26775
rect 58173 26741 58207 26775
rect 58207 26741 58216 26775
rect 58164 26732 58216 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 4712 26528 4764 26580
rect 4620 26460 4672 26512
rect 3884 26392 3936 26444
rect 7932 26528 7984 26580
rect 11612 26528 11664 26580
rect 13820 26528 13872 26580
rect 8116 26460 8168 26512
rect 19248 26528 19300 26580
rect 20812 26528 20864 26580
rect 22100 26528 22152 26580
rect 3056 26367 3108 26376
rect 3056 26333 3065 26367
rect 3065 26333 3099 26367
rect 3099 26333 3108 26367
rect 3056 26324 3108 26333
rect 3240 26367 3292 26376
rect 3240 26333 3249 26367
rect 3249 26333 3283 26367
rect 3283 26333 3292 26367
rect 3240 26324 3292 26333
rect 4068 26367 4120 26376
rect 4068 26333 4077 26367
rect 4077 26333 4111 26367
rect 4111 26333 4120 26367
rect 4068 26324 4120 26333
rect 3976 26256 4028 26308
rect 4712 26324 4764 26376
rect 3792 26231 3844 26240
rect 3792 26197 3801 26231
rect 3801 26197 3835 26231
rect 3835 26197 3844 26231
rect 3792 26188 3844 26197
rect 6736 26324 6788 26376
rect 7564 26324 7616 26376
rect 22192 26460 22244 26512
rect 12164 26392 12216 26444
rect 17224 26392 17276 26444
rect 17868 26392 17920 26444
rect 5448 26256 5500 26308
rect 7748 26256 7800 26308
rect 8392 26367 8444 26376
rect 8392 26333 8401 26367
rect 8401 26333 8435 26367
rect 8435 26333 8444 26367
rect 8392 26324 8444 26333
rect 12440 26324 12492 26376
rect 16764 26367 16816 26376
rect 16764 26333 16773 26367
rect 16773 26333 16807 26367
rect 16807 26333 16816 26367
rect 16764 26324 16816 26333
rect 9312 26299 9364 26308
rect 9312 26265 9321 26299
rect 9321 26265 9355 26299
rect 9355 26265 9364 26299
rect 9312 26256 9364 26265
rect 12624 26299 12676 26308
rect 12624 26265 12633 26299
rect 12633 26265 12667 26299
rect 12667 26265 12676 26299
rect 12624 26256 12676 26265
rect 7012 26188 7064 26240
rect 14004 26188 14056 26240
rect 16672 26188 16724 26240
rect 17960 26324 18012 26376
rect 18880 26392 18932 26444
rect 20904 26392 20956 26444
rect 18328 26367 18380 26376
rect 18328 26333 18337 26367
rect 18337 26333 18371 26367
rect 18371 26333 18380 26367
rect 18328 26324 18380 26333
rect 18696 26324 18748 26376
rect 20812 26324 20864 26376
rect 24308 26460 24360 26512
rect 25044 26528 25096 26580
rect 25228 26460 25280 26512
rect 24584 26392 24636 26444
rect 25596 26435 25648 26444
rect 20904 26188 20956 26240
rect 24492 26367 24544 26376
rect 22192 26256 22244 26308
rect 24492 26333 24501 26367
rect 24501 26333 24535 26367
rect 24535 26333 24544 26367
rect 24492 26324 24544 26333
rect 24676 26367 24728 26376
rect 24676 26333 24685 26367
rect 24685 26333 24719 26367
rect 24719 26333 24728 26367
rect 24676 26324 24728 26333
rect 25596 26401 25605 26435
rect 25605 26401 25639 26435
rect 25639 26401 25648 26435
rect 25596 26392 25648 26401
rect 29368 26392 29420 26444
rect 29736 26392 29788 26444
rect 29828 26435 29880 26444
rect 29828 26401 29837 26435
rect 29837 26401 29871 26435
rect 29871 26401 29880 26435
rect 29828 26392 29880 26401
rect 25228 26324 25280 26376
rect 27436 26299 27488 26308
rect 22744 26188 22796 26240
rect 27436 26265 27445 26299
rect 27445 26265 27479 26299
rect 27479 26265 27488 26299
rect 27436 26256 27488 26265
rect 29000 26256 29052 26308
rect 32588 26324 32640 26376
rect 26976 26231 27028 26240
rect 26976 26197 26985 26231
rect 26985 26197 27019 26231
rect 27019 26197 27028 26231
rect 26976 26188 27028 26197
rect 30380 26256 30432 26308
rect 30840 26256 30892 26308
rect 33140 26324 33192 26376
rect 33416 26324 33468 26376
rect 33692 26367 33744 26376
rect 33692 26333 33701 26367
rect 33701 26333 33735 26367
rect 33735 26333 33744 26367
rect 35992 26392 36044 26444
rect 33692 26324 33744 26333
rect 34796 26324 34848 26376
rect 29644 26188 29696 26240
rect 33048 26188 33100 26240
rect 33232 26231 33284 26240
rect 33232 26197 33241 26231
rect 33241 26197 33275 26231
rect 33275 26197 33284 26231
rect 33232 26188 33284 26197
rect 34244 26256 34296 26308
rect 38752 26324 38804 26376
rect 36084 26256 36136 26308
rect 37556 26256 37608 26308
rect 41052 26299 41104 26308
rect 41052 26265 41061 26299
rect 41061 26265 41095 26299
rect 41095 26265 41104 26299
rect 41052 26256 41104 26265
rect 40408 26231 40460 26240
rect 40408 26197 40417 26231
rect 40417 26197 40451 26231
rect 40451 26197 40460 26231
rect 40408 26188 40460 26197
rect 40500 26188 40552 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 3608 25984 3660 26036
rect 7472 26027 7524 26036
rect 7472 25993 7481 26027
rect 7481 25993 7515 26027
rect 7515 25993 7524 26027
rect 7472 25984 7524 25993
rect 8392 26027 8444 26036
rect 8392 25993 8401 26027
rect 8401 25993 8435 26027
rect 8435 25993 8444 26027
rect 8392 25984 8444 25993
rect 17500 26027 17552 26036
rect 17500 25993 17509 26027
rect 17509 25993 17543 26027
rect 17543 25993 17552 26027
rect 17500 25984 17552 25993
rect 17868 25984 17920 26036
rect 3792 25916 3844 25968
rect 5448 25959 5500 25968
rect 5448 25925 5457 25959
rect 5457 25925 5491 25959
rect 5491 25925 5500 25959
rect 5448 25916 5500 25925
rect 5632 25959 5684 25968
rect 5632 25925 5641 25959
rect 5641 25925 5675 25959
rect 5675 25925 5684 25959
rect 5632 25916 5684 25925
rect 2412 25848 2464 25900
rect 6092 25848 6144 25900
rect 6552 25848 6604 25900
rect 6705 25894 6757 25903
rect 6705 25860 6726 25894
rect 6726 25860 6757 25894
rect 6705 25851 6757 25860
rect 7012 25891 7064 25900
rect 7012 25857 7021 25891
rect 7021 25857 7055 25891
rect 7055 25857 7064 25891
rect 9772 25916 9824 25968
rect 10048 25916 10100 25968
rect 13912 25916 13964 25968
rect 7012 25848 7064 25857
rect 9680 25848 9732 25900
rect 9496 25780 9548 25832
rect 18328 25916 18380 25968
rect 22100 25984 22152 26036
rect 25228 25984 25280 26036
rect 27988 25984 28040 26036
rect 30840 26027 30892 26036
rect 30840 25993 30849 26027
rect 30849 25993 30883 26027
rect 30883 25993 30892 26027
rect 30840 25984 30892 25993
rect 33140 25984 33192 26036
rect 34520 25984 34572 26036
rect 39948 25984 40000 26036
rect 40592 26027 40644 26036
rect 40592 25993 40601 26027
rect 40601 25993 40635 26027
rect 40635 25993 40644 26027
rect 40592 25984 40644 25993
rect 20628 25916 20680 25968
rect 12992 25848 13044 25900
rect 16580 25848 16632 25900
rect 17224 25848 17276 25900
rect 17684 25848 17736 25900
rect 12624 25712 12676 25764
rect 4160 25644 4212 25696
rect 4988 25644 5040 25696
rect 6460 25644 6512 25696
rect 9036 25644 9088 25696
rect 12992 25644 13044 25696
rect 15108 25780 15160 25832
rect 14188 25644 14240 25696
rect 15292 25644 15344 25696
rect 18880 25848 18932 25900
rect 19156 25848 19208 25900
rect 19984 25848 20036 25900
rect 20996 25916 21048 25968
rect 22192 25848 22244 25900
rect 24584 25916 24636 25968
rect 26884 25916 26936 25968
rect 33232 25916 33284 25968
rect 36084 25959 36136 25968
rect 36084 25925 36102 25959
rect 36102 25925 36136 25959
rect 36084 25916 36136 25925
rect 38660 25916 38712 25968
rect 18880 25712 18932 25764
rect 21824 25712 21876 25764
rect 22100 25712 22152 25764
rect 24492 25848 24544 25900
rect 25780 25891 25832 25900
rect 25780 25857 25784 25891
rect 25784 25857 25818 25891
rect 25818 25857 25832 25891
rect 25780 25848 25832 25857
rect 25872 25891 25924 25900
rect 25872 25857 25881 25891
rect 25881 25857 25915 25891
rect 25915 25857 25924 25891
rect 25872 25848 25924 25857
rect 29000 25848 29052 25900
rect 30932 25848 30984 25900
rect 33048 25848 33100 25900
rect 40040 25848 40092 25900
rect 40408 25916 40460 25968
rect 40868 25891 40920 25900
rect 40868 25857 40877 25891
rect 40877 25857 40911 25891
rect 40911 25857 40920 25891
rect 40868 25848 40920 25857
rect 36360 25823 36412 25832
rect 36360 25789 36369 25823
rect 36369 25789 36403 25823
rect 36403 25789 36412 25823
rect 36360 25780 36412 25789
rect 40592 25780 40644 25832
rect 40960 25712 41012 25764
rect 20996 25644 21048 25696
rect 23204 25687 23256 25696
rect 23204 25653 23213 25687
rect 23213 25653 23247 25687
rect 23247 25653 23256 25687
rect 23204 25644 23256 25653
rect 28172 25687 28224 25696
rect 28172 25653 28181 25687
rect 28181 25653 28215 25687
rect 28215 25653 28224 25687
rect 28172 25644 28224 25653
rect 33324 25644 33376 25696
rect 38844 25644 38896 25696
rect 41052 25644 41104 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 5632 25440 5684 25492
rect 6552 25440 6604 25492
rect 21456 25440 21508 25492
rect 23572 25440 23624 25492
rect 24124 25440 24176 25492
rect 24860 25440 24912 25492
rect 37648 25440 37700 25492
rect 38292 25440 38344 25492
rect 40040 25483 40092 25492
rect 40040 25449 40049 25483
rect 40049 25449 40083 25483
rect 40083 25449 40092 25483
rect 40040 25440 40092 25449
rect 8392 25372 8444 25424
rect 11704 25372 11756 25424
rect 25228 25372 25280 25424
rect 29184 25372 29236 25424
rect 3884 25304 3936 25356
rect 2872 25236 2924 25288
rect 4068 25279 4120 25288
rect 4068 25245 4077 25279
rect 4077 25245 4111 25279
rect 4111 25245 4120 25279
rect 4068 25236 4120 25245
rect 4620 25304 4672 25356
rect 8208 25304 8260 25356
rect 16672 25304 16724 25356
rect 19248 25304 19300 25356
rect 22928 25347 22980 25356
rect 22928 25313 22937 25347
rect 22937 25313 22971 25347
rect 22971 25313 22980 25347
rect 22928 25304 22980 25313
rect 4712 25236 4764 25288
rect 6460 25279 6512 25288
rect 6460 25245 6478 25279
rect 6478 25245 6512 25279
rect 6460 25236 6512 25245
rect 9772 25236 9824 25288
rect 13728 25236 13780 25288
rect 15292 25279 15344 25288
rect 15292 25245 15301 25279
rect 15301 25245 15335 25279
rect 15335 25245 15344 25279
rect 15292 25236 15344 25245
rect 10048 25211 10100 25220
rect 10048 25177 10057 25211
rect 10057 25177 10091 25211
rect 10091 25177 10100 25211
rect 10048 25168 10100 25177
rect 3608 25100 3660 25152
rect 9956 25100 10008 25152
rect 10692 25100 10744 25152
rect 12716 25100 12768 25152
rect 13452 25143 13504 25152
rect 13452 25109 13461 25143
rect 13461 25109 13495 25143
rect 13495 25109 13504 25143
rect 13452 25100 13504 25109
rect 14188 25100 14240 25152
rect 14740 25100 14792 25152
rect 15200 25168 15252 25220
rect 16672 25168 16724 25220
rect 17776 25236 17828 25288
rect 23204 25236 23256 25288
rect 26976 25236 27028 25288
rect 30932 25236 30984 25288
rect 33048 25304 33100 25356
rect 36360 25236 36412 25288
rect 38660 25236 38712 25288
rect 17316 25168 17368 25220
rect 24492 25168 24544 25220
rect 25964 25211 26016 25220
rect 25964 25177 25973 25211
rect 25973 25177 26007 25211
rect 26007 25177 26016 25211
rect 25964 25168 26016 25177
rect 27436 25168 27488 25220
rect 28264 25168 28316 25220
rect 17408 25100 17460 25152
rect 17960 25100 18012 25152
rect 22192 25100 22244 25152
rect 23020 25100 23072 25152
rect 29092 25100 29144 25152
rect 30288 25100 30340 25152
rect 31760 25168 31812 25220
rect 37280 25168 37332 25220
rect 40500 25279 40552 25288
rect 40500 25245 40509 25279
rect 40509 25245 40543 25279
rect 40543 25245 40552 25279
rect 40500 25236 40552 25245
rect 40960 25236 41012 25288
rect 58164 25279 58216 25288
rect 58164 25245 58173 25279
rect 58173 25245 58207 25279
rect 58207 25245 58216 25279
rect 58164 25236 58216 25245
rect 40592 25168 40644 25220
rect 35992 25143 36044 25152
rect 35992 25109 36001 25143
rect 36001 25109 36035 25143
rect 36035 25109 36044 25143
rect 35992 25100 36044 25109
rect 39212 25143 39264 25152
rect 39212 25109 39221 25143
rect 39221 25109 39255 25143
rect 39255 25109 39264 25143
rect 39212 25100 39264 25109
rect 40868 25100 40920 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 4712 24939 4764 24948
rect 4712 24905 4721 24939
rect 4721 24905 4755 24939
rect 4755 24905 4764 24939
rect 4712 24896 4764 24905
rect 7840 24896 7892 24948
rect 10416 24896 10468 24948
rect 10784 24896 10836 24948
rect 11336 24896 11388 24948
rect 12624 24939 12676 24948
rect 12624 24905 12633 24939
rect 12633 24905 12667 24939
rect 12667 24905 12676 24939
rect 12624 24896 12676 24905
rect 2412 24760 2464 24812
rect 3608 24803 3660 24812
rect 3608 24769 3626 24803
rect 3626 24769 3660 24803
rect 3608 24760 3660 24769
rect 4068 24760 4120 24812
rect 3884 24735 3936 24744
rect 3884 24701 3893 24735
rect 3893 24701 3927 24735
rect 3927 24701 3936 24735
rect 3884 24692 3936 24701
rect 5264 24624 5316 24676
rect 10232 24803 10284 24812
rect 10232 24769 10241 24803
rect 10241 24769 10275 24803
rect 10275 24769 10284 24803
rect 10876 24828 10928 24880
rect 14556 24896 14608 24948
rect 15108 24896 15160 24948
rect 15200 24896 15252 24948
rect 10232 24760 10284 24769
rect 11704 24760 11756 24812
rect 12716 24760 12768 24812
rect 12808 24760 12860 24812
rect 14924 24828 14976 24880
rect 24032 24896 24084 24948
rect 27528 24896 27580 24948
rect 30472 24896 30524 24948
rect 11428 24692 11480 24744
rect 13084 24806 13136 24812
rect 13084 24772 13093 24806
rect 13093 24772 13127 24806
rect 13127 24772 13136 24806
rect 13084 24760 13136 24772
rect 13452 24760 13504 24812
rect 14280 24760 14332 24812
rect 16764 24760 16816 24812
rect 17408 24760 17460 24812
rect 18328 24828 18380 24880
rect 21456 24828 21508 24880
rect 2964 24556 3016 24608
rect 7196 24556 7248 24608
rect 9772 24599 9824 24608
rect 9772 24565 9781 24599
rect 9781 24565 9815 24599
rect 9815 24565 9824 24599
rect 9772 24556 9824 24565
rect 11980 24556 12032 24608
rect 12348 24624 12400 24676
rect 12808 24624 12860 24676
rect 12164 24556 12216 24608
rect 13820 24599 13872 24608
rect 13820 24565 13829 24599
rect 13829 24565 13863 24599
rect 13863 24565 13872 24599
rect 13820 24556 13872 24565
rect 18512 24760 18564 24812
rect 18696 24803 18748 24812
rect 18696 24769 18705 24803
rect 18705 24769 18739 24803
rect 18739 24769 18748 24803
rect 18696 24760 18748 24769
rect 21824 24803 21876 24812
rect 21824 24769 21855 24803
rect 21855 24769 21876 24803
rect 21824 24760 21876 24769
rect 22008 24803 22060 24812
rect 22008 24769 22012 24803
rect 22012 24769 22046 24803
rect 22046 24769 22060 24803
rect 22008 24760 22060 24769
rect 23572 24828 23624 24880
rect 28172 24828 28224 24880
rect 31024 24828 31076 24880
rect 32956 24828 33008 24880
rect 38292 24871 38344 24880
rect 38292 24837 38301 24871
rect 38301 24837 38335 24871
rect 38335 24837 38344 24871
rect 38292 24828 38344 24837
rect 22836 24760 22888 24812
rect 23020 24803 23072 24812
rect 23020 24769 23030 24803
rect 23030 24769 23064 24803
rect 23064 24769 23072 24803
rect 23204 24803 23256 24812
rect 23020 24760 23072 24769
rect 23204 24769 23213 24803
rect 23213 24769 23247 24803
rect 23247 24769 23256 24803
rect 23204 24760 23256 24769
rect 23388 24803 23440 24812
rect 23388 24769 23402 24803
rect 23402 24769 23436 24803
rect 23436 24769 23440 24803
rect 23388 24760 23440 24769
rect 28264 24760 28316 24812
rect 29460 24760 29512 24812
rect 30932 24760 30984 24812
rect 28908 24692 28960 24744
rect 17132 24624 17184 24676
rect 17684 24624 17736 24676
rect 22100 24624 22152 24676
rect 15476 24556 15528 24608
rect 20904 24556 20956 24608
rect 20996 24556 21048 24608
rect 26056 24624 26108 24676
rect 28356 24624 28408 24676
rect 29092 24624 29144 24676
rect 23480 24556 23532 24608
rect 23572 24599 23624 24608
rect 23572 24565 23581 24599
rect 23581 24565 23615 24599
rect 23615 24565 23624 24599
rect 26240 24599 26292 24608
rect 23572 24556 23624 24565
rect 26240 24565 26249 24599
rect 26249 24565 26283 24599
rect 26283 24565 26292 24599
rect 26240 24556 26292 24565
rect 28816 24599 28868 24608
rect 28816 24565 28825 24599
rect 28825 24565 28859 24599
rect 28859 24565 28868 24599
rect 28816 24556 28868 24565
rect 37372 24599 37424 24608
rect 37372 24565 37381 24599
rect 37381 24565 37415 24599
rect 37415 24565 37424 24599
rect 37372 24556 37424 24565
rect 38660 24556 38712 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 3884 24352 3936 24404
rect 7840 24352 7892 24404
rect 10140 24352 10192 24404
rect 16580 24352 16632 24404
rect 17684 24352 17736 24404
rect 11336 24284 11388 24336
rect 14280 24327 14332 24336
rect 14280 24293 14289 24327
rect 14289 24293 14323 24327
rect 14323 24293 14332 24327
rect 14280 24284 14332 24293
rect 8208 24216 8260 24268
rect 6920 24191 6972 24200
rect 6920 24157 6929 24191
rect 6929 24157 6963 24191
rect 6963 24157 6972 24191
rect 6920 24148 6972 24157
rect 7196 24191 7248 24200
rect 7196 24157 7205 24191
rect 7205 24157 7239 24191
rect 7239 24157 7248 24191
rect 7196 24148 7248 24157
rect 9772 24148 9824 24200
rect 4160 24123 4212 24132
rect 4160 24089 4169 24123
rect 4169 24089 4203 24123
rect 4203 24089 4212 24123
rect 4160 24080 4212 24089
rect 11428 24191 11480 24200
rect 11428 24157 11437 24191
rect 11437 24157 11471 24191
rect 11471 24157 11480 24191
rect 11428 24148 11480 24157
rect 9864 24080 9916 24132
rect 6552 24012 6604 24064
rect 10784 24080 10836 24132
rect 11704 24191 11756 24200
rect 11704 24157 11713 24191
rect 11713 24157 11747 24191
rect 11747 24157 11756 24191
rect 11704 24148 11756 24157
rect 12900 24148 12952 24200
rect 13820 24148 13872 24200
rect 20168 24284 20220 24336
rect 18328 24216 18380 24268
rect 11796 24080 11848 24132
rect 12624 24080 12676 24132
rect 14740 24188 14792 24200
rect 14740 24154 14749 24188
rect 14749 24154 14783 24188
rect 14783 24154 14792 24188
rect 14740 24148 14792 24154
rect 14924 24191 14976 24200
rect 14924 24157 14933 24191
rect 14933 24157 14967 24191
rect 14967 24157 14976 24191
rect 16672 24191 16724 24200
rect 14924 24148 14976 24157
rect 16672 24157 16681 24191
rect 16681 24157 16715 24191
rect 16715 24157 16724 24191
rect 16672 24148 16724 24157
rect 17500 24191 17552 24200
rect 17500 24157 17509 24191
rect 17509 24157 17543 24191
rect 17543 24157 17552 24191
rect 17500 24148 17552 24157
rect 15108 24080 15160 24132
rect 16764 24080 16816 24132
rect 17224 24080 17276 24132
rect 18236 24080 18288 24132
rect 19156 24080 19208 24132
rect 10324 24055 10376 24064
rect 10324 24021 10333 24055
rect 10333 24021 10367 24055
rect 10367 24021 10376 24055
rect 10324 24012 10376 24021
rect 11060 24055 11112 24064
rect 11060 24021 11069 24055
rect 11069 24021 11103 24055
rect 11103 24021 11112 24055
rect 11060 24012 11112 24021
rect 13544 24055 13596 24064
rect 13544 24021 13553 24055
rect 13553 24021 13587 24055
rect 13587 24021 13596 24055
rect 13544 24012 13596 24021
rect 14556 24012 14608 24064
rect 15292 24012 15344 24064
rect 20904 24191 20956 24200
rect 20904 24157 20914 24191
rect 20914 24157 20948 24191
rect 20948 24157 20956 24191
rect 28172 24352 28224 24404
rect 29000 24352 29052 24404
rect 31760 24352 31812 24404
rect 37280 24395 37332 24404
rect 37280 24361 37289 24395
rect 37289 24361 37323 24395
rect 37323 24361 37332 24395
rect 37280 24352 37332 24361
rect 22744 24284 22796 24336
rect 26240 24284 26292 24336
rect 22192 24216 22244 24268
rect 20904 24148 20956 24157
rect 21640 24148 21692 24200
rect 25872 24216 25924 24268
rect 22652 24148 22704 24200
rect 24492 24148 24544 24200
rect 20996 24080 21048 24132
rect 21548 24080 21600 24132
rect 21824 24012 21876 24064
rect 21916 24055 21968 24064
rect 21916 24021 21925 24055
rect 21925 24021 21959 24055
rect 21959 24021 21968 24055
rect 23204 24080 23256 24132
rect 24584 24080 24636 24132
rect 24952 24191 25004 24200
rect 24952 24157 24961 24191
rect 24961 24157 24995 24191
rect 24995 24157 25004 24191
rect 24952 24148 25004 24157
rect 25412 24148 25464 24200
rect 26056 24191 26108 24200
rect 26056 24157 26065 24191
rect 26065 24157 26099 24191
rect 26099 24157 26108 24191
rect 26056 24148 26108 24157
rect 26240 24191 26292 24200
rect 26240 24157 26249 24191
rect 26249 24157 26283 24191
rect 26283 24157 26292 24191
rect 29276 24284 29328 24336
rect 30012 24216 30064 24268
rect 26240 24148 26292 24157
rect 28356 24080 28408 24132
rect 28448 24080 28500 24132
rect 28816 24191 28868 24200
rect 28816 24157 28825 24191
rect 28825 24157 28859 24191
rect 28859 24157 28868 24191
rect 28816 24148 28868 24157
rect 30104 24191 30156 24200
rect 25320 24055 25372 24064
rect 21916 24012 21968 24021
rect 25320 24021 25329 24055
rect 25329 24021 25363 24055
rect 25363 24021 25372 24055
rect 25320 24012 25372 24021
rect 25872 24012 25924 24064
rect 28816 24012 28868 24064
rect 30104 24157 30113 24191
rect 30113 24157 30147 24191
rect 30147 24157 30156 24191
rect 30104 24148 30156 24157
rect 30288 24191 30340 24200
rect 30288 24157 30297 24191
rect 30297 24157 30331 24191
rect 30331 24157 30340 24191
rect 30288 24148 30340 24157
rect 33600 24284 33652 24336
rect 40868 24352 40920 24404
rect 35992 24148 36044 24200
rect 37372 24148 37424 24200
rect 40960 24284 41012 24336
rect 38752 24216 38804 24268
rect 31576 24012 31628 24064
rect 37556 24012 37608 24064
rect 38568 24148 38620 24200
rect 58164 24191 58216 24200
rect 58164 24157 58173 24191
rect 58173 24157 58207 24191
rect 58207 24157 58216 24191
rect 58164 24148 58216 24157
rect 39580 24080 39632 24132
rect 39856 24080 39908 24132
rect 40592 24012 40644 24064
rect 41052 24012 41104 24064
rect 41512 24055 41564 24064
rect 41512 24021 41521 24055
rect 41521 24021 41555 24055
rect 41555 24021 41564 24055
rect 41512 24012 41564 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 4160 23808 4212 23860
rect 9312 23808 9364 23860
rect 9772 23851 9824 23860
rect 9772 23817 9781 23851
rect 9781 23817 9815 23851
rect 9815 23817 9824 23851
rect 9772 23808 9824 23817
rect 10048 23808 10100 23860
rect 13084 23808 13136 23860
rect 13452 23808 13504 23860
rect 14924 23808 14976 23860
rect 11060 23740 11112 23792
rect 1952 23672 2004 23724
rect 3240 23672 3292 23724
rect 7840 23715 7892 23724
rect 7840 23681 7849 23715
rect 7849 23681 7883 23715
rect 7883 23681 7892 23715
rect 7840 23672 7892 23681
rect 8208 23672 8260 23724
rect 10508 23715 10560 23724
rect 10508 23681 10517 23715
rect 10517 23681 10551 23715
rect 10551 23681 10560 23715
rect 10508 23672 10560 23681
rect 3792 23604 3844 23656
rect 6736 23604 6788 23656
rect 10692 23718 10744 23724
rect 10692 23684 10701 23718
rect 10701 23684 10735 23718
rect 10735 23684 10744 23718
rect 10692 23672 10744 23684
rect 10876 23715 10928 23724
rect 10876 23681 10885 23715
rect 10885 23681 10919 23715
rect 10919 23681 10928 23715
rect 10876 23672 10928 23681
rect 11244 23672 11296 23724
rect 13544 23715 13596 23724
rect 13544 23681 13553 23715
rect 13553 23681 13587 23715
rect 13587 23681 13596 23715
rect 13544 23672 13596 23681
rect 13728 23715 13780 23724
rect 13728 23681 13737 23715
rect 13737 23681 13771 23715
rect 13771 23681 13780 23715
rect 13728 23672 13780 23681
rect 15200 23783 15252 23792
rect 15200 23749 15209 23783
rect 15209 23749 15243 23783
rect 15243 23749 15252 23783
rect 15200 23740 15252 23749
rect 18512 23808 18564 23860
rect 23112 23808 23164 23860
rect 24584 23808 24636 23860
rect 15108 23715 15160 23724
rect 15108 23681 15117 23715
rect 15117 23681 15151 23715
rect 15151 23681 15160 23715
rect 15108 23672 15160 23681
rect 15292 23715 15344 23724
rect 15292 23681 15301 23715
rect 15301 23681 15335 23715
rect 15335 23681 15344 23715
rect 15292 23672 15344 23681
rect 18604 23672 18656 23724
rect 22468 23715 22520 23724
rect 22468 23681 22477 23715
rect 22477 23681 22511 23715
rect 22511 23681 22520 23715
rect 22468 23672 22520 23681
rect 22560 23715 22612 23724
rect 22560 23681 22570 23715
rect 22570 23681 22604 23715
rect 22604 23681 22612 23715
rect 22560 23672 22612 23681
rect 11428 23604 11480 23656
rect 12900 23647 12952 23656
rect 12900 23613 12909 23647
rect 12909 23613 12943 23647
rect 12943 23613 12952 23647
rect 12900 23604 12952 23613
rect 15476 23604 15528 23656
rect 15660 23604 15712 23656
rect 20996 23604 21048 23656
rect 23204 23740 23256 23792
rect 24492 23783 24544 23792
rect 24492 23749 24501 23783
rect 24501 23749 24535 23783
rect 24535 23749 24544 23783
rect 24492 23740 24544 23749
rect 23388 23672 23440 23724
rect 25596 23740 25648 23792
rect 29092 23808 29144 23860
rect 29460 23851 29512 23860
rect 29460 23817 29469 23851
rect 29469 23817 29503 23851
rect 29503 23817 29512 23851
rect 29460 23808 29512 23817
rect 25320 23715 25372 23724
rect 25320 23681 25354 23715
rect 25354 23681 25372 23715
rect 25320 23672 25372 23681
rect 17408 23536 17460 23588
rect 19156 23536 19208 23588
rect 21640 23536 21692 23588
rect 23388 23536 23440 23588
rect 2688 23468 2740 23520
rect 11612 23468 11664 23520
rect 13636 23468 13688 23520
rect 15384 23468 15436 23520
rect 22836 23468 22888 23520
rect 27620 23740 27672 23792
rect 28908 23740 28960 23792
rect 38752 23808 38804 23860
rect 40868 23808 40920 23860
rect 26056 23468 26108 23520
rect 28264 23672 28316 23724
rect 38660 23740 38712 23792
rect 39764 23740 39816 23792
rect 30104 23715 30156 23724
rect 30104 23681 30113 23715
rect 30113 23681 30147 23715
rect 30147 23681 30156 23715
rect 35900 23715 35952 23724
rect 30104 23672 30156 23681
rect 35900 23681 35909 23715
rect 35909 23681 35943 23715
rect 35943 23681 35952 23715
rect 35900 23672 35952 23681
rect 36176 23672 36228 23724
rect 30012 23604 30064 23656
rect 36360 23672 36412 23724
rect 39580 23672 39632 23724
rect 38844 23604 38896 23656
rect 40868 23715 40920 23724
rect 40868 23681 40877 23715
rect 40877 23681 40911 23715
rect 40911 23681 40920 23715
rect 40868 23672 40920 23681
rect 40776 23604 40828 23656
rect 41052 23715 41104 23724
rect 41052 23681 41061 23715
rect 41061 23681 41095 23715
rect 41095 23681 41104 23715
rect 41052 23672 41104 23681
rect 41236 23715 41288 23724
rect 41236 23681 41245 23715
rect 41245 23681 41279 23715
rect 41279 23681 41288 23715
rect 41236 23672 41288 23681
rect 30012 23468 30064 23520
rect 31576 23536 31628 23588
rect 37188 23536 37240 23588
rect 37464 23536 37516 23588
rect 38568 23536 38620 23588
rect 33784 23468 33836 23520
rect 37740 23468 37792 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 4068 23264 4120 23316
rect 4528 23264 4580 23316
rect 4804 23307 4856 23316
rect 4804 23273 4813 23307
rect 4813 23273 4847 23307
rect 4847 23273 4856 23307
rect 4804 23264 4856 23273
rect 5080 23264 5132 23316
rect 10232 23307 10284 23316
rect 10232 23273 10241 23307
rect 10241 23273 10275 23307
rect 10275 23273 10284 23307
rect 10232 23264 10284 23273
rect 11796 23264 11848 23316
rect 20444 23264 20496 23316
rect 20996 23264 21048 23316
rect 21364 23264 21416 23316
rect 5540 23196 5592 23248
rect 5724 23196 5776 23248
rect 7840 23239 7892 23248
rect 2780 23103 2832 23112
rect 2780 23069 2789 23103
rect 2789 23069 2823 23103
rect 2823 23069 2832 23103
rect 2780 23060 2832 23069
rect 2964 23103 3016 23112
rect 2964 23069 2973 23103
rect 2973 23069 3007 23103
rect 3007 23069 3016 23103
rect 2964 23060 3016 23069
rect 7840 23205 7849 23239
rect 7849 23205 7883 23239
rect 7883 23205 7892 23239
rect 7840 23196 7892 23205
rect 11244 23196 11296 23248
rect 11336 23239 11388 23248
rect 11336 23205 11345 23239
rect 11345 23205 11379 23239
rect 11379 23205 11388 23239
rect 11336 23196 11388 23205
rect 12256 23196 12308 23248
rect 16672 23196 16724 23248
rect 9312 23128 9364 23180
rect 2320 22967 2372 22976
rect 2320 22933 2329 22967
rect 2329 22933 2363 22967
rect 2363 22933 2372 22967
rect 2320 22924 2372 22933
rect 2596 22924 2648 22976
rect 4896 22924 4948 22976
rect 6092 23060 6144 23112
rect 9220 23060 9272 23112
rect 5908 22992 5960 23044
rect 10324 23060 10376 23112
rect 11244 23103 11296 23112
rect 11244 23069 11253 23103
rect 11253 23069 11287 23103
rect 11287 23069 11296 23103
rect 11244 23060 11296 23069
rect 11428 23103 11480 23112
rect 11428 23069 11437 23103
rect 11437 23069 11471 23103
rect 11471 23069 11480 23103
rect 11428 23060 11480 23069
rect 6920 22924 6972 22976
rect 11612 22992 11664 23044
rect 13728 23060 13780 23112
rect 19340 23060 19392 23112
rect 18604 22992 18656 23044
rect 22836 23103 22888 23112
rect 22836 23069 22845 23103
rect 22845 23069 22879 23103
rect 22879 23069 22888 23103
rect 22836 23060 22888 23069
rect 25596 23103 25648 23112
rect 25596 23069 25605 23103
rect 25605 23069 25639 23103
rect 25639 23069 25648 23103
rect 25596 23060 25648 23069
rect 25872 23103 25924 23112
rect 25872 23069 25906 23103
rect 25906 23069 25924 23103
rect 25872 23060 25924 23069
rect 26976 23060 27028 23112
rect 32220 23264 32272 23316
rect 34244 23264 34296 23316
rect 33048 23128 33100 23180
rect 35900 23128 35952 23180
rect 24492 22992 24544 23044
rect 25320 22992 25372 23044
rect 31852 22992 31904 23044
rect 33416 23060 33468 23112
rect 35348 23103 35400 23112
rect 35348 23069 35357 23103
rect 35357 23069 35391 23103
rect 35391 23069 35400 23103
rect 35348 23060 35400 23069
rect 35624 23060 35676 23112
rect 35992 23060 36044 23112
rect 36360 23264 36412 23316
rect 37188 23264 37240 23316
rect 39212 23307 39264 23316
rect 39212 23273 39221 23307
rect 39221 23273 39255 23307
rect 39255 23273 39264 23307
rect 39212 23264 39264 23273
rect 38660 23060 38712 23112
rect 41512 23128 41564 23180
rect 15476 22967 15528 22976
rect 15476 22933 15485 22967
rect 15485 22933 15519 22967
rect 15519 22933 15528 22967
rect 15476 22924 15528 22933
rect 16672 22924 16724 22976
rect 18052 22924 18104 22976
rect 22928 22924 22980 22976
rect 26976 22967 27028 22976
rect 26976 22933 26985 22967
rect 26985 22933 27019 22967
rect 27019 22933 27028 22967
rect 26976 22924 27028 22933
rect 28172 22924 28224 22976
rect 28816 22924 28868 22976
rect 33232 22992 33284 23044
rect 33324 22992 33376 23044
rect 37280 23035 37332 23044
rect 32772 22967 32824 22976
rect 32772 22933 32781 22967
rect 32781 22933 32815 22967
rect 32815 22933 32824 22967
rect 32772 22924 32824 22933
rect 34520 22924 34572 22976
rect 37280 23001 37298 23035
rect 37298 23001 37332 23035
rect 37280 22992 37332 23001
rect 41236 23060 41288 23112
rect 36360 22924 36412 22976
rect 40040 22924 40092 22976
rect 40776 22924 40828 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 2780 22720 2832 22772
rect 5724 22763 5776 22772
rect 5724 22729 5733 22763
rect 5733 22729 5767 22763
rect 5767 22729 5776 22763
rect 5724 22720 5776 22729
rect 5908 22720 5960 22772
rect 1952 22695 2004 22704
rect 1952 22661 1961 22695
rect 1961 22661 1995 22695
rect 1995 22661 2004 22695
rect 1952 22652 2004 22661
rect 2320 22652 2372 22704
rect 3792 22652 3844 22704
rect 2412 22627 2464 22636
rect 2412 22593 2421 22627
rect 2421 22593 2455 22627
rect 2455 22593 2464 22627
rect 2412 22584 2464 22593
rect 4528 22627 4580 22636
rect 4528 22593 4537 22627
rect 4537 22593 4571 22627
rect 4571 22593 4580 22627
rect 4528 22584 4580 22593
rect 4712 22627 4764 22636
rect 4712 22593 4721 22627
rect 4721 22593 4755 22627
rect 4755 22593 4764 22627
rect 4712 22584 4764 22593
rect 4896 22627 4948 22636
rect 4896 22593 4905 22627
rect 4905 22593 4939 22627
rect 4939 22593 4948 22627
rect 9864 22720 9916 22772
rect 10508 22720 10560 22772
rect 11244 22720 11296 22772
rect 13820 22720 13872 22772
rect 15108 22720 15160 22772
rect 19340 22720 19392 22772
rect 20444 22720 20496 22772
rect 7840 22652 7892 22704
rect 14556 22695 14608 22704
rect 14556 22661 14565 22695
rect 14565 22661 14599 22695
rect 14599 22661 14608 22695
rect 14556 22652 14608 22661
rect 22284 22720 22336 22772
rect 26240 22720 26292 22772
rect 27620 22720 27672 22772
rect 33324 22763 33376 22772
rect 4896 22584 4948 22593
rect 5540 22516 5592 22568
rect 6644 22516 6696 22568
rect 14832 22627 14884 22636
rect 14832 22593 14841 22627
rect 14841 22593 14875 22627
rect 14875 22593 14884 22627
rect 14832 22584 14884 22593
rect 15292 22584 15344 22636
rect 18512 22627 18564 22636
rect 18512 22593 18546 22627
rect 18546 22593 18564 22627
rect 18512 22584 18564 22593
rect 21824 22627 21876 22636
rect 16672 22516 16724 22568
rect 21824 22593 21833 22627
rect 21833 22593 21867 22627
rect 21867 22593 21876 22627
rect 21824 22584 21876 22593
rect 22008 22627 22060 22636
rect 22008 22593 22017 22627
rect 22017 22593 22051 22627
rect 22051 22593 22060 22627
rect 22008 22584 22060 22593
rect 23572 22584 23624 22636
rect 24952 22584 25004 22636
rect 23112 22516 23164 22568
rect 4620 22380 4672 22432
rect 16120 22448 16172 22500
rect 8392 22380 8444 22432
rect 14280 22423 14332 22432
rect 14280 22389 14289 22423
rect 14289 22389 14323 22423
rect 14323 22389 14332 22423
rect 14280 22380 14332 22389
rect 15752 22380 15804 22432
rect 17408 22380 17460 22432
rect 17776 22380 17828 22432
rect 21088 22423 21140 22432
rect 21088 22389 21097 22423
rect 21097 22389 21131 22423
rect 21131 22389 21140 22423
rect 21088 22380 21140 22389
rect 21732 22380 21784 22432
rect 22468 22380 22520 22432
rect 22560 22380 22612 22432
rect 23388 22380 23440 22432
rect 26976 22652 27028 22704
rect 32588 22652 32640 22704
rect 33324 22729 33333 22763
rect 33333 22729 33367 22763
rect 33367 22729 33376 22763
rect 33324 22720 33376 22729
rect 33508 22720 33560 22772
rect 37280 22763 37332 22772
rect 25964 22627 26016 22636
rect 25964 22593 25973 22627
rect 25973 22593 26007 22627
rect 26007 22593 26016 22627
rect 25964 22584 26016 22593
rect 27988 22627 28040 22636
rect 27988 22593 28022 22627
rect 28022 22593 28040 22627
rect 27988 22584 28040 22593
rect 31852 22584 31904 22636
rect 32496 22584 32548 22636
rect 32864 22627 32916 22636
rect 32864 22593 32873 22627
rect 32873 22593 32907 22627
rect 32907 22593 32916 22627
rect 32864 22584 32916 22593
rect 25596 22516 25648 22568
rect 32128 22516 32180 22568
rect 33140 22584 33192 22636
rect 34060 22627 34112 22636
rect 34060 22593 34069 22627
rect 34069 22593 34103 22627
rect 34103 22593 34112 22627
rect 34060 22584 34112 22593
rect 34244 22584 34296 22636
rect 37280 22729 37289 22763
rect 37289 22729 37323 22763
rect 37323 22729 37332 22763
rect 37280 22720 37332 22729
rect 37464 22652 37516 22704
rect 35900 22627 35952 22636
rect 35900 22593 35909 22627
rect 35909 22593 35943 22627
rect 35943 22593 35952 22627
rect 35900 22584 35952 22593
rect 33600 22516 33652 22568
rect 34612 22516 34664 22568
rect 35624 22516 35676 22568
rect 36176 22584 36228 22636
rect 36268 22627 36320 22636
rect 36268 22593 36277 22627
rect 36277 22593 36311 22627
rect 36311 22593 36320 22627
rect 36268 22584 36320 22593
rect 37372 22584 37424 22636
rect 40776 22720 40828 22772
rect 39764 22652 39816 22704
rect 37740 22627 37792 22636
rect 37740 22593 37749 22627
rect 37749 22593 37783 22627
rect 37783 22593 37792 22627
rect 37740 22584 37792 22593
rect 36636 22516 36688 22568
rect 40040 22584 40092 22636
rect 29092 22423 29144 22432
rect 29092 22389 29101 22423
rect 29101 22389 29135 22423
rect 29135 22389 29144 22423
rect 29092 22380 29144 22389
rect 30012 22380 30064 22432
rect 32128 22423 32180 22432
rect 32128 22389 32137 22423
rect 32137 22389 32171 22423
rect 32171 22389 32180 22423
rect 32128 22380 32180 22389
rect 32680 22448 32732 22500
rect 32864 22448 32916 22500
rect 38752 22491 38804 22500
rect 38752 22457 38761 22491
rect 38761 22457 38795 22491
rect 38795 22457 38804 22491
rect 38752 22448 38804 22457
rect 58164 22491 58216 22500
rect 58164 22457 58173 22491
rect 58173 22457 58207 22491
rect 58207 22457 58216 22491
rect 58164 22448 58216 22457
rect 33508 22380 33560 22432
rect 34428 22380 34480 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 2596 22176 2648 22228
rect 5540 22176 5592 22228
rect 9680 22176 9732 22228
rect 6000 22083 6052 22092
rect 6000 22049 6009 22083
rect 6009 22049 6043 22083
rect 6043 22049 6052 22083
rect 6000 22040 6052 22049
rect 14832 22108 14884 22160
rect 16580 22176 16632 22228
rect 17408 22108 17460 22160
rect 17868 22108 17920 22160
rect 18512 22151 18564 22160
rect 18512 22117 18521 22151
rect 18521 22117 18555 22151
rect 18555 22117 18564 22151
rect 18512 22108 18564 22117
rect 20352 22176 20404 22228
rect 22652 22176 22704 22228
rect 23388 22176 23440 22228
rect 33508 22219 33560 22228
rect 33508 22185 33517 22219
rect 33517 22185 33551 22219
rect 33551 22185 33560 22219
rect 33508 22176 33560 22185
rect 37372 22176 37424 22228
rect 28080 22108 28132 22160
rect 3884 21972 3936 22024
rect 2228 21904 2280 21956
rect 4620 21904 4672 21956
rect 5632 21904 5684 21956
rect 8392 21972 8444 22024
rect 10416 21972 10468 22024
rect 11244 22015 11296 22024
rect 11244 21981 11253 22015
rect 11253 21981 11287 22015
rect 11287 21981 11296 22015
rect 11520 22015 11572 22024
rect 11244 21972 11296 21981
rect 11520 21981 11529 22015
rect 11529 21981 11563 22015
rect 11563 21981 11572 22015
rect 11520 21972 11572 21981
rect 11704 22040 11756 22092
rect 14096 21972 14148 22024
rect 17776 22040 17828 22092
rect 15752 22015 15804 22024
rect 15752 21981 15761 22015
rect 15761 21981 15795 22015
rect 15795 21981 15804 22015
rect 15752 21972 15804 21981
rect 17224 21972 17276 22024
rect 17868 22015 17920 22024
rect 17868 21981 17877 22015
rect 17877 21981 17911 22015
rect 17911 21981 17920 22015
rect 17868 21972 17920 21981
rect 18052 22015 18104 22024
rect 18052 21981 18061 22015
rect 18061 21981 18095 22015
rect 18095 21981 18104 22015
rect 18052 21972 18104 21981
rect 32956 22040 33008 22092
rect 6368 21904 6420 21956
rect 8944 21904 8996 21956
rect 10048 21947 10100 21956
rect 10048 21913 10057 21947
rect 10057 21913 10091 21947
rect 10091 21913 10100 21947
rect 10048 21904 10100 21913
rect 10324 21904 10376 21956
rect 11428 21947 11480 21956
rect 11428 21913 11437 21947
rect 11437 21913 11471 21947
rect 11471 21913 11480 21947
rect 11428 21904 11480 21913
rect 11704 21904 11756 21956
rect 16120 21904 16172 21956
rect 17500 21904 17552 21956
rect 18880 21972 18932 22024
rect 3240 21879 3292 21888
rect 3240 21845 3249 21879
rect 3249 21845 3283 21879
rect 3283 21845 3292 21879
rect 3240 21836 3292 21845
rect 3976 21836 4028 21888
rect 9956 21836 10008 21888
rect 10968 21836 11020 21888
rect 12624 21836 12676 21888
rect 14924 21879 14976 21888
rect 14924 21845 14933 21879
rect 14933 21845 14967 21879
rect 14967 21845 14976 21879
rect 14924 21836 14976 21845
rect 16948 21836 17000 21888
rect 19340 21836 19392 21888
rect 21916 21972 21968 22024
rect 20260 21904 20312 21956
rect 22560 21972 22612 22024
rect 23112 21975 23118 22002
rect 23118 21975 23152 22002
rect 23152 21975 23164 22002
rect 23112 21950 23164 21975
rect 23204 22015 23256 22024
rect 23204 21981 23213 22015
rect 23213 21981 23247 22015
rect 23247 21981 23256 22015
rect 23388 22015 23440 22024
rect 23204 21972 23256 21981
rect 23388 21981 23397 22015
rect 23397 21981 23431 22015
rect 23431 21981 23440 22015
rect 23388 21972 23440 21981
rect 24400 21972 24452 22024
rect 29092 21972 29144 22024
rect 30472 21972 30524 22024
rect 32220 22015 32272 22024
rect 32220 21981 32229 22015
rect 32229 21981 32263 22015
rect 32263 21981 32272 22015
rect 32220 21972 32272 21981
rect 32404 22015 32456 22024
rect 32404 21981 32413 22015
rect 32413 21981 32447 22015
rect 32447 21981 32456 22015
rect 32404 21972 32456 21981
rect 33048 21972 33100 22024
rect 34520 22040 34572 22092
rect 33324 22015 33376 22024
rect 33324 21981 33333 22015
rect 33333 21981 33367 22015
rect 33367 21981 33376 22015
rect 33324 21972 33376 21981
rect 34244 21972 34296 22024
rect 28264 21947 28316 21956
rect 28264 21913 28273 21947
rect 28273 21913 28307 21947
rect 28307 21913 28316 21947
rect 28264 21904 28316 21913
rect 32772 21904 32824 21956
rect 22744 21879 22796 21888
rect 22744 21845 22753 21879
rect 22753 21845 22787 21879
rect 22787 21845 22796 21879
rect 22744 21836 22796 21845
rect 25964 21836 26016 21888
rect 28724 21836 28776 21888
rect 34428 21904 34480 21956
rect 33048 21879 33100 21888
rect 33048 21845 33057 21879
rect 33057 21845 33091 21879
rect 33091 21845 33100 21879
rect 33048 21836 33100 21845
rect 36636 21836 36688 21888
rect 40684 21836 40736 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 2228 21675 2280 21684
rect 2228 21641 2237 21675
rect 2237 21641 2271 21675
rect 2271 21641 2280 21675
rect 2228 21632 2280 21641
rect 2596 21632 2648 21684
rect 4712 21632 4764 21684
rect 6368 21675 6420 21684
rect 6368 21641 6377 21675
rect 6377 21641 6411 21675
rect 6411 21641 6420 21675
rect 6368 21632 6420 21641
rect 6460 21632 6512 21684
rect 6828 21632 6880 21684
rect 10048 21632 10100 21684
rect 11428 21632 11480 21684
rect 12164 21675 12216 21684
rect 12164 21641 12173 21675
rect 12173 21641 12207 21675
rect 12207 21641 12216 21675
rect 12164 21632 12216 21641
rect 17868 21632 17920 21684
rect 22100 21632 22152 21684
rect 23204 21632 23256 21684
rect 27988 21632 28040 21684
rect 2504 21539 2556 21548
rect 2504 21505 2513 21539
rect 2513 21505 2547 21539
rect 2547 21505 2556 21539
rect 2504 21496 2556 21505
rect 3976 21607 4028 21616
rect 3976 21573 3985 21607
rect 3985 21573 4019 21607
rect 4019 21573 4028 21607
rect 3976 21564 4028 21573
rect 5632 21607 5684 21616
rect 5632 21573 5641 21607
rect 5641 21573 5675 21607
rect 5675 21573 5684 21607
rect 5632 21564 5684 21573
rect 2688 21539 2740 21548
rect 2688 21505 2697 21539
rect 2697 21505 2731 21539
rect 2731 21505 2740 21539
rect 2688 21496 2740 21505
rect 2964 21496 3016 21548
rect 3792 21539 3844 21548
rect 3792 21505 3801 21539
rect 3801 21505 3835 21539
rect 3835 21505 3844 21539
rect 3792 21496 3844 21505
rect 6460 21496 6512 21548
rect 6736 21539 6788 21548
rect 6736 21505 6745 21539
rect 6745 21505 6779 21539
rect 6779 21505 6788 21539
rect 6736 21496 6788 21505
rect 9772 21564 9824 21616
rect 7012 21539 7064 21548
rect 7012 21505 7021 21539
rect 7021 21505 7055 21539
rect 7055 21505 7064 21539
rect 7012 21496 7064 21505
rect 9956 21539 10008 21548
rect 9956 21505 9965 21539
rect 9965 21505 9999 21539
rect 9999 21505 10008 21539
rect 9956 21496 10008 21505
rect 10048 21496 10100 21548
rect 10416 21496 10468 21548
rect 12164 21496 12216 21548
rect 18604 21564 18656 21616
rect 15476 21539 15528 21548
rect 15476 21505 15485 21539
rect 15485 21505 15519 21539
rect 15519 21505 15528 21539
rect 15476 21496 15528 21505
rect 16948 21539 17000 21548
rect 16948 21505 16982 21539
rect 16982 21505 17000 21539
rect 16948 21496 17000 21505
rect 3240 21428 3292 21480
rect 11244 21428 11296 21480
rect 14924 21428 14976 21480
rect 16672 21471 16724 21480
rect 16672 21437 16681 21471
rect 16681 21437 16715 21471
rect 16715 21437 16724 21471
rect 16672 21428 16724 21437
rect 20352 21496 20404 21548
rect 21088 21496 21140 21548
rect 22652 21539 22704 21548
rect 22652 21505 22661 21539
rect 22661 21505 22695 21539
rect 22695 21505 22704 21539
rect 22652 21496 22704 21505
rect 22836 21539 22888 21548
rect 22836 21505 22845 21539
rect 22845 21505 22879 21539
rect 22879 21505 22888 21539
rect 22836 21496 22888 21505
rect 23112 21564 23164 21616
rect 23664 21564 23716 21616
rect 24400 21564 24452 21616
rect 24492 21564 24544 21616
rect 23940 21539 23992 21548
rect 11520 21360 11572 21412
rect 18880 21428 18932 21480
rect 23940 21505 23949 21539
rect 23949 21505 23983 21539
rect 23983 21505 23992 21539
rect 23940 21496 23992 21505
rect 8944 21335 8996 21344
rect 8944 21301 8953 21335
rect 8953 21301 8987 21335
rect 8987 21301 8996 21335
rect 8944 21292 8996 21301
rect 10784 21292 10836 21344
rect 14464 21292 14516 21344
rect 14648 21335 14700 21344
rect 14648 21301 14657 21335
rect 14657 21301 14691 21335
rect 14691 21301 14700 21335
rect 14648 21292 14700 21301
rect 18880 21335 18932 21344
rect 18880 21301 18889 21335
rect 18889 21301 18923 21335
rect 18923 21301 18932 21335
rect 18880 21292 18932 21301
rect 19248 21360 19300 21412
rect 20260 21360 20312 21412
rect 21088 21292 21140 21344
rect 21180 21292 21232 21344
rect 23848 21428 23900 21480
rect 23204 21360 23256 21412
rect 23296 21335 23348 21344
rect 23296 21301 23305 21335
rect 23305 21301 23339 21335
rect 23339 21301 23348 21335
rect 23296 21292 23348 21301
rect 25688 21292 25740 21344
rect 25964 21292 26016 21344
rect 27620 21496 27672 21548
rect 28445 21539 28497 21548
rect 28445 21505 28454 21539
rect 28454 21505 28488 21539
rect 28488 21505 28497 21539
rect 28445 21496 28497 21505
rect 28724 21632 28776 21684
rect 32680 21632 32732 21684
rect 32956 21632 33008 21684
rect 27712 21428 27764 21480
rect 30932 21496 30984 21548
rect 32772 21564 32824 21616
rect 34704 21632 34756 21684
rect 34336 21564 34388 21616
rect 30288 21471 30340 21480
rect 30288 21437 30297 21471
rect 30297 21437 30331 21471
rect 30331 21437 30340 21471
rect 30288 21428 30340 21437
rect 33784 21496 33836 21548
rect 39396 21496 39448 21548
rect 40684 21539 40736 21548
rect 32772 21428 32824 21480
rect 33692 21428 33744 21480
rect 40684 21505 40693 21539
rect 40693 21505 40727 21539
rect 40727 21505 40736 21539
rect 40684 21496 40736 21505
rect 40592 21428 40644 21480
rect 40868 21539 40920 21548
rect 40868 21505 40877 21539
rect 40877 21505 40911 21539
rect 40911 21505 40920 21539
rect 40868 21496 40920 21505
rect 40500 21360 40552 21412
rect 40960 21360 41012 21412
rect 27620 21335 27672 21344
rect 27620 21301 27629 21335
rect 27629 21301 27663 21335
rect 27663 21301 27672 21335
rect 27620 21292 27672 21301
rect 30104 21335 30156 21344
rect 30104 21301 30113 21335
rect 30113 21301 30147 21335
rect 30147 21301 30156 21335
rect 30104 21292 30156 21301
rect 33232 21335 33284 21344
rect 33232 21301 33241 21335
rect 33241 21301 33275 21335
rect 33275 21301 33284 21335
rect 33232 21292 33284 21301
rect 38568 21335 38620 21344
rect 38568 21301 38577 21335
rect 38577 21301 38611 21335
rect 38611 21301 38620 21335
rect 38568 21292 38620 21301
rect 58164 21335 58216 21344
rect 58164 21301 58173 21335
rect 58173 21301 58207 21335
rect 58207 21301 58216 21335
rect 58164 21292 58216 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 10876 21131 10928 21140
rect 10876 21097 10885 21131
rect 10885 21097 10919 21131
rect 10919 21097 10928 21131
rect 10876 21088 10928 21097
rect 13176 21088 13228 21140
rect 13636 21088 13688 21140
rect 16856 21088 16908 21140
rect 16948 21088 17000 21140
rect 22008 21088 22060 21140
rect 30104 21131 30156 21140
rect 13268 21020 13320 21072
rect 13728 21020 13780 21072
rect 13636 20952 13688 21004
rect 10784 20927 10836 20936
rect 10784 20893 10793 20927
rect 10793 20893 10827 20927
rect 10827 20893 10836 20927
rect 10784 20884 10836 20893
rect 11428 20927 11480 20936
rect 11428 20893 11437 20927
rect 11437 20893 11471 20927
rect 11471 20893 11480 20927
rect 11428 20884 11480 20893
rect 12348 20816 12400 20868
rect 14648 20884 14700 20936
rect 15384 20927 15436 20936
rect 15384 20893 15393 20927
rect 15393 20893 15427 20927
rect 15427 20893 15436 20927
rect 15384 20884 15436 20893
rect 15660 20927 15712 20936
rect 15660 20893 15669 20927
rect 15669 20893 15703 20927
rect 15703 20893 15712 20927
rect 15660 20884 15712 20893
rect 21640 21020 21692 21072
rect 30104 21097 30113 21131
rect 30113 21097 30147 21131
rect 30147 21097 30156 21131
rect 30104 21088 30156 21097
rect 30932 21088 30984 21140
rect 33048 21020 33100 21072
rect 18880 20952 18932 21004
rect 13636 20816 13688 20868
rect 14464 20816 14516 20868
rect 15752 20859 15804 20868
rect 15752 20825 15761 20859
rect 15761 20825 15795 20859
rect 15795 20825 15804 20859
rect 15752 20816 15804 20825
rect 16856 20816 16908 20868
rect 17868 20884 17920 20936
rect 19984 20884 20036 20936
rect 20444 20927 20496 20936
rect 20444 20893 20489 20927
rect 20489 20893 20496 20927
rect 20444 20884 20496 20893
rect 20628 20927 20680 20936
rect 20628 20893 20637 20927
rect 20637 20893 20671 20927
rect 20671 20893 20680 20927
rect 24584 20952 24636 21004
rect 26700 20952 26752 21004
rect 27068 20952 27120 21004
rect 30840 20952 30892 21004
rect 20628 20884 20680 20893
rect 23204 20884 23256 20936
rect 25780 20884 25832 20936
rect 29644 20884 29696 20936
rect 29920 20927 29972 20936
rect 29920 20893 29929 20927
rect 29929 20893 29963 20927
rect 29963 20893 29972 20927
rect 29920 20884 29972 20893
rect 37004 20884 37056 20936
rect 38568 21088 38620 21140
rect 37556 20884 37608 20936
rect 38200 20884 38252 20936
rect 39396 20884 39448 20936
rect 40868 21088 40920 21140
rect 2504 20748 2556 20800
rect 4988 20748 5040 20800
rect 12164 20791 12216 20800
rect 12164 20757 12173 20791
rect 12173 20757 12207 20791
rect 12207 20757 12216 20791
rect 12164 20748 12216 20757
rect 13084 20748 13136 20800
rect 13268 20748 13320 20800
rect 20260 20859 20312 20868
rect 20260 20825 20269 20859
rect 20269 20825 20303 20859
rect 20303 20825 20312 20859
rect 20260 20816 20312 20825
rect 22744 20859 22796 20868
rect 22744 20825 22778 20859
rect 22778 20825 22796 20859
rect 17500 20748 17552 20800
rect 17960 20748 18012 20800
rect 20168 20748 20220 20800
rect 22744 20816 22796 20825
rect 23388 20816 23440 20868
rect 28264 20816 28316 20868
rect 31116 20816 31168 20868
rect 22652 20748 22704 20800
rect 23940 20748 23992 20800
rect 24492 20748 24544 20800
rect 26240 20748 26292 20800
rect 27252 20791 27304 20800
rect 27252 20757 27261 20791
rect 27261 20757 27295 20791
rect 27295 20757 27304 20791
rect 27252 20748 27304 20757
rect 29644 20748 29696 20800
rect 30104 20748 30156 20800
rect 31392 20748 31444 20800
rect 32864 20748 32916 20800
rect 33324 20748 33376 20800
rect 33876 20748 33928 20800
rect 37188 20816 37240 20868
rect 40132 20816 40184 20868
rect 40408 20748 40460 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 11980 20544 12032 20596
rect 13636 20587 13688 20596
rect 13636 20553 13645 20587
rect 13645 20553 13679 20587
rect 13679 20553 13688 20587
rect 13636 20544 13688 20553
rect 15660 20587 15712 20596
rect 15660 20553 15669 20587
rect 15669 20553 15703 20587
rect 15703 20553 15712 20587
rect 15660 20544 15712 20553
rect 20168 20544 20220 20596
rect 29092 20544 29144 20596
rect 29368 20544 29420 20596
rect 31116 20544 31168 20596
rect 31668 20544 31720 20596
rect 40132 20544 40184 20596
rect 40776 20544 40828 20596
rect 5356 20476 5408 20528
rect 12164 20476 12216 20528
rect 7748 20408 7800 20460
rect 13728 20476 13780 20528
rect 12532 20451 12584 20460
rect 12532 20417 12566 20451
rect 12566 20417 12584 20451
rect 12532 20408 12584 20417
rect 13268 20408 13320 20460
rect 15200 20408 15252 20460
rect 15476 20408 15528 20460
rect 19800 20476 19852 20528
rect 23296 20519 23348 20528
rect 23296 20485 23330 20519
rect 23330 20485 23348 20519
rect 23296 20476 23348 20485
rect 17684 20451 17736 20460
rect 17684 20417 17693 20451
rect 17693 20417 17727 20451
rect 17727 20417 17736 20451
rect 17684 20408 17736 20417
rect 19524 20408 19576 20460
rect 19892 20408 19944 20460
rect 20168 20451 20220 20460
rect 20168 20417 20177 20451
rect 20177 20417 20211 20451
rect 20211 20417 20220 20451
rect 20168 20408 20220 20417
rect 20352 20451 20404 20460
rect 20352 20417 20397 20451
rect 20397 20417 20404 20451
rect 20352 20408 20404 20417
rect 20536 20451 20588 20460
rect 20536 20417 20545 20451
rect 20545 20417 20579 20451
rect 20579 20417 20588 20451
rect 20536 20408 20588 20417
rect 23112 20408 23164 20460
rect 27436 20476 27488 20528
rect 12256 20383 12308 20392
rect 9128 20272 9180 20324
rect 9220 20247 9272 20256
rect 9220 20213 9229 20247
rect 9229 20213 9263 20247
rect 9263 20213 9272 20247
rect 9220 20204 9272 20213
rect 12256 20349 12265 20383
rect 12265 20349 12299 20383
rect 12299 20349 12308 20383
rect 12256 20340 12308 20349
rect 14096 20383 14148 20392
rect 14096 20349 14105 20383
rect 14105 20349 14139 20383
rect 14139 20349 14148 20383
rect 14096 20340 14148 20349
rect 17500 20340 17552 20392
rect 24860 20340 24912 20392
rect 26240 20451 26292 20460
rect 26240 20417 26249 20451
rect 26249 20417 26283 20451
rect 26283 20417 26292 20451
rect 26240 20408 26292 20417
rect 26424 20451 26476 20460
rect 26424 20417 26433 20451
rect 26433 20417 26467 20451
rect 26467 20417 26476 20451
rect 26424 20408 26476 20417
rect 26884 20408 26936 20460
rect 27252 20408 27304 20460
rect 28632 20451 28684 20460
rect 28632 20417 28641 20451
rect 28641 20417 28675 20451
rect 28675 20417 28684 20451
rect 28632 20408 28684 20417
rect 29460 20408 29512 20460
rect 32404 20476 32456 20528
rect 32588 20476 32640 20528
rect 31760 20408 31812 20460
rect 32036 20408 32088 20460
rect 32496 20451 32548 20460
rect 32496 20417 32505 20451
rect 32505 20417 32539 20451
rect 32539 20417 32548 20451
rect 32496 20408 32548 20417
rect 32680 20451 32732 20460
rect 32680 20417 32689 20451
rect 32689 20417 32723 20451
rect 32723 20417 32732 20451
rect 32680 20408 32732 20417
rect 32864 20451 32916 20460
rect 32864 20417 32873 20451
rect 32873 20417 32907 20451
rect 32907 20417 32916 20451
rect 40684 20476 40736 20528
rect 32864 20408 32916 20417
rect 36268 20408 36320 20460
rect 40960 20451 41012 20460
rect 40960 20417 40969 20451
rect 40969 20417 41003 20451
rect 41003 20417 41012 20451
rect 40960 20408 41012 20417
rect 41236 20408 41288 20460
rect 28448 20340 28500 20392
rect 29000 20340 29052 20392
rect 29920 20340 29972 20392
rect 27620 20272 27672 20324
rect 32864 20272 32916 20324
rect 11060 20204 11112 20256
rect 11428 20204 11480 20256
rect 16764 20204 16816 20256
rect 16856 20204 16908 20256
rect 17592 20247 17644 20256
rect 17592 20213 17601 20247
rect 17601 20213 17635 20247
rect 17635 20213 17644 20247
rect 17592 20204 17644 20213
rect 19984 20204 20036 20256
rect 24400 20247 24452 20256
rect 24400 20213 24409 20247
rect 24409 20213 24443 20247
rect 24443 20213 24452 20247
rect 24400 20204 24452 20213
rect 25872 20204 25924 20256
rect 26148 20204 26200 20256
rect 29000 20204 29052 20256
rect 29368 20204 29420 20256
rect 30196 20204 30248 20256
rect 32220 20204 32272 20256
rect 33600 20204 33652 20256
rect 37188 20340 37240 20392
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 5724 20000 5776 20052
rect 12532 20043 12584 20052
rect 9588 19796 9640 19848
rect 12532 20009 12541 20043
rect 12541 20009 12575 20043
rect 12575 20009 12584 20043
rect 12532 20000 12584 20009
rect 15016 20000 15068 20052
rect 19524 20043 19576 20052
rect 19524 20009 19533 20043
rect 19533 20009 19567 20043
rect 19567 20009 19576 20043
rect 19524 20000 19576 20009
rect 22836 20000 22888 20052
rect 25780 20000 25832 20052
rect 12716 19864 12768 19916
rect 13268 19864 13320 19916
rect 19892 19864 19944 19916
rect 20536 19864 20588 19916
rect 4804 19728 4856 19780
rect 4620 19703 4672 19712
rect 4620 19669 4629 19703
rect 4629 19669 4663 19703
rect 4663 19669 4672 19703
rect 4620 19660 4672 19669
rect 5356 19660 5408 19712
rect 7840 19728 7892 19780
rect 13084 19796 13136 19848
rect 13176 19839 13228 19848
rect 13176 19805 13185 19839
rect 13185 19805 13219 19839
rect 13219 19805 13228 19839
rect 14832 19839 14884 19848
rect 13176 19796 13228 19805
rect 14832 19805 14841 19839
rect 14841 19805 14875 19839
rect 14875 19805 14884 19839
rect 14832 19796 14884 19805
rect 17960 19796 18012 19848
rect 20076 19839 20128 19848
rect 20076 19805 20084 19839
rect 20084 19805 20118 19839
rect 20118 19805 20128 19839
rect 20076 19796 20128 19805
rect 21180 19796 21232 19848
rect 13728 19728 13780 19780
rect 7656 19660 7708 19712
rect 15016 19660 15068 19712
rect 19892 19771 19944 19780
rect 19892 19737 19901 19771
rect 19901 19737 19935 19771
rect 19935 19737 19944 19771
rect 26976 19864 27028 19916
rect 24400 19796 24452 19848
rect 25688 19796 25740 19848
rect 25872 19839 25924 19848
rect 25872 19805 25906 19839
rect 25906 19805 25924 19839
rect 25872 19796 25924 19805
rect 29736 20000 29788 20052
rect 32128 20000 32180 20052
rect 32680 20000 32732 20052
rect 35348 20000 35400 20052
rect 36084 20000 36136 20052
rect 40960 20000 41012 20052
rect 30196 19932 30248 19984
rect 29000 19796 29052 19848
rect 29644 19839 29696 19848
rect 29644 19805 29653 19839
rect 29653 19805 29687 19839
rect 29687 19805 29696 19839
rect 29644 19796 29696 19805
rect 23664 19771 23716 19780
rect 19892 19728 19944 19737
rect 23664 19737 23673 19771
rect 23673 19737 23707 19771
rect 23707 19737 23716 19771
rect 23664 19728 23716 19737
rect 24676 19728 24728 19780
rect 21088 19660 21140 19712
rect 25872 19660 25924 19712
rect 26424 19660 26476 19712
rect 27620 19660 27672 19712
rect 31116 19932 31168 19984
rect 30472 19796 30524 19848
rect 31760 19864 31812 19916
rect 31484 19839 31536 19848
rect 31484 19805 31493 19839
rect 31493 19805 31527 19839
rect 31527 19805 31536 19839
rect 31484 19796 31536 19805
rect 31668 19796 31720 19848
rect 35348 19839 35400 19848
rect 35348 19805 35357 19839
rect 35357 19805 35391 19839
rect 35391 19805 35400 19839
rect 35348 19796 35400 19805
rect 37832 19932 37884 19984
rect 37004 19796 37056 19848
rect 39304 19839 39356 19848
rect 39304 19805 39313 19839
rect 39313 19805 39347 19839
rect 39347 19805 39356 19839
rect 39304 19796 39356 19805
rect 39856 19796 39908 19848
rect 40408 19839 40460 19848
rect 40408 19805 40417 19839
rect 40417 19805 40451 19839
rect 40451 19805 40460 19839
rect 40408 19796 40460 19805
rect 58164 19839 58216 19848
rect 58164 19805 58173 19839
rect 58173 19805 58207 19839
rect 58207 19805 58216 19839
rect 58164 19796 58216 19805
rect 31208 19771 31260 19780
rect 31208 19737 31217 19771
rect 31217 19737 31251 19771
rect 31251 19737 31260 19771
rect 31208 19728 31260 19737
rect 32128 19728 32180 19780
rect 32772 19771 32824 19780
rect 32772 19737 32781 19771
rect 32781 19737 32815 19771
rect 32815 19737 32824 19771
rect 32772 19728 32824 19737
rect 30932 19703 30984 19712
rect 30932 19669 30941 19703
rect 30941 19669 30975 19703
rect 30975 19669 30984 19703
rect 30932 19660 30984 19669
rect 34520 19660 34572 19712
rect 36268 19728 36320 19780
rect 40132 19728 40184 19780
rect 37372 19660 37424 19712
rect 37924 19703 37976 19712
rect 37924 19669 37933 19703
rect 37933 19669 37967 19703
rect 37967 19669 37976 19703
rect 37924 19660 37976 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 5724 19456 5776 19508
rect 7840 19499 7892 19508
rect 7840 19465 7849 19499
rect 7849 19465 7883 19499
rect 7883 19465 7892 19499
rect 7840 19456 7892 19465
rect 14096 19499 14148 19508
rect 14096 19465 14105 19499
rect 14105 19465 14139 19499
rect 14139 19465 14148 19499
rect 14096 19456 14148 19465
rect 16764 19456 16816 19508
rect 17592 19456 17644 19508
rect 18052 19499 18104 19508
rect 18052 19465 18061 19499
rect 18061 19465 18095 19499
rect 18095 19465 18104 19499
rect 18052 19456 18104 19465
rect 21088 19456 21140 19508
rect 21916 19456 21968 19508
rect 23020 19456 23072 19508
rect 26700 19456 26752 19508
rect 26976 19499 27028 19508
rect 26976 19465 26985 19499
rect 26985 19465 27019 19499
rect 27019 19465 27028 19499
rect 26976 19456 27028 19465
rect 5356 19388 5408 19440
rect 2412 19363 2464 19372
rect 2412 19329 2421 19363
rect 2421 19329 2455 19363
rect 2455 19329 2464 19363
rect 2412 19320 2464 19329
rect 4712 19320 4764 19372
rect 6920 19320 6972 19372
rect 9220 19388 9272 19440
rect 13820 19388 13872 19440
rect 7656 19363 7708 19372
rect 7656 19329 7665 19363
rect 7665 19329 7699 19363
rect 7699 19329 7708 19363
rect 7656 19320 7708 19329
rect 11980 19320 12032 19372
rect 16672 19363 16724 19372
rect 5632 19252 5684 19304
rect 4896 19184 4948 19236
rect 2136 19116 2188 19168
rect 5448 19116 5500 19168
rect 7288 19184 7340 19236
rect 8208 19184 8260 19236
rect 13912 19252 13964 19304
rect 16672 19329 16681 19363
rect 16681 19329 16715 19363
rect 16715 19329 16724 19363
rect 16672 19320 16724 19329
rect 16764 19320 16816 19372
rect 24676 19388 24728 19440
rect 25872 19388 25924 19440
rect 14556 19252 14608 19304
rect 22100 19363 22152 19372
rect 22100 19329 22109 19363
rect 22109 19329 22143 19363
rect 22143 19329 22152 19363
rect 22100 19320 22152 19329
rect 24400 19320 24452 19372
rect 25688 19363 25740 19372
rect 25688 19329 25697 19363
rect 25697 19329 25731 19363
rect 25731 19329 25740 19363
rect 25688 19320 25740 19329
rect 22376 19252 22428 19304
rect 24952 19252 25004 19304
rect 26148 19320 26200 19372
rect 26424 19320 26476 19372
rect 27160 19363 27212 19372
rect 27160 19329 27169 19363
rect 27169 19329 27203 19363
rect 27203 19329 27212 19363
rect 27528 19388 27580 19440
rect 29736 19431 29788 19440
rect 29736 19397 29745 19431
rect 29745 19397 29779 19431
rect 29779 19397 29788 19431
rect 29736 19388 29788 19397
rect 30380 19388 30432 19440
rect 39304 19499 39356 19508
rect 31024 19431 31076 19440
rect 31024 19397 31033 19431
rect 31033 19397 31067 19431
rect 31067 19397 31076 19431
rect 31024 19388 31076 19397
rect 27160 19320 27212 19329
rect 29828 19363 29880 19372
rect 29828 19329 29837 19363
rect 29837 19329 29871 19363
rect 29871 19329 29880 19363
rect 29828 19320 29880 19329
rect 30472 19320 30524 19372
rect 34428 19388 34480 19440
rect 39304 19465 39313 19499
rect 39313 19465 39347 19499
rect 39347 19465 39356 19499
rect 39304 19456 39356 19465
rect 40132 19456 40184 19508
rect 36268 19431 36320 19440
rect 36268 19397 36277 19431
rect 36277 19397 36311 19431
rect 36311 19397 36320 19431
rect 36268 19388 36320 19397
rect 33324 19363 33376 19372
rect 33324 19329 33342 19363
rect 33342 19329 33376 19363
rect 33324 19320 33376 19329
rect 33600 19363 33652 19372
rect 33600 19329 33609 19363
rect 33609 19329 33643 19363
rect 33643 19329 33652 19363
rect 33600 19320 33652 19329
rect 35900 19320 35952 19372
rect 36084 19363 36136 19372
rect 36084 19329 36093 19363
rect 36093 19329 36127 19363
rect 36127 19329 36136 19363
rect 36084 19320 36136 19329
rect 38108 19388 38160 19440
rect 40684 19388 40736 19440
rect 37280 19320 37332 19372
rect 37648 19320 37700 19372
rect 40868 19363 40920 19372
rect 40868 19329 40877 19363
rect 40877 19329 40911 19363
rect 40911 19329 40920 19363
rect 40868 19320 40920 19329
rect 41052 19363 41104 19372
rect 41052 19329 41061 19363
rect 41061 19329 41095 19363
rect 41095 19329 41104 19363
rect 41052 19320 41104 19329
rect 41236 19363 41288 19372
rect 41236 19329 41245 19363
rect 41245 19329 41279 19363
rect 41279 19329 41288 19363
rect 41236 19320 41288 19329
rect 30840 19295 30892 19304
rect 8300 19159 8352 19168
rect 8300 19125 8309 19159
rect 8309 19125 8343 19159
rect 8343 19125 8352 19159
rect 8300 19116 8352 19125
rect 10784 19184 10836 19236
rect 10692 19116 10744 19168
rect 11060 19184 11112 19236
rect 11612 19116 11664 19168
rect 12716 19116 12768 19168
rect 20628 19184 20680 19236
rect 30840 19261 30849 19295
rect 30849 19261 30883 19295
rect 30883 19261 30892 19295
rect 30840 19252 30892 19261
rect 31484 19184 31536 19236
rect 32220 19227 32272 19236
rect 32220 19193 32229 19227
rect 32229 19193 32263 19227
rect 32263 19193 32272 19227
rect 32220 19184 32272 19193
rect 19248 19116 19300 19168
rect 27344 19159 27396 19168
rect 27344 19125 27353 19159
rect 27353 19125 27387 19159
rect 27387 19125 27396 19159
rect 27344 19116 27396 19125
rect 30472 19116 30524 19168
rect 30656 19116 30708 19168
rect 31116 19116 31168 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 5632 18955 5684 18964
rect 5632 18921 5641 18955
rect 5641 18921 5675 18955
rect 5675 18921 5684 18955
rect 5632 18912 5684 18921
rect 6828 18912 6880 18964
rect 12532 18912 12584 18964
rect 13636 18912 13688 18964
rect 15844 18955 15896 18964
rect 15844 18921 15853 18955
rect 15853 18921 15887 18955
rect 15887 18921 15896 18955
rect 15844 18912 15896 18921
rect 16764 18912 16816 18964
rect 20628 18955 20680 18964
rect 20628 18921 20637 18955
rect 20637 18921 20671 18955
rect 20671 18921 20680 18955
rect 20628 18912 20680 18921
rect 26700 18912 26752 18964
rect 27344 18912 27396 18964
rect 6736 18844 6788 18896
rect 1860 18751 1912 18760
rect 1860 18717 1869 18751
rect 1869 18717 1903 18751
rect 1903 18717 1912 18751
rect 1860 18708 1912 18717
rect 2136 18751 2188 18760
rect 2136 18717 2170 18751
rect 2170 18717 2188 18751
rect 2136 18708 2188 18717
rect 4620 18776 4672 18828
rect 7380 18776 7432 18828
rect 5540 18708 5592 18760
rect 6920 18751 6972 18760
rect 6920 18717 6929 18751
rect 6929 18717 6963 18751
rect 6963 18717 6972 18751
rect 6920 18708 6972 18717
rect 7012 18708 7064 18760
rect 4068 18640 4120 18692
rect 4896 18640 4948 18692
rect 3332 18572 3384 18624
rect 4160 18615 4212 18624
rect 4160 18581 4169 18615
rect 4169 18581 4203 18615
rect 4203 18581 4212 18615
rect 4160 18572 4212 18581
rect 5632 18572 5684 18624
rect 7288 18751 7340 18760
rect 7288 18717 7297 18751
rect 7297 18717 7331 18751
rect 7331 18717 7340 18751
rect 10876 18844 10928 18896
rect 7288 18708 7340 18717
rect 9588 18751 9640 18760
rect 9588 18717 9597 18751
rect 9597 18717 9631 18751
rect 9631 18717 9640 18751
rect 9588 18708 9640 18717
rect 11612 18776 11664 18828
rect 23020 18844 23072 18896
rect 27620 18844 27672 18896
rect 30472 18912 30524 18964
rect 30932 18844 30984 18896
rect 11704 18751 11756 18760
rect 11704 18717 11713 18751
rect 11713 18717 11747 18751
rect 11747 18717 11756 18751
rect 11704 18708 11756 18717
rect 11888 18751 11940 18760
rect 11888 18717 11897 18751
rect 11897 18717 11931 18751
rect 11931 18717 11940 18751
rect 13728 18776 13780 18828
rect 11888 18708 11940 18717
rect 15844 18708 15896 18760
rect 10600 18640 10652 18692
rect 16856 18751 16908 18760
rect 16856 18717 16865 18751
rect 16865 18717 16899 18751
rect 16899 18717 16908 18751
rect 16856 18708 16908 18717
rect 17316 18708 17368 18760
rect 18236 18751 18288 18760
rect 18236 18717 18245 18751
rect 18245 18717 18279 18751
rect 18279 18717 18288 18751
rect 18236 18708 18288 18717
rect 17132 18640 17184 18692
rect 18696 18708 18748 18760
rect 20904 18776 20956 18828
rect 21916 18819 21968 18828
rect 21916 18785 21925 18819
rect 21925 18785 21959 18819
rect 21959 18785 21968 18819
rect 21916 18776 21968 18785
rect 23388 18776 23440 18828
rect 30380 18776 30432 18828
rect 30104 18751 30156 18760
rect 6920 18572 6972 18624
rect 7196 18572 7248 18624
rect 7656 18615 7708 18624
rect 7656 18581 7665 18615
rect 7665 18581 7699 18615
rect 7699 18581 7708 18615
rect 7656 18572 7708 18581
rect 11060 18572 11112 18624
rect 20812 18640 20864 18692
rect 26792 18640 26844 18692
rect 25504 18572 25556 18624
rect 26516 18572 26568 18624
rect 27988 18640 28040 18692
rect 30104 18717 30113 18751
rect 30113 18717 30147 18751
rect 30147 18717 30156 18751
rect 30104 18708 30156 18717
rect 30564 18708 30616 18760
rect 30932 18708 30984 18760
rect 31944 18708 31996 18760
rect 32496 18844 32548 18896
rect 33324 18912 33376 18964
rect 34428 18912 34480 18964
rect 41052 18912 41104 18964
rect 34520 18844 34572 18896
rect 32680 18776 32732 18828
rect 27436 18615 27488 18624
rect 27436 18581 27445 18615
rect 27445 18581 27479 18615
rect 27479 18581 27488 18615
rect 27436 18572 27488 18581
rect 28816 18572 28868 18624
rect 29644 18615 29696 18624
rect 29644 18581 29653 18615
rect 29653 18581 29687 18615
rect 29687 18581 29696 18615
rect 29644 18572 29696 18581
rect 30564 18615 30616 18624
rect 30564 18581 30573 18615
rect 30573 18581 30607 18615
rect 30607 18581 30616 18615
rect 30564 18572 30616 18581
rect 31668 18615 31720 18624
rect 31668 18581 31677 18615
rect 31677 18581 31711 18615
rect 31711 18581 31720 18615
rect 37004 18708 37056 18760
rect 37924 18776 37976 18828
rect 38936 18708 38988 18760
rect 58164 18751 58216 18760
rect 58164 18717 58173 18751
rect 58173 18717 58207 18751
rect 58207 18717 58216 18751
rect 58164 18708 58216 18717
rect 37188 18640 37240 18692
rect 38752 18640 38804 18692
rect 39856 18683 39908 18692
rect 39856 18649 39865 18683
rect 39865 18649 39899 18683
rect 39899 18649 39908 18683
rect 39856 18640 39908 18649
rect 31668 18572 31720 18581
rect 40868 18572 40920 18624
rect 41052 18572 41104 18624
rect 41328 18572 41380 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 2412 18368 2464 18420
rect 7196 18368 7248 18420
rect 4068 18300 4120 18352
rect 5632 18300 5684 18352
rect 7012 18300 7064 18352
rect 8300 18368 8352 18420
rect 7656 18300 7708 18352
rect 1676 18275 1728 18284
rect 1676 18241 1685 18275
rect 1685 18241 1719 18275
rect 1719 18241 1728 18275
rect 1676 18232 1728 18241
rect 3332 18232 3384 18284
rect 2412 18164 2464 18216
rect 3240 18164 3292 18216
rect 7380 18232 7432 18284
rect 8208 18232 8260 18284
rect 9220 18232 9272 18284
rect 11612 18368 11664 18420
rect 11888 18411 11940 18420
rect 11888 18377 11897 18411
rect 11897 18377 11931 18411
rect 11931 18377 11940 18411
rect 11888 18368 11940 18377
rect 11980 18368 12032 18420
rect 16856 18368 16908 18420
rect 18236 18368 18288 18420
rect 19248 18368 19300 18420
rect 29644 18368 29696 18420
rect 32496 18411 32548 18420
rect 32496 18377 32505 18411
rect 32505 18377 32539 18411
rect 32539 18377 32548 18411
rect 32496 18368 32548 18377
rect 40592 18368 40644 18420
rect 11060 18300 11112 18352
rect 12716 18300 12768 18352
rect 4620 18164 4672 18216
rect 5540 18164 5592 18216
rect 6092 18164 6144 18216
rect 9588 18164 9640 18216
rect 10876 18232 10928 18284
rect 12348 18232 12400 18284
rect 12532 18232 12584 18284
rect 13176 18275 13228 18284
rect 13176 18241 13185 18275
rect 13185 18241 13219 18275
rect 13219 18241 13228 18275
rect 13176 18232 13228 18241
rect 13912 18300 13964 18352
rect 30564 18300 30616 18352
rect 31944 18300 31996 18352
rect 32772 18300 32824 18352
rect 33416 18300 33468 18352
rect 34428 18300 34480 18352
rect 37188 18300 37240 18352
rect 37556 18300 37608 18352
rect 39304 18300 39356 18352
rect 11428 18164 11480 18216
rect 13636 18232 13688 18284
rect 14280 18275 14332 18284
rect 14280 18241 14289 18275
rect 14289 18241 14323 18275
rect 14323 18241 14332 18275
rect 14280 18232 14332 18241
rect 14372 18275 14424 18284
rect 14372 18241 14382 18275
rect 14382 18241 14416 18275
rect 14416 18241 14424 18275
rect 14556 18275 14608 18284
rect 14372 18232 14424 18241
rect 14556 18241 14565 18275
rect 14565 18241 14599 18275
rect 14599 18241 14608 18275
rect 14556 18232 14608 18241
rect 14740 18275 14792 18284
rect 14740 18241 14754 18275
rect 14754 18241 14788 18275
rect 14788 18241 14792 18275
rect 14740 18232 14792 18241
rect 5816 18139 5868 18148
rect 5816 18105 5825 18139
rect 5825 18105 5859 18139
rect 5859 18105 5868 18139
rect 5816 18096 5868 18105
rect 1952 18028 2004 18080
rect 3332 18071 3384 18080
rect 3332 18037 3341 18071
rect 3341 18037 3375 18071
rect 3375 18037 3384 18071
rect 3332 18028 3384 18037
rect 6736 18071 6788 18080
rect 6736 18037 6745 18071
rect 6745 18037 6779 18071
rect 6779 18037 6788 18071
rect 6736 18028 6788 18037
rect 10876 18096 10928 18148
rect 16948 18164 17000 18216
rect 17960 18232 18012 18284
rect 18052 18164 18104 18216
rect 13912 18096 13964 18148
rect 19248 18232 19300 18284
rect 20628 18164 20680 18216
rect 19248 18096 19300 18148
rect 22100 18232 22152 18284
rect 23388 18275 23440 18284
rect 23388 18241 23397 18275
rect 23397 18241 23431 18275
rect 23431 18241 23440 18275
rect 23388 18232 23440 18241
rect 24492 18275 24544 18284
rect 24492 18241 24501 18275
rect 24501 18241 24535 18275
rect 24535 18241 24544 18275
rect 24492 18232 24544 18241
rect 24676 18275 24728 18284
rect 24676 18241 24685 18275
rect 24685 18241 24719 18275
rect 24719 18241 24728 18275
rect 24676 18232 24728 18241
rect 21916 18164 21968 18216
rect 24400 18164 24452 18216
rect 24952 18232 25004 18284
rect 25780 18232 25832 18284
rect 26976 18232 27028 18284
rect 29276 18232 29328 18284
rect 32220 18232 32272 18284
rect 26240 18164 26292 18216
rect 28816 18164 28868 18216
rect 31668 18164 31720 18216
rect 36452 18275 36504 18284
rect 36452 18241 36461 18275
rect 36461 18241 36495 18275
rect 36495 18241 36504 18275
rect 36452 18232 36504 18241
rect 37464 18232 37516 18284
rect 37004 18164 37056 18216
rect 41052 18275 41104 18284
rect 41052 18241 41061 18275
rect 41061 18241 41095 18275
rect 41095 18241 41104 18275
rect 41052 18232 41104 18241
rect 41236 18275 41288 18284
rect 41236 18241 41245 18275
rect 41245 18241 41279 18275
rect 41279 18241 41288 18275
rect 41236 18232 41288 18241
rect 41328 18164 41380 18216
rect 6920 18028 6972 18080
rect 7748 18028 7800 18080
rect 9220 18071 9272 18080
rect 9220 18037 9229 18071
rect 9229 18037 9263 18071
rect 9263 18037 9272 18071
rect 9220 18028 9272 18037
rect 10324 18071 10376 18080
rect 10324 18037 10333 18071
rect 10333 18037 10367 18071
rect 10367 18037 10376 18071
rect 10324 18028 10376 18037
rect 13820 18071 13872 18080
rect 13820 18037 13829 18071
rect 13829 18037 13863 18071
rect 13863 18037 13872 18071
rect 13820 18028 13872 18037
rect 14924 18028 14976 18080
rect 21916 18028 21968 18080
rect 23664 18096 23716 18148
rect 27160 18096 27212 18148
rect 24860 18028 24912 18080
rect 25044 18071 25096 18080
rect 25044 18037 25053 18071
rect 25053 18037 25087 18071
rect 25087 18037 25096 18071
rect 25044 18028 25096 18037
rect 29736 18071 29788 18080
rect 29736 18037 29745 18071
rect 29745 18037 29779 18071
rect 29779 18037 29788 18071
rect 29736 18028 29788 18037
rect 30012 18028 30064 18080
rect 32588 18028 32640 18080
rect 38936 18071 38988 18080
rect 38936 18037 38945 18071
rect 38945 18037 38979 18071
rect 38979 18037 38988 18071
rect 38936 18028 38988 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1676 17824 1728 17876
rect 4068 17824 4120 17876
rect 5816 17824 5868 17876
rect 6184 17824 6236 17876
rect 9864 17824 9916 17876
rect 12716 17824 12768 17876
rect 4896 17799 4948 17808
rect 4896 17765 4905 17799
rect 4905 17765 4939 17799
rect 4939 17765 4948 17799
rect 4896 17756 4948 17765
rect 5080 17756 5132 17808
rect 9220 17756 9272 17808
rect 12992 17756 13044 17808
rect 3332 17688 3384 17740
rect 2412 17663 2464 17672
rect 2412 17629 2421 17663
rect 2421 17629 2455 17663
rect 2455 17629 2464 17663
rect 2412 17620 2464 17629
rect 4712 17663 4764 17672
rect 4712 17629 4721 17663
rect 4721 17629 4755 17663
rect 4755 17629 4764 17663
rect 4712 17620 4764 17629
rect 5172 17620 5224 17672
rect 9680 17620 9732 17672
rect 10600 17663 10652 17672
rect 10600 17629 10609 17663
rect 10609 17629 10643 17663
rect 10643 17629 10652 17663
rect 10600 17620 10652 17629
rect 13636 17688 13688 17740
rect 16028 17688 16080 17740
rect 24860 17824 24912 17876
rect 25688 17824 25740 17876
rect 13268 17660 13320 17672
rect 13268 17626 13277 17660
rect 13277 17626 13311 17660
rect 13311 17626 13320 17660
rect 13452 17663 13504 17672
rect 13268 17620 13320 17626
rect 13452 17629 13461 17663
rect 13461 17629 13495 17663
rect 13495 17629 13504 17663
rect 13452 17620 13504 17629
rect 13820 17620 13872 17672
rect 19984 17620 20036 17672
rect 20260 17620 20312 17672
rect 23112 17620 23164 17672
rect 24400 17620 24452 17672
rect 25412 17620 25464 17672
rect 29368 17824 29420 17876
rect 30380 17824 30432 17876
rect 31944 17756 31996 17808
rect 32772 17756 32824 17808
rect 4896 17552 4948 17604
rect 12716 17552 12768 17604
rect 12072 17527 12124 17536
rect 12072 17493 12081 17527
rect 12081 17493 12115 17527
rect 12115 17493 12124 17527
rect 12072 17484 12124 17493
rect 12808 17527 12860 17536
rect 12808 17493 12817 17527
rect 12817 17493 12851 17527
rect 12851 17493 12860 17527
rect 12808 17484 12860 17493
rect 12992 17484 13044 17536
rect 14096 17484 14148 17536
rect 14372 17484 14424 17536
rect 20444 17484 20496 17536
rect 20904 17484 20956 17536
rect 21824 17552 21876 17604
rect 25688 17552 25740 17604
rect 29092 17620 29144 17672
rect 31300 17620 31352 17672
rect 31944 17663 31996 17672
rect 31944 17629 31953 17663
rect 31953 17629 31987 17663
rect 31987 17629 31996 17663
rect 31944 17620 31996 17629
rect 32404 17620 32456 17672
rect 37464 17867 37516 17876
rect 37464 17833 37473 17867
rect 37473 17833 37507 17867
rect 37507 17833 37516 17867
rect 37464 17824 37516 17833
rect 41236 17824 41288 17876
rect 35900 17688 35952 17740
rect 38200 17731 38252 17740
rect 38200 17697 38209 17731
rect 38209 17697 38243 17731
rect 38243 17697 38252 17731
rect 38200 17688 38252 17697
rect 41052 17688 41104 17740
rect 37924 17663 37976 17672
rect 37924 17629 37933 17663
rect 37933 17629 37967 17663
rect 37967 17629 37976 17663
rect 37924 17620 37976 17629
rect 22192 17484 22244 17536
rect 25504 17484 25556 17536
rect 27436 17552 27488 17604
rect 34060 17552 34112 17604
rect 36360 17595 36412 17604
rect 36360 17561 36394 17595
rect 36394 17561 36412 17595
rect 38936 17620 38988 17672
rect 36360 17552 36412 17561
rect 26148 17484 26200 17536
rect 33416 17527 33468 17536
rect 33416 17493 33425 17527
rect 33425 17493 33459 17527
rect 33459 17493 33468 17527
rect 33416 17484 33468 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 11428 17280 11480 17332
rect 13268 17280 13320 17332
rect 13912 17323 13964 17332
rect 13912 17289 13921 17323
rect 13921 17289 13955 17323
rect 13955 17289 13964 17323
rect 13912 17280 13964 17289
rect 14096 17280 14148 17332
rect 16856 17280 16908 17332
rect 21824 17323 21876 17332
rect 21824 17289 21833 17323
rect 21833 17289 21867 17323
rect 21867 17289 21876 17323
rect 21824 17280 21876 17289
rect 1860 17212 1912 17264
rect 2780 17212 2832 17264
rect 6552 17212 6604 17264
rect 12072 17212 12124 17264
rect 12348 17212 12400 17264
rect 4988 17144 5040 17196
rect 6000 17144 6052 17196
rect 9588 17187 9640 17196
rect 9588 17153 9597 17187
rect 9597 17153 9631 17187
rect 9631 17153 9640 17187
rect 9588 17144 9640 17153
rect 10324 17144 10376 17196
rect 11612 17144 11664 17196
rect 12532 17144 12584 17196
rect 14372 17144 14424 17196
rect 15200 17187 15252 17196
rect 15200 17153 15209 17187
rect 15209 17153 15243 17187
rect 15243 17153 15252 17187
rect 15200 17144 15252 17153
rect 15292 17144 15344 17196
rect 25504 17280 25556 17332
rect 25688 17323 25740 17332
rect 25688 17289 25697 17323
rect 25697 17289 25731 17323
rect 25731 17289 25740 17323
rect 25688 17280 25740 17289
rect 23388 17212 23440 17264
rect 26700 17280 26752 17332
rect 27252 17280 27304 17332
rect 29184 17280 29236 17332
rect 33508 17280 33560 17332
rect 34612 17280 34664 17332
rect 36360 17323 36412 17332
rect 26608 17212 26660 17264
rect 30656 17212 30708 17264
rect 34428 17212 34480 17264
rect 13268 17076 13320 17128
rect 14464 17076 14516 17128
rect 14924 17119 14976 17128
rect 14924 17085 14933 17119
rect 14933 17085 14967 17119
rect 14967 17085 14976 17119
rect 14924 17076 14976 17085
rect 16580 17076 16632 17128
rect 21916 17076 21968 17128
rect 11704 17008 11756 17060
rect 18144 17008 18196 17060
rect 5172 16983 5224 16992
rect 5172 16949 5181 16983
rect 5181 16949 5215 16983
rect 5215 16949 5224 16983
rect 5172 16940 5224 16949
rect 6000 16940 6052 16992
rect 10600 16940 10652 16992
rect 19340 16940 19392 16992
rect 21272 16983 21324 16992
rect 21272 16949 21281 16983
rect 21281 16949 21315 16983
rect 21315 16949 21324 16983
rect 22284 17190 22336 17196
rect 22284 17156 22293 17190
rect 22293 17156 22327 17190
rect 22327 17156 22336 17190
rect 22284 17144 22336 17156
rect 22560 17144 22612 17196
rect 23020 17119 23072 17128
rect 23020 17085 23029 17119
rect 23029 17085 23063 17119
rect 23063 17085 23072 17119
rect 23020 17076 23072 17085
rect 23664 17119 23716 17128
rect 23664 17085 23673 17119
rect 23673 17085 23707 17119
rect 23707 17085 23716 17119
rect 23664 17076 23716 17085
rect 24952 17076 25004 17128
rect 22284 17008 22336 17060
rect 22560 17008 22612 17060
rect 26148 17187 26200 17196
rect 26148 17153 26157 17187
rect 26157 17153 26191 17187
rect 26191 17153 26200 17187
rect 26148 17144 26200 17153
rect 25320 17008 25372 17060
rect 26148 17008 26200 17060
rect 26792 17144 26844 17196
rect 29828 17144 29880 17196
rect 30012 17187 30064 17196
rect 30012 17153 30021 17187
rect 30021 17153 30055 17187
rect 30055 17153 30064 17187
rect 30012 17144 30064 17153
rect 31392 17144 31444 17196
rect 32404 17144 32456 17196
rect 32588 17144 32640 17196
rect 32772 17187 32824 17196
rect 32772 17153 32781 17187
rect 32781 17153 32815 17187
rect 32815 17153 32824 17187
rect 32772 17144 32824 17153
rect 26976 17119 27028 17128
rect 26976 17085 26985 17119
rect 26985 17085 27019 17119
rect 27019 17085 27028 17119
rect 26976 17076 27028 17085
rect 28724 17076 28776 17128
rect 30932 17076 30984 17128
rect 31576 17076 31628 17128
rect 35624 17144 35676 17196
rect 33600 17119 33652 17128
rect 33600 17085 33609 17119
rect 33609 17085 33643 17119
rect 33643 17085 33652 17119
rect 33600 17076 33652 17085
rect 36084 17187 36136 17196
rect 36084 17153 36113 17187
rect 36113 17153 36136 17187
rect 36360 17289 36369 17323
rect 36369 17289 36403 17323
rect 36403 17289 36412 17323
rect 36360 17280 36412 17289
rect 37464 17255 37516 17264
rect 37464 17221 37473 17255
rect 37473 17221 37507 17255
rect 37507 17221 37516 17255
rect 37464 17212 37516 17221
rect 37924 17212 37976 17264
rect 36084 17144 36136 17153
rect 37556 17144 37608 17196
rect 38752 17187 38804 17196
rect 38752 17153 38761 17187
rect 38761 17153 38795 17187
rect 38795 17153 38804 17187
rect 38752 17144 38804 17153
rect 39856 17076 39908 17128
rect 58164 17051 58216 17060
rect 21272 16940 21324 16949
rect 25504 16940 25556 16992
rect 28356 16983 28408 16992
rect 28356 16949 28365 16983
rect 28365 16949 28399 16983
rect 28399 16949 28408 16983
rect 28356 16940 28408 16949
rect 29368 16940 29420 16992
rect 31576 16983 31628 16992
rect 31576 16949 31585 16983
rect 31585 16949 31619 16983
rect 31619 16949 31628 16983
rect 31576 16940 31628 16949
rect 58164 17017 58173 17051
rect 58173 17017 58207 17051
rect 58207 17017 58216 17051
rect 58164 17008 58216 17017
rect 33968 16940 34020 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 3240 16779 3292 16788
rect 3240 16745 3249 16779
rect 3249 16745 3283 16779
rect 3283 16745 3292 16779
rect 3240 16736 3292 16745
rect 4988 16779 5040 16788
rect 4988 16745 4997 16779
rect 4997 16745 5031 16779
rect 5031 16745 5040 16779
rect 4988 16736 5040 16745
rect 9680 16736 9732 16788
rect 4896 16668 4948 16720
rect 1860 16643 1912 16652
rect 1860 16609 1869 16643
rect 1869 16609 1903 16643
rect 1903 16609 1912 16643
rect 1860 16600 1912 16609
rect 9588 16600 9640 16652
rect 1952 16532 2004 16584
rect 6000 16532 6052 16584
rect 9404 16532 9456 16584
rect 22468 16736 22520 16788
rect 24860 16779 24912 16788
rect 24860 16745 24869 16779
rect 24869 16745 24903 16779
rect 24903 16745 24912 16779
rect 24860 16736 24912 16745
rect 25044 16779 25096 16788
rect 25044 16745 25053 16779
rect 25053 16745 25087 16779
rect 25087 16745 25096 16779
rect 25044 16736 25096 16745
rect 26792 16779 26844 16788
rect 26792 16745 26801 16779
rect 26801 16745 26835 16779
rect 26835 16745 26844 16779
rect 26792 16736 26844 16745
rect 27436 16779 27488 16788
rect 27436 16745 27445 16779
rect 27445 16745 27479 16779
rect 27479 16745 27488 16779
rect 27436 16736 27488 16745
rect 31300 16736 31352 16788
rect 34060 16736 34112 16788
rect 35624 16736 35676 16788
rect 36268 16779 36320 16788
rect 36268 16745 36277 16779
rect 36277 16745 36311 16779
rect 36311 16745 36320 16779
rect 36268 16736 36320 16745
rect 40684 16736 40736 16788
rect 9864 16668 9916 16720
rect 10232 16600 10284 16652
rect 12992 16668 13044 16720
rect 12716 16643 12768 16652
rect 12716 16609 12725 16643
rect 12725 16609 12759 16643
rect 12759 16609 12768 16643
rect 12716 16600 12768 16609
rect 20720 16668 20772 16720
rect 10968 16575 11020 16584
rect 10968 16541 10977 16575
rect 10977 16541 11011 16575
rect 11011 16541 11020 16575
rect 10968 16532 11020 16541
rect 11060 16575 11112 16584
rect 11060 16541 11070 16575
rect 11070 16541 11104 16575
rect 11104 16541 11112 16575
rect 11060 16532 11112 16541
rect 11704 16532 11756 16584
rect 7564 16464 7616 16516
rect 11244 16507 11296 16516
rect 11244 16473 11253 16507
rect 11253 16473 11287 16507
rect 11287 16473 11296 16507
rect 11244 16464 11296 16473
rect 13912 16464 13964 16516
rect 15844 16575 15896 16584
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 15844 16532 15896 16541
rect 16856 16575 16908 16584
rect 16856 16541 16865 16575
rect 16865 16541 16899 16575
rect 16899 16541 16908 16575
rect 16856 16532 16908 16541
rect 17132 16532 17184 16584
rect 18604 16600 18656 16652
rect 20260 16600 20312 16652
rect 22100 16600 22152 16652
rect 22744 16600 22796 16652
rect 22928 16600 22980 16652
rect 17316 16464 17368 16516
rect 17776 16575 17828 16584
rect 17776 16541 17785 16575
rect 17785 16541 17819 16575
rect 17819 16541 17828 16575
rect 17776 16532 17828 16541
rect 18144 16532 18196 16584
rect 23112 16575 23164 16584
rect 23112 16541 23121 16575
rect 23121 16541 23155 16575
rect 23155 16541 23164 16575
rect 23112 16532 23164 16541
rect 25044 16575 25096 16584
rect 25044 16541 25053 16575
rect 25053 16541 25087 16575
rect 25087 16541 25096 16575
rect 25044 16532 25096 16541
rect 25504 16532 25556 16584
rect 26148 16575 26200 16584
rect 26148 16541 26163 16575
rect 26163 16541 26197 16575
rect 26197 16541 26200 16575
rect 26332 16575 26384 16584
rect 26148 16532 26200 16541
rect 26332 16541 26341 16575
rect 26341 16541 26375 16575
rect 26375 16541 26384 16575
rect 26332 16532 26384 16541
rect 26700 16600 26752 16652
rect 27252 16600 27304 16652
rect 26608 16532 26660 16584
rect 27528 16532 27580 16584
rect 29552 16532 29604 16584
rect 26240 16464 26292 16516
rect 28356 16464 28408 16516
rect 28908 16464 28960 16516
rect 30104 16464 30156 16516
rect 32680 16532 32732 16584
rect 33600 16532 33652 16584
rect 37004 16575 37056 16584
rect 37004 16541 37013 16575
rect 37013 16541 37047 16575
rect 37047 16541 37056 16575
rect 37004 16532 37056 16541
rect 33416 16464 33468 16516
rect 37188 16507 37240 16516
rect 37188 16473 37197 16507
rect 37197 16473 37231 16507
rect 37231 16473 37240 16507
rect 37188 16464 37240 16473
rect 38660 16532 38712 16584
rect 40224 16532 40276 16584
rect 39212 16507 39264 16516
rect 39212 16473 39221 16507
rect 39221 16473 39255 16507
rect 39255 16473 39264 16507
rect 39856 16507 39908 16516
rect 39212 16464 39264 16473
rect 39856 16473 39865 16507
rect 39865 16473 39899 16507
rect 39899 16473 39908 16507
rect 39856 16464 39908 16473
rect 7380 16396 7432 16448
rect 10416 16439 10468 16448
rect 10416 16405 10425 16439
rect 10425 16405 10459 16439
rect 10459 16405 10468 16439
rect 10416 16396 10468 16405
rect 12716 16396 12768 16448
rect 15384 16439 15436 16448
rect 15384 16405 15393 16439
rect 15393 16405 15427 16439
rect 15427 16405 15436 16439
rect 15384 16396 15436 16405
rect 17132 16439 17184 16448
rect 17132 16405 17141 16439
rect 17141 16405 17175 16439
rect 17175 16405 17184 16439
rect 17132 16396 17184 16405
rect 18420 16396 18472 16448
rect 19432 16396 19484 16448
rect 30012 16396 30064 16448
rect 35900 16396 35952 16448
rect 36820 16439 36872 16448
rect 36820 16405 36829 16439
rect 36829 16405 36863 16439
rect 36863 16405 36872 16439
rect 36820 16396 36872 16405
rect 38200 16396 38252 16448
rect 40316 16396 40368 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 10140 16192 10192 16244
rect 11152 16192 11204 16244
rect 12164 16235 12216 16244
rect 12164 16201 12173 16235
rect 12173 16201 12207 16235
rect 12207 16201 12216 16235
rect 12164 16192 12216 16201
rect 12440 16192 12492 16244
rect 15844 16192 15896 16244
rect 17316 16192 17368 16244
rect 17776 16192 17828 16244
rect 20812 16192 20864 16244
rect 23112 16192 23164 16244
rect 23388 16192 23440 16244
rect 3792 16124 3844 16176
rect 2136 16056 2188 16108
rect 10416 16124 10468 16176
rect 4620 15988 4672 16040
rect 5356 15988 5408 16040
rect 2504 15852 2556 15904
rect 2596 15852 2648 15904
rect 6000 15852 6052 15904
rect 6552 15852 6604 15904
rect 8668 15852 8720 15904
rect 10232 16056 10284 16108
rect 11244 16124 11296 16176
rect 10968 16056 11020 16108
rect 11520 16099 11572 16108
rect 11520 16065 11529 16099
rect 11529 16065 11563 16099
rect 11563 16065 11572 16099
rect 11520 16056 11572 16065
rect 11612 16099 11664 16108
rect 11612 16065 11622 16099
rect 11622 16065 11656 16099
rect 11656 16065 11664 16099
rect 11612 16056 11664 16065
rect 13360 16124 13412 16176
rect 17960 16167 18012 16176
rect 17960 16133 17969 16167
rect 17969 16133 18003 16167
rect 18003 16133 18012 16167
rect 17960 16124 18012 16133
rect 11980 16099 12032 16108
rect 11980 16065 11994 16099
rect 11994 16065 12028 16099
rect 12028 16065 12032 16099
rect 11980 16056 12032 16065
rect 12716 16056 12768 16108
rect 12992 16056 13044 16108
rect 14280 16099 14332 16108
rect 14280 16065 14289 16099
rect 14289 16065 14323 16099
rect 14323 16065 14332 16099
rect 14280 16056 14332 16065
rect 14924 16056 14976 16108
rect 16856 16056 16908 16108
rect 12900 15988 12952 16040
rect 14556 16031 14608 16040
rect 14556 15997 14565 16031
rect 14565 15997 14599 16031
rect 14599 15997 14608 16031
rect 14556 15988 14608 15997
rect 19432 16056 19484 16108
rect 18236 15988 18288 16040
rect 12716 15920 12768 15972
rect 19892 15920 19944 15972
rect 20812 16099 20864 16108
rect 20812 16065 20821 16099
rect 20821 16065 20855 16099
rect 20855 16065 20864 16099
rect 20812 16056 20864 16065
rect 22100 16056 22152 16108
rect 23480 16124 23532 16176
rect 25504 16192 25556 16244
rect 26332 16192 26384 16244
rect 26608 16192 26660 16244
rect 28908 16235 28960 16244
rect 26240 16167 26292 16176
rect 13820 15895 13872 15904
rect 13820 15861 13829 15895
rect 13829 15861 13863 15895
rect 13863 15861 13872 15895
rect 13820 15852 13872 15861
rect 20352 15852 20404 15904
rect 23664 16056 23716 16108
rect 26240 16133 26249 16167
rect 26249 16133 26283 16167
rect 26283 16133 26292 16167
rect 26240 16124 26292 16133
rect 27436 16124 27488 16176
rect 28908 16201 28917 16235
rect 28917 16201 28951 16235
rect 28951 16201 28960 16235
rect 28908 16192 28960 16201
rect 33600 16192 33652 16244
rect 40224 16235 40276 16244
rect 40224 16201 40233 16235
rect 40233 16201 40267 16235
rect 40267 16201 40276 16235
rect 40224 16192 40276 16201
rect 38292 16124 38344 16176
rect 26608 16056 26660 16108
rect 23572 15988 23624 16040
rect 27528 15988 27580 16040
rect 27252 15895 27304 15904
rect 27252 15861 27261 15895
rect 27261 15861 27295 15895
rect 27295 15861 27304 15895
rect 27252 15852 27304 15861
rect 27896 15852 27948 15904
rect 29368 16099 29420 16108
rect 29368 16065 29377 16099
rect 29377 16065 29411 16099
rect 29411 16065 29420 16099
rect 29368 16056 29420 16065
rect 30196 16056 30248 16108
rect 31300 16099 31352 16108
rect 31300 16065 31309 16099
rect 31309 16065 31343 16099
rect 31343 16065 31352 16099
rect 31300 16056 31352 16065
rect 32496 16099 32548 16108
rect 32496 16065 32505 16099
rect 32505 16065 32539 16099
rect 32539 16065 32548 16099
rect 32496 16056 32548 16065
rect 37188 16056 37240 16108
rect 39304 16124 39356 16176
rect 39856 16056 39908 16108
rect 41144 16056 41196 16108
rect 30012 16031 30064 16040
rect 30012 15997 30021 16031
rect 30021 15997 30055 16031
rect 30055 15997 30064 16031
rect 30012 15988 30064 15997
rect 30104 15988 30156 16040
rect 35348 15988 35400 16040
rect 40684 16031 40736 16040
rect 40684 15997 40693 16031
rect 40693 15997 40727 16031
rect 40727 15997 40736 16031
rect 40684 15988 40736 15997
rect 31392 15852 31444 15904
rect 58164 15895 58216 15904
rect 58164 15861 58173 15895
rect 58173 15861 58207 15895
rect 58207 15861 58216 15895
rect 58164 15852 58216 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2136 15691 2188 15700
rect 2136 15657 2145 15691
rect 2145 15657 2179 15691
rect 2179 15657 2188 15691
rect 2136 15648 2188 15657
rect 7564 15691 7616 15700
rect 7564 15657 7573 15691
rect 7573 15657 7607 15691
rect 7607 15657 7616 15691
rect 7564 15648 7616 15657
rect 8484 15648 8536 15700
rect 10232 15691 10284 15700
rect 10232 15657 10241 15691
rect 10241 15657 10275 15691
rect 10275 15657 10284 15691
rect 10232 15648 10284 15657
rect 12532 15648 12584 15700
rect 14280 15691 14332 15700
rect 14280 15657 14289 15691
rect 14289 15657 14323 15691
rect 14323 15657 14332 15691
rect 14280 15648 14332 15657
rect 2596 15512 2648 15564
rect 2780 15512 2832 15564
rect 7288 15512 7340 15564
rect 2412 15487 2464 15496
rect 2412 15453 2421 15487
rect 2421 15453 2455 15487
rect 2455 15453 2464 15487
rect 2412 15444 2464 15453
rect 4252 15376 4304 15428
rect 3792 15308 3844 15360
rect 6092 15487 6144 15496
rect 6092 15453 6101 15487
rect 6101 15453 6135 15487
rect 6135 15453 6144 15487
rect 6092 15444 6144 15453
rect 6644 15444 6696 15496
rect 7012 15487 7064 15496
rect 6552 15376 6604 15428
rect 7012 15453 7021 15487
rect 7021 15453 7055 15487
rect 7055 15453 7064 15487
rect 7012 15444 7064 15453
rect 7380 15487 7432 15496
rect 7380 15453 7389 15487
rect 7389 15453 7423 15487
rect 7423 15453 7432 15487
rect 7380 15444 7432 15453
rect 8300 15487 8352 15496
rect 8300 15453 8309 15487
rect 8309 15453 8343 15487
rect 8343 15453 8352 15487
rect 8300 15444 8352 15453
rect 9864 15444 9916 15496
rect 10876 15444 10928 15496
rect 12072 15444 12124 15496
rect 13636 15444 13688 15496
rect 12808 15376 12860 15428
rect 5080 15308 5132 15360
rect 5632 15351 5684 15360
rect 5632 15317 5641 15351
rect 5641 15317 5675 15351
rect 5675 15317 5684 15351
rect 5632 15308 5684 15317
rect 6828 15308 6880 15360
rect 10968 15351 11020 15360
rect 10968 15317 10977 15351
rect 10977 15317 11011 15351
rect 11011 15317 11020 15351
rect 10968 15308 11020 15317
rect 12992 15308 13044 15360
rect 13820 15512 13872 15564
rect 14004 15444 14056 15496
rect 15108 15487 15160 15496
rect 15108 15453 15117 15487
rect 15117 15453 15151 15487
rect 15151 15453 15160 15487
rect 15108 15444 15160 15453
rect 15384 15487 15436 15496
rect 15384 15453 15418 15487
rect 15418 15453 15436 15487
rect 15384 15444 15436 15453
rect 19340 15648 19392 15700
rect 19892 15691 19944 15700
rect 19892 15657 19901 15691
rect 19901 15657 19935 15691
rect 19935 15657 19944 15691
rect 19892 15648 19944 15657
rect 22100 15691 22152 15700
rect 22100 15657 22109 15691
rect 22109 15657 22143 15691
rect 22143 15657 22152 15691
rect 22100 15648 22152 15657
rect 23664 15648 23716 15700
rect 26700 15648 26752 15700
rect 29920 15648 29972 15700
rect 31208 15648 31260 15700
rect 38292 15691 38344 15700
rect 38292 15657 38301 15691
rect 38301 15657 38335 15691
rect 38335 15657 38344 15691
rect 38292 15648 38344 15657
rect 39856 15691 39908 15700
rect 39856 15657 39865 15691
rect 39865 15657 39899 15691
rect 39899 15657 39908 15691
rect 39856 15648 39908 15657
rect 18696 15555 18748 15564
rect 18696 15521 18705 15555
rect 18705 15521 18739 15555
rect 18739 15521 18748 15555
rect 18696 15512 18748 15521
rect 19524 15512 19576 15564
rect 16028 15376 16080 15428
rect 19340 15444 19392 15496
rect 27068 15580 27120 15632
rect 20260 15512 20312 15564
rect 34704 15512 34756 15564
rect 37004 15512 37056 15564
rect 39212 15512 39264 15564
rect 20812 15444 20864 15496
rect 21640 15444 21692 15496
rect 22100 15376 22152 15428
rect 22192 15376 22244 15428
rect 27068 15444 27120 15496
rect 27528 15487 27580 15496
rect 23848 15376 23900 15428
rect 27528 15453 27537 15487
rect 27537 15453 27571 15487
rect 27571 15453 27580 15487
rect 27528 15444 27580 15453
rect 29552 15487 29604 15496
rect 29552 15453 29561 15487
rect 29561 15453 29595 15487
rect 29595 15453 29604 15487
rect 29552 15444 29604 15453
rect 31208 15444 31260 15496
rect 33048 15444 33100 15496
rect 16856 15308 16908 15360
rect 19524 15308 19576 15360
rect 21180 15308 21232 15360
rect 29644 15376 29696 15428
rect 31392 15419 31444 15428
rect 31392 15385 31401 15419
rect 31401 15385 31435 15419
rect 31435 15385 31444 15419
rect 31392 15376 31444 15385
rect 33600 15444 33652 15496
rect 37740 15444 37792 15496
rect 37924 15444 37976 15496
rect 38292 15444 38344 15496
rect 38660 15376 38712 15428
rect 40316 15487 40368 15496
rect 40316 15453 40325 15487
rect 40325 15453 40359 15487
rect 40359 15453 40368 15487
rect 40316 15444 40368 15453
rect 41144 15444 41196 15496
rect 30012 15308 30064 15360
rect 30196 15308 30248 15360
rect 30472 15308 30524 15360
rect 31760 15351 31812 15360
rect 31760 15317 31769 15351
rect 31769 15317 31803 15351
rect 31803 15317 31812 15351
rect 31760 15308 31812 15317
rect 32496 15308 32548 15360
rect 37924 15308 37976 15360
rect 38752 15308 38804 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 3792 15147 3844 15156
rect 3792 15113 3801 15147
rect 3801 15113 3835 15147
rect 3835 15113 3844 15147
rect 3792 15104 3844 15113
rect 4252 15147 4304 15156
rect 4252 15113 4261 15147
rect 4261 15113 4295 15147
rect 4295 15113 4304 15147
rect 4252 15104 4304 15113
rect 7012 15147 7064 15156
rect 7012 15113 7021 15147
rect 7021 15113 7055 15147
rect 7055 15113 7064 15147
rect 7012 15104 7064 15113
rect 8300 15104 8352 15156
rect 17224 15147 17276 15156
rect 2780 15036 2832 15088
rect 3240 15036 3292 15088
rect 6736 15036 6788 15088
rect 9496 15079 9548 15088
rect 9496 15045 9505 15079
rect 9505 15045 9539 15079
rect 9539 15045 9548 15079
rect 9496 15036 9548 15045
rect 12532 15036 12584 15088
rect 2504 14968 2556 15020
rect 4712 14968 4764 15020
rect 9588 15011 9640 15020
rect 2412 14764 2464 14816
rect 5908 14764 5960 14816
rect 9588 14977 9597 15011
rect 9597 14977 9631 15011
rect 9631 14977 9640 15011
rect 9588 14968 9640 14977
rect 12164 14968 12216 15020
rect 12624 15011 12676 15020
rect 12624 14977 12633 15011
rect 12633 14977 12667 15011
rect 12667 14977 12676 15011
rect 12624 14968 12676 14977
rect 12808 15036 12860 15088
rect 14004 15036 14056 15088
rect 17224 15113 17233 15147
rect 17233 15113 17267 15147
rect 17267 15113 17276 15147
rect 17224 15104 17276 15113
rect 18696 15036 18748 15088
rect 9772 14900 9824 14952
rect 11336 14900 11388 14952
rect 11704 14900 11756 14952
rect 13912 14968 13964 15020
rect 14648 14900 14700 14952
rect 17316 15011 17368 15020
rect 17316 14977 17325 15011
rect 17325 14977 17359 15011
rect 17359 14977 17368 15011
rect 18328 15011 18380 15020
rect 17316 14968 17368 14977
rect 18328 14977 18337 15011
rect 18337 14977 18371 15011
rect 18371 14977 18380 15011
rect 18328 14968 18380 14977
rect 18420 14968 18472 15020
rect 19432 15104 19484 15156
rect 20904 15104 20956 15156
rect 21180 15147 21232 15156
rect 21180 15113 21189 15147
rect 21189 15113 21223 15147
rect 21223 15113 21232 15147
rect 21180 15104 21232 15113
rect 29644 15147 29696 15156
rect 29644 15113 29653 15147
rect 29653 15113 29687 15147
rect 29687 15113 29696 15147
rect 29644 15104 29696 15113
rect 29920 15104 29972 15156
rect 8760 14764 8812 14816
rect 8852 14807 8904 14816
rect 8852 14773 8861 14807
rect 8861 14773 8895 14807
rect 8895 14773 8904 14807
rect 8852 14764 8904 14773
rect 9588 14764 9640 14816
rect 10048 14807 10100 14816
rect 10048 14773 10057 14807
rect 10057 14773 10091 14807
rect 10091 14773 10100 14807
rect 10048 14764 10100 14773
rect 10508 14764 10560 14816
rect 13912 14807 13964 14816
rect 13912 14773 13921 14807
rect 13921 14773 13955 14807
rect 13955 14773 13964 14807
rect 13912 14764 13964 14773
rect 15200 14764 15252 14816
rect 16028 14807 16080 14816
rect 16028 14773 16037 14807
rect 16037 14773 16071 14807
rect 16071 14773 16080 14807
rect 16028 14764 16080 14773
rect 16304 14764 16356 14816
rect 17316 14764 17368 14816
rect 19892 14900 19944 14952
rect 20628 14968 20680 15020
rect 21180 14968 21232 15020
rect 22100 14968 22152 15020
rect 22744 15036 22796 15088
rect 23480 14968 23532 15020
rect 23848 15011 23900 15020
rect 23572 14900 23624 14952
rect 23848 14977 23857 15011
rect 23857 14977 23891 15011
rect 23891 14977 23900 15011
rect 23848 14968 23900 14977
rect 25044 14968 25096 15020
rect 28632 14968 28684 15020
rect 29092 14968 29144 15020
rect 31760 15036 31812 15088
rect 37740 15104 37792 15156
rect 38568 15104 38620 15156
rect 38660 15104 38712 15156
rect 24400 14900 24452 14952
rect 27068 14900 27120 14952
rect 22192 14875 22244 14884
rect 19432 14764 19484 14816
rect 20260 14764 20312 14816
rect 22192 14841 22201 14875
rect 22201 14841 22235 14875
rect 22235 14841 22244 14875
rect 22192 14832 22244 14841
rect 23112 14764 23164 14816
rect 23572 14764 23624 14816
rect 23848 14807 23900 14816
rect 23848 14773 23857 14807
rect 23857 14773 23891 14807
rect 23891 14773 23900 14807
rect 23848 14764 23900 14773
rect 27344 14764 27396 14816
rect 27712 14764 27764 14816
rect 29092 14807 29144 14816
rect 29092 14773 29101 14807
rect 29101 14773 29135 14807
rect 29135 14773 29144 14807
rect 29092 14764 29144 14773
rect 30472 14968 30524 15020
rect 32404 14968 32456 15020
rect 33600 15011 33652 15020
rect 33600 14977 33609 15011
rect 33609 14977 33643 15011
rect 33643 14977 33652 15011
rect 33600 14968 33652 14977
rect 35440 14968 35492 15020
rect 36268 14968 36320 15020
rect 37924 15011 37976 15020
rect 37924 14977 37928 15011
rect 37928 14977 37962 15011
rect 37962 14977 37976 15011
rect 37924 14968 37976 14977
rect 35348 14943 35400 14952
rect 35348 14909 35357 14943
rect 35357 14909 35391 14943
rect 35391 14909 35400 14943
rect 35348 14900 35400 14909
rect 35808 14943 35860 14952
rect 35808 14909 35817 14943
rect 35817 14909 35851 14943
rect 35851 14909 35860 14943
rect 35808 14900 35860 14909
rect 37556 14900 37608 14952
rect 38292 14968 38344 15020
rect 38568 14968 38620 15020
rect 38752 14968 38804 15020
rect 41328 15036 41380 15088
rect 40316 14968 40368 15020
rect 40684 14968 40736 15020
rect 38660 14900 38712 14952
rect 30104 14764 30156 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 4712 14560 4764 14612
rect 7380 14560 7432 14612
rect 10048 14560 10100 14612
rect 4988 14492 5040 14544
rect 5080 14467 5132 14476
rect 5080 14433 5089 14467
rect 5089 14433 5123 14467
rect 5123 14433 5132 14467
rect 5080 14424 5132 14433
rect 9404 14492 9456 14544
rect 9588 14492 9640 14544
rect 14924 14560 14976 14612
rect 6644 14356 6696 14408
rect 7656 14399 7708 14408
rect 7656 14365 7665 14399
rect 7665 14365 7699 14399
rect 7699 14365 7708 14399
rect 7656 14356 7708 14365
rect 8208 14399 8260 14408
rect 8208 14365 8217 14399
rect 8217 14365 8251 14399
rect 8251 14365 8260 14399
rect 8208 14356 8260 14365
rect 11980 14356 12032 14408
rect 9588 14288 9640 14340
rect 9772 14331 9824 14340
rect 9772 14297 9781 14331
rect 9781 14297 9815 14331
rect 9815 14297 9824 14331
rect 9772 14288 9824 14297
rect 10140 14288 10192 14340
rect 20352 14560 20404 14612
rect 21088 14560 21140 14612
rect 22284 14560 22336 14612
rect 18236 14535 18288 14544
rect 18236 14501 18245 14535
rect 18245 14501 18279 14535
rect 18279 14501 18288 14535
rect 18236 14492 18288 14501
rect 20536 14424 20588 14476
rect 20628 14424 20680 14476
rect 15108 14356 15160 14408
rect 18328 14356 18380 14408
rect 19432 14356 19484 14408
rect 20076 14356 20128 14408
rect 15936 14288 15988 14340
rect 17132 14331 17184 14340
rect 5540 14220 5592 14272
rect 5632 14220 5684 14272
rect 7472 14263 7524 14272
rect 7472 14229 7481 14263
rect 7481 14229 7515 14263
rect 7515 14229 7524 14263
rect 7472 14220 7524 14229
rect 15292 14220 15344 14272
rect 15844 14220 15896 14272
rect 16304 14263 16356 14272
rect 16304 14229 16313 14263
rect 16313 14229 16347 14263
rect 16347 14229 16356 14263
rect 16304 14220 16356 14229
rect 17132 14297 17166 14331
rect 17166 14297 17184 14331
rect 17132 14288 17184 14297
rect 19892 14288 19944 14340
rect 21732 14399 21784 14408
rect 21732 14365 21741 14399
rect 21741 14365 21775 14399
rect 21775 14365 21784 14399
rect 21732 14356 21784 14365
rect 21916 14399 21968 14408
rect 21916 14365 21925 14399
rect 21925 14365 21959 14399
rect 21959 14365 21968 14399
rect 22744 14492 22796 14544
rect 23848 14560 23900 14612
rect 24400 14492 24452 14544
rect 24584 14492 24636 14544
rect 25044 14535 25096 14544
rect 25044 14501 25053 14535
rect 25053 14501 25087 14535
rect 25087 14501 25096 14535
rect 25044 14492 25096 14501
rect 37556 14560 37608 14612
rect 34704 14492 34756 14544
rect 34796 14492 34848 14544
rect 35348 14492 35400 14544
rect 28264 14424 28316 14476
rect 35808 14424 35860 14476
rect 21916 14356 21968 14365
rect 23480 14356 23532 14408
rect 25412 14356 25464 14408
rect 28632 14356 28684 14408
rect 31392 14356 31444 14408
rect 34704 14399 34756 14408
rect 19340 14220 19392 14272
rect 20076 14220 20128 14272
rect 20628 14220 20680 14272
rect 23664 14220 23716 14272
rect 23848 14263 23900 14272
rect 23848 14229 23857 14263
rect 23857 14229 23891 14263
rect 23891 14229 23900 14263
rect 23848 14220 23900 14229
rect 26976 14288 27028 14340
rect 27160 14331 27212 14340
rect 27160 14297 27194 14331
rect 27194 14297 27212 14331
rect 27160 14288 27212 14297
rect 29644 14288 29696 14340
rect 34704 14365 34713 14399
rect 34713 14365 34747 14399
rect 34747 14365 34756 14399
rect 34704 14356 34756 14365
rect 35532 14356 35584 14408
rect 37280 14492 37332 14544
rect 35440 14288 35492 14340
rect 37464 14356 37516 14408
rect 37740 14356 37792 14408
rect 38384 14399 38436 14408
rect 38384 14365 38393 14399
rect 38393 14365 38427 14399
rect 38427 14365 38436 14399
rect 38384 14356 38436 14365
rect 58164 14399 58216 14408
rect 58164 14365 58173 14399
rect 58173 14365 58207 14399
rect 58207 14365 58216 14399
rect 58164 14356 58216 14365
rect 39028 14331 39080 14340
rect 39028 14297 39037 14331
rect 39037 14297 39071 14331
rect 39071 14297 39080 14331
rect 39028 14288 39080 14297
rect 40316 14331 40368 14340
rect 40316 14297 40325 14331
rect 40325 14297 40359 14331
rect 40359 14297 40368 14331
rect 40316 14288 40368 14297
rect 28448 14220 28500 14272
rect 29828 14220 29880 14272
rect 36728 14220 36780 14272
rect 38568 14263 38620 14272
rect 38568 14229 38577 14263
rect 38577 14229 38611 14263
rect 38611 14229 38620 14263
rect 38568 14220 38620 14229
rect 40408 14263 40460 14272
rect 40408 14229 40417 14263
rect 40417 14229 40451 14263
rect 40451 14229 40460 14263
rect 40408 14220 40460 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 7656 14016 7708 14068
rect 9772 14016 9824 14068
rect 14004 14016 14056 14068
rect 16856 14016 16908 14068
rect 7472 13948 7524 14000
rect 7564 13948 7616 14000
rect 14924 13948 14976 14000
rect 19340 13948 19392 14000
rect 19432 13948 19484 14000
rect 20536 13991 20588 14000
rect 20536 13957 20545 13991
rect 20545 13957 20579 13991
rect 20579 13957 20588 13991
rect 20536 13948 20588 13957
rect 21916 14016 21968 14068
rect 22744 14016 22796 14068
rect 23112 14016 23164 14068
rect 25412 14016 25464 14068
rect 27160 14059 27212 14068
rect 27160 14025 27169 14059
rect 27169 14025 27203 14059
rect 27203 14025 27212 14059
rect 27160 14016 27212 14025
rect 10048 13880 10100 13932
rect 10876 13923 10928 13932
rect 10876 13889 10885 13923
rect 10885 13889 10919 13923
rect 10919 13889 10928 13923
rect 10876 13880 10928 13889
rect 11980 13923 12032 13932
rect 11980 13889 11989 13923
rect 11989 13889 12023 13923
rect 12023 13889 12032 13923
rect 11980 13880 12032 13889
rect 12164 13923 12216 13932
rect 12164 13889 12173 13923
rect 12173 13889 12207 13923
rect 12207 13889 12216 13923
rect 12164 13880 12216 13889
rect 14280 13923 14332 13932
rect 14280 13889 14298 13923
rect 14298 13889 14332 13923
rect 14280 13880 14332 13889
rect 15108 13880 15160 13932
rect 16304 13880 16356 13932
rect 22100 13880 22152 13932
rect 29644 14016 29696 14068
rect 30012 14016 30064 14068
rect 34796 14016 34848 14068
rect 23480 13880 23532 13932
rect 5540 13855 5592 13864
rect 5540 13821 5549 13855
rect 5549 13821 5583 13855
rect 5583 13821 5592 13855
rect 5540 13812 5592 13821
rect 7104 13855 7156 13864
rect 7104 13821 7113 13855
rect 7113 13821 7147 13855
rect 7147 13821 7156 13855
rect 7104 13812 7156 13821
rect 14648 13812 14700 13864
rect 21732 13812 21784 13864
rect 8760 13744 8812 13796
rect 9864 13744 9916 13796
rect 17592 13744 17644 13796
rect 17776 13744 17828 13796
rect 23756 13855 23808 13864
rect 23756 13821 23765 13855
rect 23765 13821 23799 13855
rect 23799 13821 23808 13855
rect 23756 13812 23808 13821
rect 25964 13880 26016 13932
rect 27068 13880 27120 13932
rect 27528 13923 27580 13932
rect 27528 13889 27552 13923
rect 27552 13889 27580 13923
rect 27528 13880 27580 13889
rect 28448 13991 28500 14000
rect 28448 13957 28457 13991
rect 28457 13957 28491 13991
rect 28491 13957 28500 13991
rect 28448 13948 28500 13957
rect 28632 13991 28684 14000
rect 28632 13957 28641 13991
rect 28641 13957 28675 13991
rect 28675 13957 28684 13991
rect 28632 13948 28684 13957
rect 28080 13880 28132 13932
rect 29092 13923 29144 13932
rect 29092 13889 29101 13923
rect 29101 13889 29135 13923
rect 29135 13889 29144 13923
rect 29092 13880 29144 13889
rect 30196 13948 30248 14000
rect 36452 13948 36504 14000
rect 37648 13991 37700 14000
rect 37648 13957 37657 13991
rect 37657 13957 37691 13991
rect 37691 13957 37700 13991
rect 37648 13948 37700 13957
rect 29828 13923 29880 13932
rect 29828 13889 29837 13923
rect 29837 13889 29871 13923
rect 29871 13889 29880 13923
rect 29828 13880 29880 13889
rect 24584 13812 24636 13864
rect 30104 13812 30156 13864
rect 23848 13744 23900 13796
rect 24308 13744 24360 13796
rect 29092 13744 29144 13796
rect 36268 13880 36320 13932
rect 36728 13923 36780 13932
rect 36728 13889 36737 13923
rect 36737 13889 36771 13923
rect 36771 13889 36780 13923
rect 36728 13880 36780 13889
rect 37464 13880 37516 13932
rect 38200 13880 38252 13932
rect 30748 13812 30800 13864
rect 33600 13812 33652 13864
rect 40316 13812 40368 13864
rect 9496 13719 9548 13728
rect 9496 13685 9505 13719
rect 9505 13685 9539 13719
rect 9539 13685 9548 13719
rect 9496 13676 9548 13685
rect 23204 13676 23256 13728
rect 23572 13719 23624 13728
rect 23572 13685 23581 13719
rect 23581 13685 23615 13719
rect 23615 13685 23624 13719
rect 23572 13676 23624 13685
rect 23940 13676 23992 13728
rect 27804 13676 27856 13728
rect 29276 13676 29328 13728
rect 30840 13676 30892 13728
rect 36084 13676 36136 13728
rect 38660 13676 38712 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 2412 13472 2464 13524
rect 4620 13472 4672 13524
rect 9588 13472 9640 13524
rect 9404 13404 9456 13456
rect 6644 13336 6696 13388
rect 10048 13472 10100 13524
rect 10600 13472 10652 13524
rect 17776 13472 17828 13524
rect 20536 13515 20588 13524
rect 20536 13481 20545 13515
rect 20545 13481 20579 13515
rect 20579 13481 20588 13515
rect 20536 13472 20588 13481
rect 23204 13515 23256 13524
rect 23204 13481 23213 13515
rect 23213 13481 23247 13515
rect 23247 13481 23256 13515
rect 23204 13472 23256 13481
rect 23664 13472 23716 13524
rect 25964 13515 26016 13524
rect 25964 13481 25973 13515
rect 25973 13481 26007 13515
rect 26007 13481 26016 13515
rect 25964 13472 26016 13481
rect 32496 13472 32548 13524
rect 37648 13515 37700 13524
rect 37648 13481 37657 13515
rect 37657 13481 37691 13515
rect 37691 13481 37700 13515
rect 37648 13472 37700 13481
rect 9864 13404 9916 13456
rect 26976 13447 27028 13456
rect 11336 13336 11388 13388
rect 26976 13413 26985 13447
rect 26985 13413 27019 13447
rect 27019 13413 27028 13447
rect 26976 13404 27028 13413
rect 3884 13268 3936 13320
rect 5080 13268 5132 13320
rect 8208 13268 8260 13320
rect 9864 13268 9916 13320
rect 14004 13268 14056 13320
rect 10600 13200 10652 13252
rect 14096 13243 14148 13252
rect 14096 13209 14105 13243
rect 14105 13209 14139 13243
rect 14139 13209 14148 13243
rect 19432 13268 19484 13320
rect 23204 13311 23256 13320
rect 23204 13277 23213 13311
rect 23213 13277 23247 13311
rect 23247 13277 23256 13311
rect 23204 13268 23256 13277
rect 24216 13268 24268 13320
rect 24584 13268 24636 13320
rect 14096 13200 14148 13209
rect 17868 13243 17920 13252
rect 17868 13209 17877 13243
rect 17877 13209 17911 13243
rect 17911 13209 17920 13243
rect 17868 13200 17920 13209
rect 6368 13175 6420 13184
rect 6368 13141 6377 13175
rect 6377 13141 6411 13175
rect 6411 13141 6420 13175
rect 6368 13132 6420 13141
rect 6920 13132 6972 13184
rect 7472 13175 7524 13184
rect 7472 13141 7481 13175
rect 7481 13141 7515 13175
rect 7515 13141 7524 13175
rect 7472 13132 7524 13141
rect 9036 13132 9088 13184
rect 9496 13132 9548 13184
rect 9864 13132 9916 13184
rect 14648 13132 14700 13184
rect 17776 13132 17828 13184
rect 22100 13200 22152 13252
rect 23388 13200 23440 13252
rect 23940 13200 23992 13252
rect 18512 13132 18564 13184
rect 23112 13132 23164 13184
rect 25228 13268 25280 13320
rect 27528 13404 27580 13456
rect 29644 13447 29696 13456
rect 29644 13413 29653 13447
rect 29653 13413 29687 13447
rect 29687 13413 29696 13447
rect 29644 13404 29696 13413
rect 27436 13308 27488 13320
rect 27436 13274 27445 13308
rect 27445 13274 27479 13308
rect 27479 13274 27488 13308
rect 27436 13268 27488 13274
rect 27804 13268 27856 13320
rect 28080 13268 28132 13320
rect 29920 13336 29972 13388
rect 29552 13268 29604 13320
rect 24860 13132 24912 13184
rect 29368 13200 29420 13252
rect 30104 13200 30156 13252
rect 30748 13243 30800 13252
rect 30748 13209 30766 13243
rect 30766 13209 30800 13243
rect 31944 13243 31996 13252
rect 30748 13200 30800 13209
rect 31944 13209 31953 13243
rect 31953 13209 31987 13243
rect 31987 13209 31996 13243
rect 31944 13200 31996 13209
rect 32128 13243 32180 13252
rect 32128 13209 32137 13243
rect 32137 13209 32171 13243
rect 32171 13209 32180 13243
rect 32128 13200 32180 13209
rect 29184 13132 29236 13184
rect 29552 13132 29604 13184
rect 32404 13132 32456 13184
rect 32956 13200 33008 13252
rect 35348 13268 35400 13320
rect 40408 13404 40460 13456
rect 35532 13200 35584 13252
rect 35624 13200 35676 13252
rect 35256 13175 35308 13184
rect 35256 13141 35265 13175
rect 35265 13141 35299 13175
rect 35299 13141 35308 13175
rect 35256 13132 35308 13141
rect 36452 13132 36504 13184
rect 38568 13311 38620 13320
rect 38568 13277 38577 13311
rect 38577 13277 38611 13311
rect 38611 13277 38620 13311
rect 38568 13268 38620 13277
rect 38844 13336 38896 13388
rect 39028 13336 39080 13388
rect 38752 13311 38804 13320
rect 38752 13277 38761 13311
rect 38761 13277 38795 13311
rect 38795 13277 38804 13311
rect 38752 13268 38804 13277
rect 58164 13311 58216 13320
rect 58164 13277 58173 13311
rect 58173 13277 58207 13311
rect 58207 13277 58216 13311
rect 58164 13268 58216 13277
rect 38660 13132 38712 13184
rect 39028 13175 39080 13184
rect 39028 13141 39037 13175
rect 39037 13141 39071 13175
rect 39071 13141 39080 13175
rect 39028 13132 39080 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 5080 12971 5132 12980
rect 5080 12937 5089 12971
rect 5089 12937 5123 12971
rect 5123 12937 5132 12971
rect 5080 12928 5132 12937
rect 14280 12928 14332 12980
rect 15752 12928 15804 12980
rect 17868 12928 17920 12980
rect 6552 12860 6604 12912
rect 3792 12792 3844 12844
rect 4620 12792 4672 12844
rect 4804 12792 4856 12844
rect 7472 12860 7524 12912
rect 6828 12835 6880 12844
rect 6828 12801 6837 12835
rect 6837 12801 6871 12835
rect 6871 12801 6880 12835
rect 6828 12792 6880 12801
rect 6920 12835 6972 12844
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 7196 12835 7248 12844
rect 6920 12792 6972 12801
rect 7196 12801 7205 12835
rect 7205 12801 7239 12835
rect 7239 12801 7248 12835
rect 7196 12792 7248 12801
rect 8208 12792 8260 12844
rect 12164 12792 12216 12844
rect 2412 12724 2464 12776
rect 2780 12767 2832 12776
rect 2780 12733 2789 12767
rect 2789 12733 2823 12767
rect 2823 12733 2832 12767
rect 2780 12724 2832 12733
rect 5356 12724 5408 12776
rect 7288 12724 7340 12776
rect 10508 12767 10560 12776
rect 3884 12656 3936 12708
rect 10508 12733 10517 12767
rect 10517 12733 10551 12767
rect 10551 12733 10560 12767
rect 10508 12724 10560 12733
rect 2504 12588 2556 12640
rect 5264 12588 5316 12640
rect 8760 12588 8812 12640
rect 9588 12656 9640 12708
rect 11980 12656 12032 12708
rect 11060 12588 11112 12640
rect 20260 12860 20312 12912
rect 24952 12860 25004 12912
rect 25228 12928 25280 12980
rect 27804 12971 27856 12980
rect 27804 12937 27813 12971
rect 27813 12937 27847 12971
rect 27847 12937 27856 12971
rect 27804 12928 27856 12937
rect 29552 12928 29604 12980
rect 29092 12860 29144 12912
rect 31576 12928 31628 12980
rect 32956 12971 33008 12980
rect 14464 12835 14516 12844
rect 14464 12801 14473 12835
rect 14473 12801 14507 12835
rect 14507 12801 14516 12835
rect 14464 12792 14516 12801
rect 14648 12835 14700 12844
rect 14648 12801 14657 12835
rect 14657 12801 14691 12835
rect 14691 12801 14700 12835
rect 14648 12792 14700 12801
rect 15108 12792 15160 12844
rect 18144 12835 18196 12844
rect 18144 12801 18162 12835
rect 18162 12801 18196 12835
rect 18144 12792 18196 12801
rect 18328 12792 18380 12844
rect 19156 12835 19208 12844
rect 19156 12801 19165 12835
rect 19165 12801 19199 12835
rect 19199 12801 19208 12835
rect 19156 12792 19208 12801
rect 14924 12724 14976 12776
rect 18420 12656 18472 12708
rect 20904 12792 20956 12844
rect 22100 12835 22152 12844
rect 22100 12801 22109 12835
rect 22109 12801 22143 12835
rect 22143 12801 22152 12835
rect 24124 12835 24176 12844
rect 22100 12792 22152 12801
rect 24124 12801 24133 12835
rect 24133 12801 24167 12835
rect 24167 12801 24176 12835
rect 24124 12792 24176 12801
rect 24676 12835 24728 12844
rect 24676 12801 24685 12835
rect 24685 12801 24719 12835
rect 24719 12801 24728 12835
rect 24676 12792 24728 12801
rect 31300 12792 31352 12844
rect 32404 12792 32456 12844
rect 32956 12937 32965 12971
rect 32965 12937 32999 12971
rect 32999 12937 33008 12971
rect 32956 12928 33008 12937
rect 35348 12928 35400 12980
rect 35624 12971 35676 12980
rect 35624 12937 35633 12971
rect 35633 12937 35667 12971
rect 35667 12937 35676 12971
rect 35624 12928 35676 12937
rect 38384 12928 38436 12980
rect 35256 12860 35308 12912
rect 35900 12835 35952 12844
rect 20536 12724 20588 12776
rect 24032 12724 24084 12776
rect 24308 12724 24360 12776
rect 17684 12588 17736 12640
rect 18880 12631 18932 12640
rect 18880 12597 18889 12631
rect 18889 12597 18923 12631
rect 18923 12597 18932 12631
rect 18880 12588 18932 12597
rect 19340 12656 19392 12708
rect 19432 12656 19484 12708
rect 24584 12656 24636 12708
rect 31852 12724 31904 12776
rect 35900 12801 35909 12835
rect 35909 12801 35943 12835
rect 35943 12801 35952 12835
rect 35900 12792 35952 12801
rect 36084 12835 36136 12844
rect 36084 12801 36093 12835
rect 36093 12801 36127 12835
rect 36127 12801 36136 12835
rect 36084 12792 36136 12801
rect 36268 12835 36320 12844
rect 36268 12801 36277 12835
rect 36277 12801 36311 12835
rect 36311 12801 36320 12835
rect 36268 12792 36320 12801
rect 38660 12792 38712 12844
rect 39028 12860 39080 12912
rect 39212 12792 39264 12844
rect 20812 12588 20864 12640
rect 22008 12588 22060 12640
rect 27068 12631 27120 12640
rect 27068 12597 27077 12631
rect 27077 12597 27111 12631
rect 27111 12597 27120 12631
rect 27068 12588 27120 12597
rect 34612 12656 34664 12708
rect 34704 12588 34756 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 2780 12384 2832 12436
rect 7104 12384 7156 12436
rect 7932 12427 7984 12436
rect 7932 12393 7941 12427
rect 7941 12393 7975 12427
rect 7975 12393 7984 12427
rect 7932 12384 7984 12393
rect 14832 12384 14884 12436
rect 19340 12384 19392 12436
rect 22560 12384 22612 12436
rect 23940 12384 23992 12436
rect 24952 12427 25004 12436
rect 24952 12393 24961 12427
rect 24961 12393 24995 12427
rect 24995 12393 25004 12427
rect 24952 12384 25004 12393
rect 29736 12384 29788 12436
rect 9496 12316 9548 12368
rect 12164 12359 12216 12368
rect 12164 12325 12173 12359
rect 12173 12325 12207 12359
rect 12207 12325 12216 12359
rect 12164 12316 12216 12325
rect 13728 12316 13780 12368
rect 28172 12359 28224 12368
rect 28172 12325 28181 12359
rect 28181 12325 28215 12359
rect 28215 12325 28224 12359
rect 28172 12316 28224 12325
rect 37648 12384 37700 12436
rect 37924 12384 37976 12436
rect 5356 12291 5408 12300
rect 5356 12257 5365 12291
rect 5365 12257 5399 12291
rect 5399 12257 5408 12291
rect 5356 12248 5408 12257
rect 12440 12248 12492 12300
rect 13268 12248 13320 12300
rect 16672 12248 16724 12300
rect 19432 12248 19484 12300
rect 20812 12291 20864 12300
rect 20812 12257 20821 12291
rect 20821 12257 20855 12291
rect 20855 12257 20864 12291
rect 20812 12248 20864 12257
rect 21088 12291 21140 12300
rect 21088 12257 21097 12291
rect 21097 12257 21131 12291
rect 21131 12257 21140 12291
rect 21088 12248 21140 12257
rect 2504 12223 2556 12232
rect 2504 12189 2513 12223
rect 2513 12189 2547 12223
rect 2547 12189 2556 12223
rect 2504 12180 2556 12189
rect 7932 12180 7984 12232
rect 11060 12223 11112 12232
rect 11060 12189 11094 12223
rect 11094 12189 11112 12223
rect 11060 12180 11112 12189
rect 14096 12180 14148 12232
rect 5172 12155 5224 12164
rect 5172 12121 5181 12155
rect 5181 12121 5215 12155
rect 5215 12121 5224 12155
rect 5172 12112 5224 12121
rect 5816 12112 5868 12164
rect 9680 12112 9732 12164
rect 13360 12155 13412 12164
rect 13360 12121 13369 12155
rect 13369 12121 13403 12155
rect 13403 12121 13412 12155
rect 13360 12112 13412 12121
rect 2688 12087 2740 12096
rect 2688 12053 2697 12087
rect 2697 12053 2731 12087
rect 2731 12053 2740 12087
rect 2688 12044 2740 12053
rect 4620 12044 4672 12096
rect 4896 12044 4948 12096
rect 5264 12087 5316 12096
rect 5264 12053 5273 12087
rect 5273 12053 5307 12087
rect 5307 12053 5316 12087
rect 5264 12044 5316 12053
rect 14280 12044 14332 12096
rect 14372 12087 14424 12096
rect 14372 12053 14381 12087
rect 14381 12053 14415 12087
rect 14415 12053 14424 12087
rect 14832 12223 14884 12232
rect 14832 12189 14841 12223
rect 14841 12189 14875 12223
rect 14875 12189 14884 12223
rect 14832 12180 14884 12189
rect 15108 12180 15160 12232
rect 15476 12180 15528 12232
rect 21824 12223 21876 12232
rect 21824 12189 21833 12223
rect 21833 12189 21867 12223
rect 21867 12189 21876 12223
rect 21824 12180 21876 12189
rect 22008 12223 22060 12232
rect 22008 12189 22017 12223
rect 22017 12189 22051 12223
rect 22051 12189 22060 12223
rect 22008 12180 22060 12189
rect 22560 12180 22612 12232
rect 24952 12180 25004 12232
rect 25044 12180 25096 12232
rect 25412 12180 25464 12232
rect 31300 12223 31352 12232
rect 31300 12189 31309 12223
rect 31309 12189 31343 12223
rect 31343 12189 31352 12223
rect 31300 12180 31352 12189
rect 31484 12223 31536 12232
rect 31484 12189 31493 12223
rect 31493 12189 31527 12223
rect 31527 12189 31536 12223
rect 31484 12180 31536 12189
rect 14924 12112 14976 12164
rect 18880 12112 18932 12164
rect 14372 12044 14424 12053
rect 14832 12044 14884 12096
rect 16948 12044 17000 12096
rect 20168 12112 20220 12164
rect 21548 12087 21600 12096
rect 21548 12053 21557 12087
rect 21557 12053 21591 12087
rect 21591 12053 21600 12087
rect 21548 12044 21600 12053
rect 25596 12112 25648 12164
rect 28356 12155 28408 12164
rect 28356 12121 28365 12155
rect 28365 12121 28399 12155
rect 28399 12121 28408 12155
rect 28356 12112 28408 12121
rect 32036 12180 32088 12232
rect 37280 12248 37332 12300
rect 37464 12248 37516 12300
rect 34796 12180 34848 12232
rect 37556 12180 37608 12232
rect 31852 12112 31904 12164
rect 35348 12112 35400 12164
rect 35532 12112 35584 12164
rect 24492 12087 24544 12096
rect 24492 12053 24501 12087
rect 24501 12053 24535 12087
rect 24535 12053 24544 12087
rect 24492 12044 24544 12053
rect 25964 12044 26016 12096
rect 27528 12087 27580 12096
rect 27528 12053 27537 12087
rect 27537 12053 27571 12087
rect 27571 12053 27580 12087
rect 27528 12044 27580 12053
rect 27712 12044 27764 12096
rect 32036 12044 32088 12096
rect 32404 12087 32456 12096
rect 32404 12053 32413 12087
rect 32413 12053 32447 12087
rect 32447 12053 32456 12087
rect 32404 12044 32456 12053
rect 35256 12044 35308 12096
rect 35900 12044 35952 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 5080 11840 5132 11892
rect 14740 11840 14792 11892
rect 2688 11772 2740 11824
rect 7932 11772 7984 11824
rect 2780 11704 2832 11756
rect 4896 11747 4948 11756
rect 4896 11713 4905 11747
rect 4905 11713 4939 11747
rect 4939 11713 4948 11747
rect 4896 11704 4948 11713
rect 6644 11747 6696 11756
rect 6644 11713 6653 11747
rect 6653 11713 6687 11747
rect 6687 11713 6696 11747
rect 6644 11704 6696 11713
rect 8760 11747 8812 11756
rect 14096 11772 14148 11824
rect 14280 11772 14332 11824
rect 14924 11840 14976 11892
rect 18144 11840 18196 11892
rect 18236 11840 18288 11892
rect 20260 11840 20312 11892
rect 21180 11840 21232 11892
rect 22468 11840 22520 11892
rect 8760 11713 8778 11747
rect 8778 11713 8812 11747
rect 8760 11704 8812 11713
rect 11980 11704 12032 11756
rect 13820 11747 13872 11756
rect 13820 11713 13829 11747
rect 13829 11713 13863 11747
rect 13863 11713 13872 11747
rect 13820 11704 13872 11713
rect 14004 11704 14056 11756
rect 4712 11636 4764 11688
rect 5080 11679 5132 11688
rect 5080 11645 5089 11679
rect 5089 11645 5123 11679
rect 5123 11645 5132 11679
rect 5080 11636 5132 11645
rect 6920 11636 6972 11688
rect 11520 11679 11572 11688
rect 11520 11645 11529 11679
rect 11529 11645 11563 11679
rect 11563 11645 11572 11679
rect 11520 11636 11572 11645
rect 14924 11750 14976 11756
rect 14924 11716 14933 11750
rect 14933 11716 14967 11750
rect 14967 11716 14976 11750
rect 14924 11704 14976 11716
rect 15108 11747 15160 11756
rect 15108 11713 15117 11747
rect 15117 11713 15151 11747
rect 15151 11713 15160 11747
rect 15108 11704 15160 11713
rect 15660 11704 15712 11756
rect 18144 11704 18196 11756
rect 18420 11747 18472 11756
rect 18420 11713 18429 11747
rect 18429 11713 18463 11747
rect 18463 11713 18472 11747
rect 18420 11704 18472 11713
rect 18512 11747 18564 11756
rect 18512 11713 18521 11747
rect 18521 11713 18555 11747
rect 18555 11713 18564 11747
rect 18512 11704 18564 11713
rect 19064 11704 19116 11756
rect 20168 11772 20220 11824
rect 21548 11772 21600 11824
rect 20536 11704 20588 11756
rect 22100 11704 22152 11756
rect 23572 11840 23624 11892
rect 25596 11883 25648 11892
rect 25596 11849 25605 11883
rect 25605 11849 25639 11883
rect 25639 11849 25648 11883
rect 25596 11840 25648 11849
rect 22652 11747 22704 11756
rect 22652 11713 22661 11747
rect 22661 11713 22695 11747
rect 22695 11713 22704 11747
rect 22652 11704 22704 11713
rect 15016 11636 15068 11688
rect 21640 11636 21692 11688
rect 22744 11636 22796 11688
rect 23664 11704 23716 11756
rect 24400 11704 24452 11756
rect 4712 11543 4764 11552
rect 4712 11509 4721 11543
rect 4721 11509 4755 11543
rect 4755 11509 4764 11543
rect 4712 11500 4764 11509
rect 4804 11500 4856 11552
rect 5448 11500 5500 11552
rect 7196 11500 7248 11552
rect 14464 11543 14516 11552
rect 14464 11509 14473 11543
rect 14473 11509 14507 11543
rect 14507 11509 14516 11543
rect 14464 11500 14516 11509
rect 15016 11500 15068 11552
rect 21272 11500 21324 11552
rect 26148 11704 26200 11756
rect 31484 11840 31536 11892
rect 34704 11840 34756 11892
rect 27528 11704 27580 11756
rect 26332 11636 26384 11688
rect 35256 11772 35308 11824
rect 36544 11840 36596 11892
rect 37280 11840 37332 11892
rect 38752 11840 38804 11892
rect 30748 11704 30800 11756
rect 31944 11704 31996 11756
rect 32404 11704 32456 11756
rect 32956 11704 33008 11756
rect 33048 11747 33100 11756
rect 33048 11713 33057 11747
rect 33057 11713 33091 11747
rect 33091 11713 33100 11747
rect 33048 11704 33100 11713
rect 35348 11747 35400 11756
rect 28356 11636 28408 11688
rect 35348 11713 35357 11747
rect 35357 11713 35391 11747
rect 35391 11713 35400 11747
rect 35348 11704 35400 11713
rect 35532 11747 35584 11756
rect 35532 11713 35541 11747
rect 35541 11713 35575 11747
rect 35575 11713 35584 11747
rect 35532 11704 35584 11713
rect 35624 11704 35676 11756
rect 36636 11772 36688 11824
rect 39212 11704 39264 11756
rect 39028 11679 39080 11688
rect 32312 11568 32364 11620
rect 39028 11645 39037 11679
rect 39037 11645 39071 11679
rect 39071 11645 39080 11679
rect 39028 11636 39080 11645
rect 58164 11611 58216 11620
rect 58164 11577 58173 11611
rect 58173 11577 58207 11611
rect 58207 11577 58216 11611
rect 58164 11568 58216 11577
rect 22192 11543 22244 11552
rect 22192 11509 22201 11543
rect 22201 11509 22235 11543
rect 22235 11509 22244 11543
rect 22192 11500 22244 11509
rect 22468 11500 22520 11552
rect 23664 11500 23716 11552
rect 24952 11500 25004 11552
rect 34520 11500 34572 11552
rect 35440 11500 35492 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 3792 11339 3844 11348
rect 3792 11305 3801 11339
rect 3801 11305 3835 11339
rect 3835 11305 3844 11339
rect 3792 11296 3844 11305
rect 3884 11160 3936 11212
rect 5264 11160 5316 11212
rect 6920 11296 6972 11348
rect 12440 11339 12492 11348
rect 12440 11305 12449 11339
rect 12449 11305 12483 11339
rect 12483 11305 12492 11339
rect 12440 11296 12492 11305
rect 13360 11296 13412 11348
rect 18144 11296 18196 11348
rect 18512 11339 18564 11348
rect 18512 11305 18521 11339
rect 18521 11305 18555 11339
rect 18555 11305 18564 11339
rect 18512 11296 18564 11305
rect 21180 11296 21232 11348
rect 6644 11228 6696 11280
rect 6736 11203 6788 11212
rect 6736 11169 6745 11203
rect 6745 11169 6779 11203
rect 6779 11169 6788 11203
rect 6736 11160 6788 11169
rect 7196 11160 7248 11212
rect 7288 11160 7340 11212
rect 2688 11092 2740 11144
rect 4712 11092 4764 11144
rect 4896 11092 4948 11144
rect 5632 11024 5684 11076
rect 4712 10956 4764 11008
rect 4988 10956 5040 11008
rect 6368 10999 6420 11008
rect 6368 10965 6377 10999
rect 6377 10965 6411 10999
rect 6411 10965 6420 10999
rect 6368 10956 6420 10965
rect 7472 11092 7524 11144
rect 15936 11228 15988 11280
rect 17224 11228 17276 11280
rect 21272 11228 21324 11280
rect 15660 11160 15712 11212
rect 22744 11296 22796 11348
rect 26148 11339 26200 11348
rect 26148 11305 26157 11339
rect 26157 11305 26191 11339
rect 26191 11305 26200 11339
rect 26148 11296 26200 11305
rect 30196 11296 30248 11348
rect 30380 11296 30432 11348
rect 24492 11228 24544 11280
rect 33048 11296 33100 11348
rect 34520 11296 34572 11348
rect 21640 11203 21692 11212
rect 21640 11169 21649 11203
rect 21649 11169 21683 11203
rect 21683 11169 21692 11203
rect 21640 11160 21692 11169
rect 23572 11203 23624 11212
rect 23572 11169 23581 11203
rect 23581 11169 23615 11203
rect 23615 11169 23624 11203
rect 23572 11160 23624 11169
rect 24584 11160 24636 11212
rect 26332 11160 26384 11212
rect 29092 11160 29144 11212
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 11520 11135 11572 11144
rect 11520 11101 11529 11135
rect 11529 11101 11563 11135
rect 11563 11101 11572 11135
rect 11520 11092 11572 11101
rect 14464 11092 14516 11144
rect 15476 11092 15528 11144
rect 14832 11024 14884 11076
rect 17776 11067 17828 11076
rect 17776 11033 17785 11067
rect 17785 11033 17819 11067
rect 17819 11033 17828 11067
rect 17776 11024 17828 11033
rect 18512 11024 18564 11076
rect 19340 11024 19392 11076
rect 20812 11024 20864 11076
rect 21456 11024 21508 11076
rect 22192 11024 22244 11076
rect 23480 11135 23532 11144
rect 23480 11101 23489 11135
rect 23489 11101 23523 11135
rect 23523 11101 23532 11135
rect 23664 11135 23716 11144
rect 23480 11092 23532 11101
rect 23664 11101 23673 11135
rect 23673 11101 23707 11135
rect 23707 11101 23716 11135
rect 23664 11092 23716 11101
rect 25964 11135 26016 11144
rect 25964 11101 25973 11135
rect 25973 11101 26007 11135
rect 26007 11101 26016 11135
rect 25964 11092 26016 11101
rect 30196 11092 30248 11144
rect 31852 11160 31904 11212
rect 30840 11135 30892 11144
rect 30840 11101 30849 11135
rect 30849 11101 30883 11135
rect 30883 11101 30892 11135
rect 30840 11092 30892 11101
rect 25044 11024 25096 11076
rect 25780 11067 25832 11076
rect 25780 11033 25789 11067
rect 25789 11033 25823 11067
rect 25823 11033 25832 11067
rect 25780 11024 25832 11033
rect 30472 11024 30524 11076
rect 30564 11024 30616 11076
rect 31300 11092 31352 11144
rect 32036 11135 32088 11144
rect 32036 11101 32045 11135
rect 32045 11101 32079 11135
rect 32079 11101 32088 11135
rect 32036 11092 32088 11101
rect 32312 11135 32364 11144
rect 32312 11101 32321 11135
rect 32321 11101 32355 11135
rect 32355 11101 32364 11135
rect 32312 11092 32364 11101
rect 35440 11160 35492 11212
rect 35256 11092 35308 11144
rect 36544 11135 36596 11144
rect 36544 11101 36553 11135
rect 36553 11101 36587 11135
rect 36587 11101 36596 11135
rect 36544 11092 36596 11101
rect 36636 11092 36688 11144
rect 39028 11228 39080 11280
rect 37556 11024 37608 11076
rect 38016 11067 38068 11076
rect 38016 11033 38025 11067
rect 38025 11033 38059 11067
rect 38059 11033 38068 11067
rect 38016 11024 38068 11033
rect 8944 10999 8996 11008
rect 8944 10965 8953 10999
rect 8953 10965 8987 10999
rect 8987 10965 8996 10999
rect 8944 10956 8996 10965
rect 14188 10956 14240 11008
rect 18236 10956 18288 11008
rect 19248 10956 19300 11008
rect 20076 10956 20128 11008
rect 23020 10999 23072 11008
rect 23020 10965 23029 10999
rect 23029 10965 23063 10999
rect 23063 10965 23072 10999
rect 23020 10956 23072 10965
rect 35348 10956 35400 11008
rect 38752 11024 38804 11076
rect 40132 11024 40184 11076
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 5356 10752 5408 10804
rect 7472 10752 7524 10804
rect 9128 10752 9180 10804
rect 14004 10795 14056 10804
rect 14004 10761 14013 10795
rect 14013 10761 14047 10795
rect 14047 10761 14056 10795
rect 14004 10752 14056 10761
rect 22652 10752 22704 10804
rect 23204 10752 23256 10804
rect 27160 10752 27212 10804
rect 4620 10684 4672 10736
rect 5264 10684 5316 10736
rect 8944 10684 8996 10736
rect 14372 10684 14424 10736
rect 23020 10684 23072 10736
rect 2044 10616 2096 10668
rect 4988 10616 5040 10668
rect 7656 10659 7708 10668
rect 7656 10625 7665 10659
rect 7665 10625 7699 10659
rect 7699 10625 7708 10659
rect 7656 10616 7708 10625
rect 7932 10616 7984 10668
rect 2688 10548 2740 10600
rect 12624 10616 12676 10668
rect 22192 10616 22244 10668
rect 28816 10684 28868 10736
rect 30840 10752 30892 10804
rect 36544 10752 36596 10804
rect 38016 10752 38068 10804
rect 24584 10659 24636 10668
rect 24584 10625 24593 10659
rect 24593 10625 24627 10659
rect 24627 10625 24636 10659
rect 24584 10616 24636 10625
rect 25044 10659 25096 10668
rect 25044 10625 25053 10659
rect 25053 10625 25087 10659
rect 25087 10625 25096 10659
rect 25044 10616 25096 10625
rect 25320 10659 25372 10668
rect 25320 10625 25354 10659
rect 25354 10625 25372 10659
rect 25320 10616 25372 10625
rect 25780 10616 25832 10668
rect 30748 10684 30800 10736
rect 37924 10684 37976 10736
rect 40132 10727 40184 10736
rect 40132 10693 40166 10727
rect 40166 10693 40184 10727
rect 40132 10684 40184 10693
rect 15384 10591 15436 10600
rect 15384 10557 15393 10591
rect 15393 10557 15427 10591
rect 15427 10557 15436 10591
rect 15384 10548 15436 10557
rect 24308 10591 24360 10600
rect 24308 10557 24317 10591
rect 24317 10557 24351 10591
rect 24351 10557 24360 10591
rect 24308 10548 24360 10557
rect 15476 10480 15528 10532
rect 22836 10480 22888 10532
rect 29092 10480 29144 10532
rect 30564 10616 30616 10668
rect 30840 10659 30892 10668
rect 30840 10625 30849 10659
rect 30849 10625 30883 10659
rect 30883 10625 30892 10659
rect 30840 10616 30892 10625
rect 34796 10616 34848 10668
rect 35348 10659 35400 10668
rect 35348 10625 35382 10659
rect 35382 10625 35400 10659
rect 35348 10616 35400 10625
rect 29368 10480 29420 10532
rect 2412 10455 2464 10464
rect 2412 10421 2421 10455
rect 2421 10421 2455 10455
rect 2455 10421 2464 10455
rect 2412 10412 2464 10421
rect 9772 10412 9824 10464
rect 10232 10455 10284 10464
rect 10232 10421 10241 10455
rect 10241 10421 10275 10455
rect 10275 10421 10284 10455
rect 10232 10412 10284 10421
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 12440 10412 12492 10421
rect 12808 10412 12860 10464
rect 16580 10412 16632 10464
rect 18420 10412 18472 10464
rect 19064 10412 19116 10464
rect 19340 10412 19392 10464
rect 19616 10455 19668 10464
rect 19616 10421 19625 10455
rect 19625 10421 19659 10455
rect 19659 10421 19668 10455
rect 19616 10412 19668 10421
rect 26332 10412 26384 10464
rect 28540 10412 28592 10464
rect 38936 10455 38988 10464
rect 38936 10421 38945 10455
rect 38945 10421 38979 10455
rect 38979 10421 38988 10455
rect 38936 10412 38988 10421
rect 58164 10455 58216 10464
rect 58164 10421 58173 10455
rect 58173 10421 58207 10455
rect 58207 10421 58216 10455
rect 58164 10412 58216 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2044 10251 2096 10260
rect 2044 10217 2053 10251
rect 2053 10217 2087 10251
rect 2087 10217 2096 10251
rect 2044 10208 2096 10217
rect 5080 10208 5132 10260
rect 5448 10208 5500 10260
rect 7012 10251 7064 10260
rect 7012 10217 7021 10251
rect 7021 10217 7055 10251
rect 7055 10217 7064 10251
rect 7012 10208 7064 10217
rect 7656 10208 7708 10260
rect 21272 10251 21324 10260
rect 21272 10217 21281 10251
rect 21281 10217 21315 10251
rect 21315 10217 21324 10251
rect 21272 10208 21324 10217
rect 22192 10251 22244 10260
rect 22192 10217 22201 10251
rect 22201 10217 22235 10251
rect 22235 10217 22244 10251
rect 22192 10208 22244 10217
rect 25320 10208 25372 10260
rect 26424 10251 26476 10260
rect 26424 10217 26433 10251
rect 26433 10217 26467 10251
rect 26467 10217 26476 10251
rect 26424 10208 26476 10217
rect 27988 10251 28040 10260
rect 27988 10217 27997 10251
rect 27997 10217 28031 10251
rect 28031 10217 28040 10251
rect 27988 10208 28040 10217
rect 29368 10208 29420 10260
rect 30656 10251 30708 10260
rect 30656 10217 30665 10251
rect 30665 10217 30699 10251
rect 30699 10217 30708 10251
rect 30656 10208 30708 10217
rect 32496 10251 32548 10260
rect 32496 10217 32505 10251
rect 32505 10217 32539 10251
rect 32539 10217 32548 10251
rect 32496 10208 32548 10217
rect 36636 10208 36688 10260
rect 3700 10072 3752 10124
rect 5172 10115 5224 10124
rect 5172 10081 5181 10115
rect 5181 10081 5215 10115
rect 5215 10081 5224 10115
rect 5172 10072 5224 10081
rect 9680 10072 9732 10124
rect 10600 10140 10652 10192
rect 15200 10140 15252 10192
rect 19616 10140 19668 10192
rect 3608 10004 3660 10056
rect 2228 9936 2280 9988
rect 2688 9936 2740 9988
rect 4988 9979 5040 9988
rect 4988 9945 4997 9979
rect 4997 9945 5031 9979
rect 5031 9945 5040 9979
rect 4988 9936 5040 9945
rect 10232 10004 10284 10056
rect 16580 10072 16632 10124
rect 20444 10072 20496 10124
rect 21272 10072 21324 10124
rect 24308 10072 24360 10124
rect 10600 10004 10652 10056
rect 12808 10004 12860 10056
rect 15568 10004 15620 10056
rect 16764 10004 16816 10056
rect 22100 10004 22152 10056
rect 23388 10004 23440 10056
rect 24032 10004 24084 10056
rect 24952 10047 25004 10056
rect 24952 10013 24961 10047
rect 24961 10013 24995 10047
rect 24995 10013 25004 10047
rect 24952 10004 25004 10013
rect 27712 10140 27764 10192
rect 28632 10140 28684 10192
rect 29276 10140 29328 10192
rect 11520 9936 11572 9988
rect 12440 9936 12492 9988
rect 20720 9936 20772 9988
rect 25964 10004 26016 10056
rect 26240 10047 26292 10056
rect 26240 10013 26249 10047
rect 26249 10013 26283 10047
rect 26283 10013 26292 10047
rect 27436 10047 27488 10056
rect 26240 10004 26292 10013
rect 27436 10013 27445 10047
rect 27445 10013 27479 10047
rect 27479 10013 27488 10047
rect 27436 10004 27488 10013
rect 28264 10072 28316 10124
rect 27804 10047 27856 10056
rect 27804 10013 27813 10047
rect 27813 10013 27847 10047
rect 27847 10013 27856 10047
rect 27804 10004 27856 10013
rect 28448 10047 28500 10056
rect 28448 10013 28457 10047
rect 28457 10013 28491 10047
rect 28491 10013 28500 10047
rect 28448 10004 28500 10013
rect 28816 10047 28868 10056
rect 28816 10013 28825 10047
rect 28825 10013 28859 10047
rect 28859 10013 28868 10047
rect 28816 10004 28868 10013
rect 30656 10004 30708 10056
rect 37924 10208 37976 10260
rect 37096 10004 37148 10056
rect 38108 10047 38160 10056
rect 38108 10013 38117 10047
rect 38117 10013 38151 10047
rect 38151 10013 38160 10047
rect 38108 10004 38160 10013
rect 39028 10072 39080 10124
rect 3424 9868 3476 9920
rect 3884 9911 3936 9920
rect 3884 9877 3893 9911
rect 3893 9877 3927 9911
rect 3927 9877 3936 9911
rect 3884 9868 3936 9877
rect 9680 9868 9732 9920
rect 12808 9868 12860 9920
rect 13268 9868 13320 9920
rect 22468 9868 22520 9920
rect 27528 9936 27580 9988
rect 26332 9868 26384 9920
rect 29644 9936 29696 9988
rect 30748 9936 30800 9988
rect 37280 9936 37332 9988
rect 38844 9868 38896 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 15016 9664 15068 9716
rect 2412 9596 2464 9648
rect 10508 9596 10560 9648
rect 20628 9596 20680 9648
rect 24952 9664 25004 9716
rect 22284 9596 22336 9648
rect 23020 9596 23072 9648
rect 5540 9571 5592 9580
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 9680 9528 9732 9580
rect 5632 9460 5684 9512
rect 5908 9460 5960 9512
rect 12624 9571 12676 9580
rect 12624 9537 12633 9571
rect 12633 9537 12667 9571
rect 12667 9537 12676 9571
rect 12624 9528 12676 9537
rect 12808 9571 12860 9580
rect 12808 9537 12817 9571
rect 12817 9537 12851 9571
rect 12851 9537 12860 9571
rect 12808 9528 12860 9537
rect 10784 9460 10836 9512
rect 10600 9392 10652 9444
rect 15292 9460 15344 9512
rect 13268 9392 13320 9444
rect 15200 9392 15252 9444
rect 20168 9528 20220 9580
rect 22468 9528 22520 9580
rect 22744 9571 22796 9580
rect 22744 9537 22753 9571
rect 22753 9537 22787 9571
rect 22787 9537 22796 9571
rect 22744 9528 22796 9537
rect 25780 9664 25832 9716
rect 29644 9707 29696 9716
rect 29644 9673 29653 9707
rect 29653 9673 29687 9707
rect 29687 9673 29696 9707
rect 29644 9664 29696 9673
rect 30840 9664 30892 9716
rect 31576 9707 31628 9716
rect 31576 9673 31585 9707
rect 31585 9673 31619 9707
rect 31619 9673 31628 9707
rect 31576 9664 31628 9673
rect 38108 9664 38160 9716
rect 26332 9596 26384 9648
rect 29828 9596 29880 9648
rect 31852 9596 31904 9648
rect 28540 9571 28592 9580
rect 28540 9537 28574 9571
rect 28574 9537 28592 9571
rect 19248 9460 19300 9512
rect 22928 9435 22980 9444
rect 22928 9401 22937 9435
rect 22937 9401 22971 9435
rect 22971 9401 22980 9435
rect 22928 9392 22980 9401
rect 28540 9528 28592 9537
rect 30472 9571 30524 9580
rect 30472 9537 30506 9571
rect 30506 9537 30524 9571
rect 30472 9528 30524 9537
rect 32036 9528 32088 9580
rect 32312 9571 32364 9580
rect 32312 9537 32321 9571
rect 32321 9537 32355 9571
rect 32355 9537 32364 9571
rect 32312 9528 32364 9537
rect 32864 9596 32916 9648
rect 34796 9596 34848 9648
rect 38936 9596 38988 9648
rect 34704 9528 34756 9580
rect 25780 9392 25832 9444
rect 2320 9324 2372 9376
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 6276 9324 6328 9376
rect 11704 9324 11756 9376
rect 13084 9324 13136 9376
rect 15660 9367 15712 9376
rect 15660 9333 15669 9367
rect 15669 9333 15703 9367
rect 15703 9333 15712 9367
rect 15660 9324 15712 9333
rect 22744 9324 22796 9376
rect 26240 9324 26292 9376
rect 27068 9324 27120 9376
rect 34520 9392 34572 9444
rect 35256 9392 35308 9444
rect 35624 9528 35676 9580
rect 37556 9528 37608 9580
rect 37372 9460 37424 9512
rect 38844 9528 38896 9580
rect 37740 9392 37792 9444
rect 32680 9324 32732 9376
rect 35440 9324 35492 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 9404 9120 9456 9172
rect 9680 9120 9732 9172
rect 12716 9120 12768 9172
rect 13268 9120 13320 9172
rect 14280 9120 14332 9172
rect 14740 9120 14792 9172
rect 18604 9120 18656 9172
rect 18972 9120 19024 9172
rect 20536 9120 20588 9172
rect 20720 9120 20772 9172
rect 22284 9120 22336 9172
rect 23664 9120 23716 9172
rect 27068 9120 27120 9172
rect 32312 9120 32364 9172
rect 33508 9120 33560 9172
rect 35624 9120 35676 9172
rect 37832 9120 37884 9172
rect 38936 9120 38988 9172
rect 9588 9095 9640 9104
rect 9588 9061 9597 9095
rect 9597 9061 9631 9095
rect 9631 9061 9640 9095
rect 9588 9052 9640 9061
rect 12256 9052 12308 9104
rect 14464 9052 14516 9104
rect 27804 9052 27856 9104
rect 3424 8984 3476 9036
rect 5724 8984 5776 9036
rect 9312 8984 9364 9036
rect 11704 9027 11756 9036
rect 5080 8959 5132 8968
rect 5080 8925 5089 8959
rect 5089 8925 5123 8959
rect 5123 8925 5132 8959
rect 5080 8916 5132 8925
rect 10600 8916 10652 8968
rect 11244 8916 11296 8968
rect 11704 8993 11713 9027
rect 11713 8993 11747 9027
rect 11747 8993 11756 9027
rect 11704 8984 11756 8993
rect 11888 8984 11940 9036
rect 21824 8984 21876 9036
rect 22744 8984 22796 9036
rect 26240 8984 26292 9036
rect 5540 8848 5592 8900
rect 6920 8848 6972 8900
rect 7472 8848 7524 8900
rect 8760 8848 8812 8900
rect 9220 8848 9272 8900
rect 12256 8916 12308 8968
rect 13084 8959 13136 8968
rect 13084 8925 13093 8959
rect 13093 8925 13127 8959
rect 13127 8925 13136 8959
rect 13084 8916 13136 8925
rect 15384 8916 15436 8968
rect 19248 8959 19300 8968
rect 19248 8925 19257 8959
rect 19257 8925 19291 8959
rect 19291 8925 19300 8959
rect 19248 8916 19300 8925
rect 20628 8916 20680 8968
rect 21272 8959 21324 8968
rect 21272 8925 21281 8959
rect 21281 8925 21315 8959
rect 21315 8925 21324 8959
rect 21272 8916 21324 8925
rect 21732 8916 21784 8968
rect 31576 8984 31628 9036
rect 33876 9052 33928 9104
rect 28816 8916 28868 8968
rect 30748 8916 30800 8968
rect 31668 8959 31720 8968
rect 31668 8925 31677 8959
rect 31677 8925 31711 8959
rect 31711 8925 31720 8959
rect 31668 8916 31720 8925
rect 32588 8984 32640 9036
rect 32404 8916 32456 8968
rect 32956 8959 33008 8968
rect 32956 8925 32965 8959
rect 32965 8925 32999 8959
rect 32999 8925 33008 8959
rect 32956 8916 33008 8925
rect 35808 8984 35860 9036
rect 34796 8916 34848 8968
rect 36268 8916 36320 8968
rect 37004 8959 37056 8968
rect 37004 8925 37013 8959
rect 37013 8925 37047 8959
rect 37047 8925 37056 8959
rect 37004 8916 37056 8925
rect 37280 8916 37332 8968
rect 38752 8916 38804 8968
rect 58164 8959 58216 8968
rect 58164 8925 58173 8959
rect 58173 8925 58207 8959
rect 58207 8925 58216 8959
rect 58164 8916 58216 8925
rect 11888 8848 11940 8900
rect 3240 8823 3292 8832
rect 3240 8789 3249 8823
rect 3249 8789 3283 8823
rect 3283 8789 3292 8823
rect 3240 8780 3292 8789
rect 4804 8780 4856 8832
rect 7196 8823 7248 8832
rect 7196 8789 7205 8823
rect 7205 8789 7239 8823
rect 7239 8789 7248 8823
rect 7196 8780 7248 8789
rect 8116 8780 8168 8832
rect 9588 8780 9640 8832
rect 12716 8780 12768 8832
rect 17684 8848 17736 8900
rect 18788 8848 18840 8900
rect 31392 8848 31444 8900
rect 16396 8780 16448 8832
rect 17960 8780 18012 8832
rect 20168 8780 20220 8832
rect 28264 8780 28316 8832
rect 32312 8848 32364 8900
rect 34980 8891 35032 8900
rect 34980 8857 35014 8891
rect 35014 8857 35032 8891
rect 34980 8848 35032 8857
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 4988 8576 5040 8628
rect 8208 8576 8260 8628
rect 9680 8619 9732 8628
rect 9680 8585 9689 8619
rect 9689 8585 9723 8619
rect 9723 8585 9732 8619
rect 9680 8576 9732 8585
rect 10140 8619 10192 8628
rect 10140 8585 10149 8619
rect 10149 8585 10183 8619
rect 10183 8585 10192 8619
rect 10140 8576 10192 8585
rect 13360 8576 13412 8628
rect 7012 8508 7064 8560
rect 9772 8508 9824 8560
rect 5632 8440 5684 8492
rect 6644 8483 6696 8492
rect 6644 8449 6653 8483
rect 6653 8449 6687 8483
rect 6687 8449 6696 8483
rect 6644 8440 6696 8449
rect 8760 8440 8812 8492
rect 5908 8372 5960 8424
rect 6368 8415 6420 8424
rect 6368 8381 6377 8415
rect 6377 8381 6411 8415
rect 6411 8381 6420 8415
rect 6368 8372 6420 8381
rect 8576 8415 8628 8424
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 10876 8440 10928 8492
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 12808 8508 12860 8560
rect 12256 8483 12308 8492
rect 12256 8449 12265 8483
rect 12265 8449 12299 8483
rect 12299 8449 12308 8483
rect 12256 8440 12308 8449
rect 14280 8576 14332 8628
rect 14464 8576 14516 8628
rect 17132 8576 17184 8628
rect 18236 8576 18288 8628
rect 14004 8483 14056 8492
rect 14004 8449 14013 8483
rect 14013 8449 14047 8483
rect 14047 8449 14056 8483
rect 14004 8440 14056 8449
rect 9312 8372 9364 8424
rect 11796 8372 11848 8424
rect 11980 8415 12032 8424
rect 11980 8381 11989 8415
rect 11989 8381 12023 8415
rect 12023 8381 12032 8415
rect 12808 8415 12860 8424
rect 11980 8372 12032 8381
rect 12808 8381 12817 8415
rect 12817 8381 12851 8415
rect 12851 8381 12860 8415
rect 15476 8508 15528 8560
rect 14832 8440 14884 8492
rect 15016 8483 15068 8492
rect 15016 8449 15050 8483
rect 15050 8449 15068 8483
rect 18144 8508 18196 8560
rect 15016 8440 15068 8449
rect 12808 8372 12860 8381
rect 1584 8347 1636 8356
rect 1584 8313 1593 8347
rect 1593 8313 1627 8347
rect 1627 8313 1636 8347
rect 1584 8304 1636 8313
rect 2136 8347 2188 8356
rect 2136 8313 2145 8347
rect 2145 8313 2179 8347
rect 2179 8313 2188 8347
rect 2136 8304 2188 8313
rect 2596 8304 2648 8356
rect 4620 8304 4672 8356
rect 7564 8304 7616 8356
rect 8760 8304 8812 8356
rect 10692 8347 10744 8356
rect 3884 8236 3936 8288
rect 5540 8236 5592 8288
rect 8024 8236 8076 8288
rect 8852 8236 8904 8288
rect 9680 8236 9732 8288
rect 10692 8313 10701 8347
rect 10701 8313 10735 8347
rect 10735 8313 10744 8347
rect 10692 8304 10744 8313
rect 11612 8304 11664 8356
rect 17132 8440 17184 8492
rect 18788 8576 18840 8628
rect 20720 8576 20772 8628
rect 21272 8576 21324 8628
rect 30288 8576 30340 8628
rect 32128 8576 32180 8628
rect 20168 8551 20220 8560
rect 20168 8517 20177 8551
rect 20177 8517 20211 8551
rect 20211 8517 20220 8551
rect 20168 8508 20220 8517
rect 16488 8372 16540 8424
rect 17500 8372 17552 8424
rect 18420 8483 18472 8492
rect 18420 8449 18429 8483
rect 18429 8449 18463 8483
rect 18463 8449 18472 8483
rect 18420 8440 18472 8449
rect 18604 8440 18656 8492
rect 19432 8440 19484 8492
rect 21364 8440 21416 8492
rect 21824 8483 21876 8492
rect 21824 8449 21833 8483
rect 21833 8449 21867 8483
rect 21867 8449 21876 8483
rect 21824 8440 21876 8449
rect 22100 8483 22152 8492
rect 22100 8449 22109 8483
rect 22109 8449 22143 8483
rect 22143 8449 22152 8483
rect 22100 8440 22152 8449
rect 22652 8440 22704 8492
rect 23664 8483 23716 8492
rect 23664 8449 23673 8483
rect 23673 8449 23707 8483
rect 23707 8449 23716 8483
rect 23664 8440 23716 8449
rect 24308 8508 24360 8560
rect 24032 8483 24084 8492
rect 16856 8304 16908 8356
rect 18144 8304 18196 8356
rect 23296 8372 23348 8424
rect 24032 8449 24041 8483
rect 24041 8449 24075 8483
rect 24075 8449 24084 8483
rect 24032 8440 24084 8449
rect 27620 8440 27672 8492
rect 28632 8508 28684 8560
rect 31392 8508 31444 8560
rect 32312 8551 32364 8560
rect 32312 8517 32321 8551
rect 32321 8517 32355 8551
rect 32355 8517 32364 8551
rect 32312 8508 32364 8517
rect 33692 8576 33744 8628
rect 34520 8619 34572 8628
rect 34520 8585 34529 8619
rect 34529 8585 34563 8619
rect 34563 8585 34572 8619
rect 34520 8576 34572 8585
rect 34980 8619 35032 8628
rect 34980 8585 34989 8619
rect 34989 8585 35023 8619
rect 35023 8585 35032 8619
rect 34980 8576 35032 8585
rect 37004 8576 37056 8628
rect 28264 8483 28316 8492
rect 28264 8449 28273 8483
rect 28273 8449 28307 8483
rect 28307 8449 28316 8483
rect 28264 8440 28316 8449
rect 29276 8483 29328 8492
rect 29276 8449 29285 8483
rect 29285 8449 29319 8483
rect 29319 8449 29328 8483
rect 29276 8440 29328 8449
rect 32128 8483 32180 8492
rect 28816 8372 28868 8424
rect 32128 8449 32137 8483
rect 32137 8449 32171 8483
rect 32171 8449 32180 8483
rect 32128 8440 32180 8449
rect 32588 8440 32640 8492
rect 35808 8508 35860 8560
rect 37832 8508 37884 8560
rect 35440 8483 35492 8492
rect 35440 8449 35449 8483
rect 35449 8449 35483 8483
rect 35483 8449 35492 8483
rect 35440 8440 35492 8449
rect 36268 8440 36320 8492
rect 23480 8304 23532 8356
rect 27620 8304 27672 8356
rect 27896 8304 27948 8356
rect 37740 8440 37792 8492
rect 37280 8372 37332 8424
rect 23204 8236 23256 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 9588 8032 9640 8084
rect 11980 8032 12032 8084
rect 17132 8075 17184 8084
rect 3424 7964 3476 8016
rect 4712 7964 4764 8016
rect 4988 7896 5040 7948
rect 5632 7964 5684 8016
rect 7932 7964 7984 8016
rect 3884 7828 3936 7880
rect 4068 7828 4120 7880
rect 5724 7896 5776 7948
rect 5448 7871 5500 7880
rect 2688 7760 2740 7812
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 5448 7828 5500 7837
rect 6736 7828 6788 7880
rect 7472 7828 7524 7880
rect 6000 7760 6052 7812
rect 8024 7760 8076 7812
rect 9220 7828 9272 7880
rect 9496 7871 9548 7880
rect 9496 7837 9505 7871
rect 9505 7837 9539 7871
rect 9539 7837 9548 7871
rect 9496 7828 9548 7837
rect 9680 7871 9732 7880
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 15108 7964 15160 8016
rect 17132 8041 17141 8075
rect 17141 8041 17175 8075
rect 17175 8041 17184 8075
rect 17132 8032 17184 8041
rect 17684 8075 17736 8084
rect 17684 8041 17693 8075
rect 17693 8041 17727 8075
rect 17727 8041 17736 8075
rect 17684 8032 17736 8041
rect 20076 8032 20128 8084
rect 27160 8032 27212 8084
rect 10600 7939 10652 7948
rect 10600 7905 10609 7939
rect 10609 7905 10643 7939
rect 10643 7905 10652 7939
rect 10600 7896 10652 7905
rect 14464 7896 14516 7948
rect 17132 7896 17184 7948
rect 9680 7828 9732 7837
rect 13360 7828 13412 7880
rect 14280 7828 14332 7880
rect 14740 7828 14792 7880
rect 10048 7760 10100 7812
rect 13912 7760 13964 7812
rect 17868 7828 17920 7880
rect 18144 7871 18196 7880
rect 18144 7837 18153 7871
rect 18153 7837 18187 7871
rect 18187 7837 18196 7871
rect 18144 7828 18196 7837
rect 19064 7828 19116 7880
rect 25964 7964 26016 8016
rect 28724 8032 28776 8084
rect 20720 7896 20772 7948
rect 20812 7828 20864 7880
rect 22100 7828 22152 7880
rect 18236 7760 18288 7812
rect 18696 7760 18748 7812
rect 23204 7828 23256 7880
rect 24952 7828 25004 7880
rect 27804 7871 27856 7880
rect 27804 7837 27813 7871
rect 27813 7837 27847 7871
rect 27847 7837 27856 7871
rect 27804 7828 27856 7837
rect 31668 7828 31720 7880
rect 35348 7896 35400 7948
rect 35532 7828 35584 7880
rect 35624 7871 35676 7880
rect 35624 7837 35633 7871
rect 35633 7837 35667 7871
rect 35667 7837 35676 7871
rect 58164 7871 58216 7880
rect 35624 7828 35676 7837
rect 58164 7837 58173 7871
rect 58173 7837 58207 7871
rect 58207 7837 58216 7871
rect 58164 7828 58216 7837
rect 25320 7760 25372 7812
rect 28264 7760 28316 7812
rect 31484 7760 31536 7812
rect 37188 7760 37240 7812
rect 1492 7735 1544 7744
rect 1492 7701 1501 7735
rect 1501 7701 1535 7735
rect 1535 7701 1544 7735
rect 1492 7692 1544 7701
rect 2504 7735 2556 7744
rect 2504 7701 2513 7735
rect 2513 7701 2547 7735
rect 2547 7701 2556 7735
rect 2504 7692 2556 7701
rect 3792 7692 3844 7744
rect 3976 7735 4028 7744
rect 3976 7701 3985 7735
rect 3985 7701 4019 7735
rect 4019 7701 4028 7735
rect 3976 7692 4028 7701
rect 4712 7735 4764 7744
rect 4712 7701 4721 7735
rect 4721 7701 4755 7735
rect 4755 7701 4764 7735
rect 4712 7692 4764 7701
rect 5172 7692 5224 7744
rect 8944 7735 8996 7744
rect 8944 7701 8953 7735
rect 8953 7701 8987 7735
rect 8987 7701 8996 7735
rect 8944 7692 8996 7701
rect 9496 7692 9548 7744
rect 10784 7692 10836 7744
rect 12072 7692 12124 7744
rect 14924 7692 14976 7744
rect 15476 7692 15528 7744
rect 16672 7735 16724 7744
rect 16672 7701 16681 7735
rect 16681 7701 16715 7735
rect 16715 7701 16724 7735
rect 16672 7692 16724 7701
rect 21272 7735 21324 7744
rect 21272 7701 21281 7735
rect 21281 7701 21315 7735
rect 21315 7701 21324 7735
rect 21272 7692 21324 7701
rect 22560 7692 22612 7744
rect 24676 7692 24728 7744
rect 26884 7735 26936 7744
rect 26884 7701 26893 7735
rect 26893 7701 26927 7735
rect 26927 7701 26936 7735
rect 26884 7692 26936 7701
rect 30656 7735 30708 7744
rect 30656 7701 30665 7735
rect 30665 7701 30699 7735
rect 30699 7701 30708 7735
rect 30656 7692 30708 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 2228 7395 2280 7404
rect 2228 7361 2237 7395
rect 2237 7361 2271 7395
rect 2271 7361 2280 7395
rect 2228 7352 2280 7361
rect 3516 7531 3568 7540
rect 3516 7497 3525 7531
rect 3525 7497 3559 7531
rect 3559 7497 3568 7531
rect 3516 7488 3568 7497
rect 5172 7531 5224 7540
rect 5172 7497 5181 7531
rect 5181 7497 5215 7531
rect 5215 7497 5224 7531
rect 5172 7488 5224 7497
rect 7932 7531 7984 7540
rect 7932 7497 7941 7531
rect 7941 7497 7975 7531
rect 7975 7497 7984 7531
rect 7932 7488 7984 7497
rect 8024 7488 8076 7540
rect 9496 7488 9548 7540
rect 10140 7488 10192 7540
rect 10324 7488 10376 7540
rect 14556 7488 14608 7540
rect 15016 7531 15068 7540
rect 15016 7497 15025 7531
rect 15025 7497 15059 7531
rect 15059 7497 15068 7531
rect 15016 7488 15068 7497
rect 3976 7420 4028 7472
rect 5540 7420 5592 7472
rect 3792 7352 3844 7404
rect 5080 7352 5132 7404
rect 3700 7327 3752 7336
rect 3700 7293 3709 7327
rect 3709 7293 3743 7327
rect 3743 7293 3752 7327
rect 3700 7284 3752 7293
rect 3884 7284 3936 7336
rect 12716 7463 12768 7472
rect 12716 7429 12734 7463
rect 12734 7429 12768 7463
rect 17868 7488 17920 7540
rect 23112 7488 23164 7540
rect 23296 7531 23348 7540
rect 23296 7497 23305 7531
rect 23305 7497 23339 7531
rect 23339 7497 23348 7531
rect 23296 7488 23348 7497
rect 12716 7420 12768 7429
rect 3148 7216 3200 7268
rect 7104 7284 7156 7336
rect 2964 7148 3016 7200
rect 5724 7191 5776 7200
rect 5724 7157 5733 7191
rect 5733 7157 5767 7191
rect 5767 7157 5776 7191
rect 5724 7148 5776 7157
rect 6184 7148 6236 7200
rect 9496 7352 9548 7404
rect 14280 7395 14332 7404
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 15292 7395 15344 7404
rect 15292 7361 15301 7395
rect 15301 7361 15335 7395
rect 15335 7361 15344 7395
rect 15292 7352 15344 7361
rect 16856 7463 16908 7472
rect 16856 7429 16865 7463
rect 16865 7429 16899 7463
rect 16899 7429 16908 7463
rect 22560 7463 22612 7472
rect 16856 7420 16908 7429
rect 8208 7284 8260 7336
rect 13820 7284 13872 7336
rect 14832 7284 14884 7336
rect 16948 7352 17000 7404
rect 17040 7395 17092 7404
rect 17040 7361 17049 7395
rect 17049 7361 17083 7395
rect 17083 7361 17092 7395
rect 17040 7352 17092 7361
rect 19340 7352 19392 7404
rect 15384 7216 15436 7268
rect 8208 7148 8260 7200
rect 8760 7148 8812 7200
rect 9220 7191 9272 7200
rect 9220 7157 9229 7191
rect 9229 7157 9263 7191
rect 9263 7157 9272 7191
rect 9220 7148 9272 7157
rect 9772 7191 9824 7200
rect 9772 7157 9781 7191
rect 9781 7157 9815 7191
rect 9815 7157 9824 7191
rect 9772 7148 9824 7157
rect 10416 7191 10468 7200
rect 10416 7157 10425 7191
rect 10425 7157 10459 7191
rect 10459 7157 10468 7191
rect 10416 7148 10468 7157
rect 11244 7148 11296 7200
rect 14280 7148 14332 7200
rect 14556 7148 14608 7200
rect 21364 7352 21416 7404
rect 22560 7429 22569 7463
rect 22569 7429 22603 7463
rect 22603 7429 22612 7463
rect 22560 7420 22612 7429
rect 23664 7463 23716 7472
rect 23664 7429 23673 7463
rect 23673 7429 23707 7463
rect 23707 7429 23716 7463
rect 23664 7420 23716 7429
rect 22652 7395 22704 7404
rect 22100 7284 22152 7336
rect 22652 7361 22661 7395
rect 22661 7361 22695 7395
rect 22695 7361 22704 7395
rect 22652 7352 22704 7361
rect 23388 7352 23440 7404
rect 24032 7352 24084 7404
rect 24768 7352 24820 7404
rect 31668 7488 31720 7540
rect 34612 7488 34664 7540
rect 34704 7420 34756 7472
rect 35624 7488 35676 7540
rect 36636 7488 36688 7540
rect 37096 7488 37148 7540
rect 39028 7488 39080 7540
rect 35532 7420 35584 7472
rect 25780 7395 25832 7404
rect 22744 7284 22796 7336
rect 23940 7284 23992 7336
rect 24308 7284 24360 7336
rect 25780 7361 25789 7395
rect 25789 7361 25823 7395
rect 25823 7361 25832 7395
rect 25780 7352 25832 7361
rect 25964 7395 26016 7404
rect 25964 7361 25973 7395
rect 25973 7361 26007 7395
rect 26007 7361 26016 7395
rect 25964 7352 26016 7361
rect 26884 7352 26936 7404
rect 25320 7327 25372 7336
rect 17040 7216 17092 7268
rect 18788 7216 18840 7268
rect 20076 7216 20128 7268
rect 25320 7293 25329 7327
rect 25329 7293 25363 7327
rect 25363 7293 25372 7327
rect 25320 7284 25372 7293
rect 26240 7284 26292 7336
rect 27804 7395 27856 7404
rect 27804 7361 27818 7395
rect 27818 7361 27852 7395
rect 27852 7361 27856 7395
rect 27804 7352 27856 7361
rect 27988 7395 28040 7404
rect 27988 7361 27997 7395
rect 27997 7361 28031 7395
rect 28031 7361 28040 7395
rect 27988 7352 28040 7361
rect 28172 7352 28224 7404
rect 30472 7395 30524 7404
rect 30472 7361 30506 7395
rect 30506 7361 30524 7395
rect 30472 7352 30524 7361
rect 34796 7352 34848 7404
rect 35256 7395 35308 7404
rect 35256 7361 35265 7395
rect 35265 7361 35299 7395
rect 35299 7361 35308 7395
rect 35256 7352 35308 7361
rect 29828 7284 29880 7336
rect 36176 7352 36228 7404
rect 37648 7352 37700 7404
rect 39672 7284 39724 7336
rect 18144 7191 18196 7200
rect 18144 7157 18153 7191
rect 18153 7157 18187 7191
rect 18187 7157 18196 7191
rect 18144 7148 18196 7157
rect 19064 7148 19116 7200
rect 27620 7216 27672 7268
rect 35348 7216 35400 7268
rect 27344 7191 27396 7200
rect 27344 7157 27353 7191
rect 27353 7157 27387 7191
rect 27387 7157 27396 7191
rect 27344 7148 27396 7157
rect 28632 7191 28684 7200
rect 28632 7157 28641 7191
rect 28641 7157 28675 7191
rect 28675 7157 28684 7191
rect 28632 7148 28684 7157
rect 38844 7148 38896 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3608 6944 3660 6996
rect 5356 6944 5408 6996
rect 6000 6987 6052 6996
rect 6000 6953 6009 6987
rect 6009 6953 6043 6987
rect 6043 6953 6052 6987
rect 6000 6944 6052 6953
rect 3976 6876 4028 6928
rect 5264 6876 5316 6928
rect 9496 6876 9548 6928
rect 14924 6876 14976 6928
rect 6092 6808 6144 6860
rect 2228 6783 2280 6792
rect 2228 6749 2237 6783
rect 2237 6749 2271 6783
rect 2271 6749 2280 6783
rect 2228 6740 2280 6749
rect 2504 6740 2556 6792
rect 2964 6740 3016 6792
rect 5264 6740 5316 6792
rect 6184 6783 6236 6792
rect 6184 6749 6193 6783
rect 6193 6749 6227 6783
rect 6227 6749 6236 6783
rect 6184 6740 6236 6749
rect 5816 6672 5868 6724
rect 2228 6604 2280 6656
rect 2964 6647 3016 6656
rect 2964 6613 2973 6647
rect 2973 6613 3007 6647
rect 3007 6613 3016 6647
rect 2964 6604 3016 6613
rect 4988 6647 5040 6656
rect 4988 6613 4997 6647
rect 4997 6613 5031 6647
rect 5031 6613 5040 6647
rect 4988 6604 5040 6613
rect 7380 6808 7432 6860
rect 7564 6740 7616 6792
rect 8760 6808 8812 6860
rect 13820 6808 13872 6860
rect 14004 6808 14056 6860
rect 8392 6740 8444 6792
rect 9220 6740 9272 6792
rect 11612 6783 11664 6792
rect 11612 6749 11630 6783
rect 11630 6749 11664 6783
rect 11612 6740 11664 6749
rect 14924 6740 14976 6792
rect 7104 6604 7156 6656
rect 8576 6672 8628 6724
rect 13084 6672 13136 6724
rect 15752 6715 15804 6724
rect 15752 6681 15761 6715
rect 15761 6681 15795 6715
rect 15795 6681 15804 6715
rect 15752 6672 15804 6681
rect 17040 6740 17092 6792
rect 18696 6851 18748 6860
rect 18696 6817 18705 6851
rect 18705 6817 18739 6851
rect 18739 6817 18748 6851
rect 18696 6808 18748 6817
rect 21272 6808 21324 6860
rect 16856 6672 16908 6724
rect 18512 6672 18564 6724
rect 18696 6672 18748 6724
rect 21732 6740 21784 6792
rect 22468 6740 22520 6792
rect 23480 6783 23532 6792
rect 23480 6749 23489 6783
rect 23489 6749 23523 6783
rect 23523 6749 23532 6783
rect 23480 6740 23532 6749
rect 23664 6783 23716 6792
rect 23664 6749 23673 6783
rect 23673 6749 23707 6783
rect 23707 6749 23716 6783
rect 23664 6740 23716 6749
rect 24032 6740 24084 6792
rect 24308 6740 24360 6792
rect 24584 6740 24636 6792
rect 8024 6604 8076 6656
rect 8944 6647 8996 6656
rect 8944 6613 8953 6647
rect 8953 6613 8987 6647
rect 8987 6613 8996 6647
rect 8944 6604 8996 6613
rect 10876 6604 10928 6656
rect 14740 6604 14792 6656
rect 15292 6604 15344 6656
rect 15568 6647 15620 6656
rect 15568 6613 15577 6647
rect 15577 6613 15611 6647
rect 15611 6613 15620 6647
rect 15568 6604 15620 6613
rect 16580 6647 16632 6656
rect 16580 6613 16589 6647
rect 16589 6613 16623 6647
rect 16623 6613 16632 6647
rect 16580 6604 16632 6613
rect 17408 6647 17460 6656
rect 17408 6613 17417 6647
rect 17417 6613 17451 6647
rect 17451 6613 17460 6647
rect 17408 6604 17460 6613
rect 19064 6604 19116 6656
rect 19984 6647 20036 6656
rect 19984 6613 19993 6647
rect 19993 6613 20027 6647
rect 20027 6613 20036 6647
rect 19984 6604 20036 6613
rect 20444 6647 20496 6656
rect 20444 6613 20453 6647
rect 20453 6613 20487 6647
rect 20487 6613 20496 6647
rect 20444 6604 20496 6613
rect 23204 6647 23256 6656
rect 23204 6613 23213 6647
rect 23213 6613 23247 6647
rect 23247 6613 23256 6647
rect 23204 6604 23256 6613
rect 23940 6672 23992 6724
rect 24860 6783 24912 6792
rect 24860 6749 24869 6783
rect 24869 6749 24903 6783
rect 24903 6749 24912 6783
rect 24860 6740 24912 6749
rect 26240 6783 26292 6792
rect 24308 6604 24360 6656
rect 24676 6604 24728 6656
rect 24768 6604 24820 6656
rect 26240 6749 26249 6783
rect 26249 6749 26283 6783
rect 26283 6749 26292 6783
rect 26240 6740 26292 6749
rect 27160 6740 27212 6792
rect 29828 6740 29880 6792
rect 30012 6783 30064 6792
rect 30012 6749 30021 6783
rect 30021 6749 30055 6783
rect 30055 6749 30064 6783
rect 30012 6740 30064 6749
rect 27344 6672 27396 6724
rect 29276 6604 29328 6656
rect 31208 6604 31260 6656
rect 32496 6740 32548 6792
rect 32680 6783 32732 6792
rect 32680 6749 32714 6783
rect 32714 6749 32732 6783
rect 32680 6740 32732 6749
rect 34336 6740 34388 6792
rect 35532 6783 35584 6792
rect 35532 6749 35541 6783
rect 35541 6749 35575 6783
rect 35575 6749 35584 6783
rect 35532 6740 35584 6749
rect 35900 6740 35952 6792
rect 36268 6740 36320 6792
rect 36636 6783 36688 6792
rect 36636 6749 36645 6783
rect 36645 6749 36679 6783
rect 36679 6749 36688 6783
rect 36636 6740 36688 6749
rect 36820 6783 36872 6792
rect 36820 6749 36829 6783
rect 36829 6749 36863 6783
rect 36863 6749 36872 6783
rect 36820 6740 36872 6749
rect 35808 6672 35860 6724
rect 37004 6783 37056 6792
rect 37004 6749 37013 6783
rect 37013 6749 37047 6783
rect 37047 6749 37056 6783
rect 37004 6740 37056 6749
rect 38844 6783 38896 6792
rect 38844 6749 38853 6783
rect 38853 6749 38887 6783
rect 38887 6749 38896 6783
rect 38844 6740 38896 6749
rect 39028 6783 39080 6792
rect 39028 6749 39037 6783
rect 39037 6749 39071 6783
rect 39071 6749 39080 6783
rect 39028 6740 39080 6749
rect 38936 6672 38988 6724
rect 31392 6604 31444 6656
rect 35440 6604 35492 6656
rect 37280 6647 37332 6656
rect 37280 6613 37289 6647
rect 37289 6613 37323 6647
rect 37323 6613 37332 6647
rect 37280 6604 37332 6613
rect 38384 6647 38436 6656
rect 38384 6613 38393 6647
rect 38393 6613 38427 6647
rect 38427 6613 38436 6647
rect 38384 6604 38436 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 3516 6400 3568 6452
rect 2964 6332 3016 6384
rect 6460 6332 6512 6384
rect 5448 6264 5500 6316
rect 2320 6239 2372 6248
rect 2320 6205 2329 6239
rect 2329 6205 2363 6239
rect 2363 6205 2372 6239
rect 2320 6196 2372 6205
rect 6000 6264 6052 6316
rect 3424 6128 3476 6180
rect 9220 6400 9272 6452
rect 16580 6400 16632 6452
rect 21272 6400 21324 6452
rect 24216 6400 24268 6452
rect 27804 6400 27856 6452
rect 29460 6400 29512 6452
rect 30104 6400 30156 6452
rect 30472 6400 30524 6452
rect 32496 6400 32548 6452
rect 35532 6400 35584 6452
rect 36820 6400 36872 6452
rect 6736 6332 6788 6384
rect 8484 6264 8536 6316
rect 15200 6332 15252 6384
rect 18788 6375 18840 6384
rect 18788 6341 18797 6375
rect 18797 6341 18831 6375
rect 18831 6341 18840 6375
rect 18788 6332 18840 6341
rect 20720 6332 20772 6384
rect 24768 6332 24820 6384
rect 26148 6332 26200 6384
rect 30012 6332 30064 6384
rect 34336 6375 34388 6384
rect 9036 6264 9088 6316
rect 9496 6264 9548 6316
rect 14740 6264 14792 6316
rect 16948 6307 17000 6316
rect 6828 6196 6880 6248
rect 7288 6196 7340 6248
rect 13268 6196 13320 6248
rect 16028 6239 16080 6248
rect 16028 6205 16037 6239
rect 16037 6205 16071 6239
rect 16071 6205 16080 6239
rect 16028 6196 16080 6205
rect 16580 6196 16632 6248
rect 16948 6273 16957 6307
rect 16957 6273 16991 6307
rect 16991 6273 17000 6307
rect 16948 6264 17000 6273
rect 18604 6307 18656 6316
rect 18604 6273 18613 6307
rect 18613 6273 18647 6307
rect 18647 6273 18656 6307
rect 18604 6264 18656 6273
rect 18144 6196 18196 6248
rect 18788 6196 18840 6248
rect 21732 6196 21784 6248
rect 23480 6307 23532 6316
rect 7012 6128 7064 6180
rect 10048 6128 10100 6180
rect 11060 6128 11112 6180
rect 13820 6128 13872 6180
rect 15752 6128 15804 6180
rect 22744 6196 22796 6248
rect 23480 6273 23489 6307
rect 23489 6273 23523 6307
rect 23523 6273 23532 6307
rect 23480 6264 23532 6273
rect 24584 6196 24636 6248
rect 26884 6196 26936 6248
rect 27988 6264 28040 6316
rect 28632 6307 28684 6316
rect 28632 6273 28641 6307
rect 28641 6273 28675 6307
rect 28675 6273 28684 6307
rect 28632 6264 28684 6273
rect 29276 6196 29328 6248
rect 30196 6264 30248 6316
rect 30288 6264 30340 6316
rect 30564 6307 30616 6316
rect 30564 6273 30573 6307
rect 30573 6273 30607 6307
rect 30607 6273 30616 6307
rect 30564 6264 30616 6273
rect 30656 6307 30708 6316
rect 30656 6273 30665 6307
rect 30665 6273 30699 6307
rect 30699 6273 30708 6307
rect 30656 6264 30708 6273
rect 31484 6196 31536 6248
rect 34336 6341 34345 6375
rect 34345 6341 34379 6375
rect 34379 6341 34388 6375
rect 34336 6332 34388 6341
rect 35808 6332 35860 6384
rect 37188 6332 37240 6384
rect 38752 6400 38804 6452
rect 39672 6443 39724 6452
rect 39672 6409 39681 6443
rect 39681 6409 39715 6443
rect 39715 6409 39724 6443
rect 39672 6400 39724 6409
rect 37648 6375 37700 6384
rect 37648 6341 37657 6375
rect 37657 6341 37691 6375
rect 37691 6341 37700 6375
rect 37648 6332 37700 6341
rect 38384 6332 38436 6384
rect 1860 6103 1912 6112
rect 1860 6069 1869 6103
rect 1869 6069 1903 6103
rect 1903 6069 1912 6103
rect 1860 6060 1912 6069
rect 5080 6103 5132 6112
rect 5080 6069 5089 6103
rect 5089 6069 5123 6103
rect 5123 6069 5132 6103
rect 5080 6060 5132 6069
rect 5632 6103 5684 6112
rect 5632 6069 5641 6103
rect 5641 6069 5675 6103
rect 5675 6069 5684 6103
rect 5632 6060 5684 6069
rect 6644 6103 6696 6112
rect 6644 6069 6653 6103
rect 6653 6069 6687 6103
rect 6687 6069 6696 6103
rect 6644 6060 6696 6069
rect 9956 6060 10008 6112
rect 10508 6060 10560 6112
rect 12164 6060 12216 6112
rect 15292 6060 15344 6112
rect 18144 6060 18196 6112
rect 19340 6060 19392 6112
rect 20168 6103 20220 6112
rect 20168 6069 20177 6103
rect 20177 6069 20211 6103
rect 20211 6069 20220 6103
rect 20168 6060 20220 6069
rect 20628 6103 20680 6112
rect 20628 6069 20637 6103
rect 20637 6069 20671 6103
rect 20671 6069 20680 6103
rect 20628 6060 20680 6069
rect 20720 6060 20772 6112
rect 21272 6060 21324 6112
rect 24952 6060 25004 6112
rect 30104 6060 30156 6112
rect 35348 6307 35400 6316
rect 35348 6273 35357 6307
rect 35357 6273 35391 6307
rect 35391 6273 35400 6307
rect 35348 6264 35400 6273
rect 35900 6264 35952 6316
rect 36176 6307 36228 6316
rect 36176 6273 36185 6307
rect 36185 6273 36219 6307
rect 36219 6273 36228 6307
rect 36176 6264 36228 6273
rect 34796 6196 34848 6248
rect 38292 6239 38344 6248
rect 38292 6205 38301 6239
rect 38301 6205 38335 6239
rect 38335 6205 38344 6239
rect 38292 6196 38344 6205
rect 37004 6128 37056 6180
rect 58164 6171 58216 6180
rect 58164 6137 58173 6171
rect 58173 6137 58207 6171
rect 58207 6137 58216 6171
rect 58164 6128 58216 6137
rect 35808 6060 35860 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 2320 5856 2372 5908
rect 6736 5856 6788 5908
rect 7748 5899 7800 5908
rect 7748 5865 7757 5899
rect 7757 5865 7791 5899
rect 7791 5865 7800 5899
rect 7748 5856 7800 5865
rect 13268 5856 13320 5908
rect 4988 5788 5040 5840
rect 9036 5788 9088 5840
rect 9220 5788 9272 5840
rect 15476 5856 15528 5908
rect 12992 5720 13044 5772
rect 15752 5856 15804 5908
rect 18604 5856 18656 5908
rect 2228 5695 2280 5704
rect 2228 5661 2237 5695
rect 2237 5661 2271 5695
rect 2271 5661 2280 5695
rect 2228 5652 2280 5661
rect 5816 5652 5868 5704
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 7012 5695 7064 5704
rect 7012 5661 7021 5695
rect 7021 5661 7055 5695
rect 7055 5661 7064 5695
rect 7012 5652 7064 5661
rect 7380 5652 7432 5704
rect 8852 5652 8904 5704
rect 9220 5652 9272 5704
rect 10232 5652 10284 5704
rect 10784 5652 10836 5704
rect 11336 5652 11388 5704
rect 11888 5652 11940 5704
rect 12440 5652 12492 5704
rect 12716 5652 12768 5704
rect 14832 5652 14884 5704
rect 16028 5652 16080 5704
rect 17316 5720 17368 5772
rect 17776 5788 17828 5840
rect 6828 5584 6880 5636
rect 13176 5584 13228 5636
rect 14556 5627 14608 5636
rect 14556 5593 14590 5627
rect 14590 5593 14608 5627
rect 14556 5584 14608 5593
rect 15384 5584 15436 5636
rect 16580 5695 16632 5704
rect 16580 5661 16589 5695
rect 16589 5661 16623 5695
rect 16623 5661 16632 5695
rect 16580 5652 16632 5661
rect 16764 5695 16816 5704
rect 16764 5661 16773 5695
rect 16773 5661 16807 5695
rect 16807 5661 16816 5695
rect 16764 5652 16816 5661
rect 16948 5652 17000 5704
rect 17868 5652 17920 5704
rect 18144 5695 18196 5704
rect 18144 5661 18153 5695
rect 18153 5661 18187 5695
rect 18187 5661 18196 5695
rect 18144 5652 18196 5661
rect 19248 5763 19300 5772
rect 19248 5729 19257 5763
rect 19257 5729 19291 5763
rect 19291 5729 19300 5763
rect 19248 5720 19300 5729
rect 23664 5856 23716 5908
rect 26148 5899 26200 5908
rect 26148 5865 26157 5899
rect 26157 5865 26191 5899
rect 26191 5865 26200 5899
rect 26148 5856 26200 5865
rect 26884 5899 26936 5908
rect 26884 5865 26893 5899
rect 26893 5865 26927 5899
rect 26927 5865 26936 5899
rect 26884 5856 26936 5865
rect 30288 5856 30340 5908
rect 32496 5856 32548 5908
rect 23756 5788 23808 5840
rect 24584 5788 24636 5840
rect 27436 5720 27488 5772
rect 18512 5584 18564 5636
rect 22744 5695 22796 5704
rect 22744 5661 22753 5695
rect 22753 5661 22787 5695
rect 22787 5661 22796 5695
rect 22744 5652 22796 5661
rect 23388 5652 23440 5704
rect 24768 5652 24820 5704
rect 25320 5695 25372 5704
rect 25320 5661 25329 5695
rect 25329 5661 25363 5695
rect 25363 5661 25372 5695
rect 25320 5652 25372 5661
rect 25780 5652 25832 5704
rect 1768 5559 1820 5568
rect 1768 5525 1777 5559
rect 1777 5525 1811 5559
rect 1811 5525 1820 5559
rect 1768 5516 1820 5525
rect 2504 5516 2556 5568
rect 6736 5559 6788 5568
rect 6736 5525 6745 5559
rect 6745 5525 6779 5559
rect 6779 5525 6788 5559
rect 6736 5516 6788 5525
rect 15292 5516 15344 5568
rect 15476 5516 15528 5568
rect 16120 5559 16172 5568
rect 16120 5525 16129 5559
rect 16129 5525 16163 5559
rect 16163 5525 16172 5559
rect 16120 5516 16172 5525
rect 17592 5516 17644 5568
rect 24584 5584 24636 5636
rect 21364 5559 21416 5568
rect 21364 5525 21373 5559
rect 21373 5525 21407 5559
rect 21407 5525 21416 5559
rect 21364 5516 21416 5525
rect 21916 5559 21968 5568
rect 21916 5525 21925 5559
rect 21925 5525 21959 5559
rect 21959 5525 21968 5559
rect 21916 5516 21968 5525
rect 23572 5516 23624 5568
rect 30104 5720 30156 5772
rect 28448 5652 28500 5704
rect 30196 5652 30248 5704
rect 34704 5831 34756 5840
rect 34704 5797 34713 5831
rect 34713 5797 34747 5831
rect 34747 5797 34756 5831
rect 34704 5788 34756 5797
rect 28632 5584 28684 5636
rect 30656 5695 30708 5704
rect 30656 5661 30685 5695
rect 30685 5661 30708 5695
rect 30656 5652 30708 5661
rect 32128 5652 32180 5704
rect 32404 5695 32456 5704
rect 32404 5661 32413 5695
rect 32413 5661 32447 5695
rect 32447 5661 32456 5695
rect 32404 5652 32456 5661
rect 35808 5695 35860 5704
rect 35808 5661 35826 5695
rect 35826 5661 35860 5695
rect 35808 5652 35860 5661
rect 27804 5516 27856 5568
rect 29552 5516 29604 5568
rect 30656 5516 30708 5568
rect 31484 5584 31536 5636
rect 35900 5584 35952 5636
rect 30932 5559 30984 5568
rect 30932 5525 30941 5559
rect 30941 5525 30975 5559
rect 30975 5525 30984 5559
rect 30932 5516 30984 5525
rect 37372 5516 37424 5568
rect 38292 5516 38344 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 3792 5312 3844 5364
rect 5080 5312 5132 5364
rect 2320 5176 2372 5228
rect 2504 5219 2556 5228
rect 2504 5185 2538 5219
rect 2538 5185 2556 5219
rect 2504 5176 2556 5185
rect 5172 5244 5224 5296
rect 6368 5287 6420 5296
rect 6368 5253 6377 5287
rect 6377 5253 6411 5287
rect 6411 5253 6420 5287
rect 6368 5244 6420 5253
rect 4896 5176 4948 5228
rect 5356 5176 5408 5228
rect 3792 5108 3844 5160
rect 6000 5176 6052 5228
rect 8852 5312 8904 5364
rect 9220 5355 9272 5364
rect 9220 5321 9229 5355
rect 9229 5321 9263 5355
rect 9263 5321 9272 5355
rect 9220 5312 9272 5321
rect 14188 5312 14240 5364
rect 14556 5355 14608 5364
rect 14556 5321 14565 5355
rect 14565 5321 14599 5355
rect 14599 5321 14608 5355
rect 14556 5312 14608 5321
rect 6736 5244 6788 5296
rect 7012 5176 7064 5228
rect 7656 5219 7708 5228
rect 7656 5185 7665 5219
rect 7665 5185 7699 5219
rect 7699 5185 7708 5219
rect 7656 5176 7708 5185
rect 7840 5176 7892 5228
rect 11428 5176 11480 5228
rect 6552 5108 6604 5160
rect 6276 5040 6328 5092
rect 11796 5108 11848 5160
rect 10140 5040 10192 5092
rect 11152 5040 11204 5092
rect 11704 5040 11756 5092
rect 14004 5176 14056 5228
rect 15384 5312 15436 5364
rect 16580 5312 16632 5364
rect 24860 5312 24912 5364
rect 15568 5244 15620 5296
rect 17040 5244 17092 5296
rect 16764 5176 16816 5228
rect 17592 5176 17644 5228
rect 17868 5176 17920 5228
rect 19340 5244 19392 5296
rect 20076 5244 20128 5296
rect 21548 5244 21600 5296
rect 24584 5287 24636 5296
rect 24584 5253 24593 5287
rect 24593 5253 24627 5287
rect 24627 5253 24636 5287
rect 24584 5244 24636 5253
rect 26240 5244 26292 5296
rect 30564 5312 30616 5364
rect 38752 5355 38804 5364
rect 38752 5321 38761 5355
rect 38761 5321 38795 5355
rect 38795 5321 38804 5355
rect 38752 5312 38804 5321
rect 18512 5219 18564 5228
rect 18512 5185 18521 5219
rect 18521 5185 18555 5219
rect 18555 5185 18564 5219
rect 18512 5176 18564 5185
rect 18788 5176 18840 5228
rect 25320 5176 25372 5228
rect 26332 5176 26384 5228
rect 26516 5176 26568 5228
rect 27804 5176 27856 5228
rect 27988 5176 28040 5228
rect 30196 5219 30248 5228
rect 30196 5185 30205 5219
rect 30205 5185 30239 5219
rect 30239 5185 30248 5219
rect 30196 5176 30248 5185
rect 30288 5176 30340 5228
rect 37280 5244 37332 5296
rect 37372 5219 37424 5228
rect 22192 5108 22244 5160
rect 29644 5151 29696 5160
rect 29644 5117 29653 5151
rect 29653 5117 29687 5151
rect 29687 5117 29696 5151
rect 37372 5185 37381 5219
rect 37381 5185 37415 5219
rect 37415 5185 37424 5219
rect 37372 5176 37424 5185
rect 29644 5108 29696 5117
rect 53748 5108 53800 5160
rect 22652 5040 22704 5092
rect 54116 5040 54168 5092
rect 4896 4972 4948 5024
rect 4988 5015 5040 5024
rect 4988 4981 4997 5015
rect 4997 4981 5031 5015
rect 5031 4981 5040 5015
rect 5724 5015 5776 5024
rect 4988 4972 5040 4981
rect 5724 4981 5733 5015
rect 5733 4981 5767 5015
rect 5767 4981 5776 5015
rect 5724 4972 5776 4981
rect 6460 4972 6512 5024
rect 7748 4972 7800 5024
rect 8024 5015 8076 5024
rect 8024 4981 8033 5015
rect 8033 4981 8067 5015
rect 8067 4981 8076 5015
rect 8024 4972 8076 4981
rect 11612 4972 11664 5024
rect 11980 4972 12032 5024
rect 13544 4972 13596 5024
rect 14372 4972 14424 5024
rect 15384 4972 15436 5024
rect 17592 5015 17644 5024
rect 17592 4981 17601 5015
rect 17601 4981 17635 5015
rect 17635 4981 17644 5015
rect 17592 4972 17644 4981
rect 18880 5015 18932 5024
rect 18880 4981 18889 5015
rect 18889 4981 18923 5015
rect 18923 4981 18932 5015
rect 18880 4972 18932 4981
rect 19340 5015 19392 5024
rect 19340 4981 19349 5015
rect 19349 4981 19383 5015
rect 19383 4981 19392 5015
rect 19340 4972 19392 4981
rect 20076 4972 20128 5024
rect 20904 4972 20956 5024
rect 21824 5015 21876 5024
rect 21824 4981 21833 5015
rect 21833 4981 21867 5015
rect 21867 4981 21876 5015
rect 21824 4972 21876 4981
rect 22284 4972 22336 5024
rect 26332 5015 26384 5024
rect 26332 4981 26341 5015
rect 26341 4981 26375 5015
rect 26375 4981 26384 5015
rect 26332 4972 26384 4981
rect 27252 5015 27304 5024
rect 27252 4981 27261 5015
rect 27261 4981 27295 5015
rect 27295 4981 27304 5015
rect 27252 4972 27304 4981
rect 30840 5015 30892 5024
rect 30840 4981 30849 5015
rect 30849 4981 30883 5015
rect 30883 4981 30892 5015
rect 30840 4972 30892 4981
rect 53656 4972 53708 5024
rect 58164 5015 58216 5024
rect 58164 4981 58173 5015
rect 58173 4981 58207 5015
rect 58207 4981 58216 5015
rect 58164 4972 58216 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 6000 4768 6052 4820
rect 6736 4768 6788 4820
rect 7656 4768 7708 4820
rect 8668 4768 8720 4820
rect 10048 4768 10100 4820
rect 10324 4811 10376 4820
rect 10324 4777 10333 4811
rect 10333 4777 10367 4811
rect 10367 4777 10376 4811
rect 10324 4768 10376 4777
rect 10968 4811 11020 4820
rect 10968 4777 10977 4811
rect 10977 4777 11011 4811
rect 11011 4777 11020 4811
rect 10968 4768 11020 4777
rect 3976 4700 4028 4752
rect 7012 4700 7064 4752
rect 7748 4700 7800 4752
rect 1768 4632 1820 4684
rect 4160 4632 4212 4684
rect 5080 4632 5132 4684
rect 2504 4564 2556 4616
rect 3056 4607 3108 4616
rect 3056 4573 3065 4607
rect 3065 4573 3099 4607
rect 3099 4573 3108 4607
rect 3056 4564 3108 4573
rect 4620 4564 4672 4616
rect 5264 4564 5316 4616
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 6276 4564 6328 4616
rect 9864 4675 9916 4684
rect 9864 4641 9870 4675
rect 9870 4641 9916 4675
rect 9864 4632 9916 4641
rect 11704 4768 11756 4820
rect 11428 4743 11480 4752
rect 11428 4709 11437 4743
rect 11437 4709 11471 4743
rect 11471 4709 11480 4743
rect 11428 4700 11480 4709
rect 16488 4700 16540 4752
rect 18972 4700 19024 4752
rect 20812 4768 20864 4820
rect 24584 4768 24636 4820
rect 28448 4768 28500 4820
rect 32404 4768 32456 4820
rect 21732 4700 21784 4752
rect 52184 4700 52236 4752
rect 53932 4700 53984 4752
rect 11520 4632 11572 4684
rect 12256 4632 12308 4684
rect 6644 4607 6696 4616
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 7104 4564 7156 4616
rect 3976 4496 4028 4548
rect 4160 4496 4212 4548
rect 6736 4496 6788 4548
rect 7932 4564 7984 4616
rect 9128 4564 9180 4616
rect 7840 4496 7892 4548
rect 11428 4564 11480 4616
rect 11796 4607 11848 4616
rect 11796 4573 11805 4607
rect 11805 4573 11839 4607
rect 11839 4573 11848 4607
rect 11796 4564 11848 4573
rect 16028 4632 16080 4684
rect 27160 4675 27212 4684
rect 27160 4641 27169 4675
rect 27169 4641 27203 4675
rect 27203 4641 27212 4675
rect 27160 4632 27212 4641
rect 31208 4675 31260 4684
rect 31208 4641 31217 4675
rect 31217 4641 31251 4675
rect 31251 4641 31260 4675
rect 31208 4632 31260 4641
rect 53196 4632 53248 4684
rect 54300 4632 54352 4684
rect 3700 4428 3752 4480
rect 4620 4428 4672 4480
rect 7104 4428 7156 4480
rect 7288 4428 7340 4480
rect 10140 4496 10192 4548
rect 14004 4564 14056 4616
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 14740 4564 14792 4616
rect 15936 4564 15988 4616
rect 16764 4564 16816 4616
rect 18604 4564 18656 4616
rect 18880 4564 18932 4616
rect 21732 4607 21784 4616
rect 21732 4573 21741 4607
rect 21741 4573 21775 4607
rect 21775 4573 21784 4607
rect 21732 4564 21784 4573
rect 22560 4564 22612 4616
rect 23112 4564 23164 4616
rect 23480 4607 23532 4616
rect 23480 4573 23489 4607
rect 23489 4573 23523 4607
rect 23523 4573 23532 4607
rect 23480 4564 23532 4573
rect 23940 4564 23992 4616
rect 24952 4564 25004 4616
rect 27252 4564 27304 4616
rect 30932 4564 30984 4616
rect 52092 4564 52144 4616
rect 52644 4564 52696 4616
rect 18144 4496 18196 4548
rect 24676 4539 24728 4548
rect 24676 4505 24710 4539
rect 24710 4505 24728 4539
rect 24676 4496 24728 4505
rect 8300 4428 8352 4480
rect 10048 4428 10100 4480
rect 11520 4428 11572 4480
rect 11980 4428 12032 4480
rect 14832 4428 14884 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 3056 4267 3108 4276
rect 3056 4233 3065 4267
rect 3065 4233 3099 4267
rect 3099 4233 3108 4267
rect 3056 4224 3108 4233
rect 3700 4224 3752 4276
rect 5540 4224 5592 4276
rect 6276 4224 6328 4276
rect 6552 4267 6604 4276
rect 6552 4233 6577 4267
rect 6577 4233 6604 4267
rect 6552 4224 6604 4233
rect 7104 4224 7156 4276
rect 7472 4224 7524 4276
rect 7656 4224 7708 4276
rect 3608 4156 3660 4208
rect 2688 4088 2740 4140
rect 3148 4088 3200 4140
rect 3884 4088 3936 4140
rect 4896 4156 4948 4208
rect 4896 4020 4948 4072
rect 7932 4088 7984 4140
rect 5816 4020 5868 4072
rect 6552 4020 6604 4072
rect 7472 4063 7524 4072
rect 7472 4029 7481 4063
rect 7481 4029 7515 4063
rect 7515 4029 7524 4063
rect 7472 4020 7524 4029
rect 7840 4020 7892 4072
rect 3700 3952 3752 4004
rect 3976 3952 4028 4004
rect 1952 3927 2004 3936
rect 1952 3893 1961 3927
rect 1961 3893 1995 3927
rect 1995 3893 2004 3927
rect 1952 3884 2004 3893
rect 6460 3884 6512 3936
rect 6920 3952 6972 4004
rect 7104 3884 7156 3936
rect 9312 4088 9364 4140
rect 9772 4088 9824 4140
rect 15568 4224 15620 4276
rect 15844 4224 15896 4276
rect 22100 4156 22152 4208
rect 8484 4020 8536 4072
rect 8668 4063 8720 4072
rect 8668 4029 8677 4063
rect 8677 4029 8711 4063
rect 8711 4029 8720 4063
rect 8668 4020 8720 4029
rect 11428 4020 11480 4072
rect 11704 4020 11756 4072
rect 12900 4020 12952 4072
rect 14648 4020 14700 4072
rect 15752 4088 15804 4140
rect 16672 4088 16724 4140
rect 17224 4088 17276 4140
rect 23204 4088 23256 4140
rect 35900 4156 35952 4208
rect 35440 4131 35492 4140
rect 35440 4097 35474 4131
rect 35474 4097 35492 4131
rect 35440 4088 35492 4097
rect 53012 4088 53064 4140
rect 17868 4020 17920 4072
rect 8760 3952 8812 4004
rect 9496 3995 9548 4004
rect 9496 3961 9505 3995
rect 9505 3961 9539 3995
rect 9539 3961 9548 3995
rect 9496 3952 9548 3961
rect 9864 3952 9916 4004
rect 11980 3995 12032 4004
rect 8944 3884 8996 3936
rect 9220 3884 9272 3936
rect 10600 3884 10652 3936
rect 11980 3961 11989 3995
rect 11989 3961 12023 3995
rect 12023 3961 12032 3995
rect 11980 3952 12032 3961
rect 15292 3952 15344 4004
rect 15844 3995 15896 4004
rect 15844 3961 15853 3995
rect 15853 3961 15887 3995
rect 15887 3961 15896 3995
rect 15844 3952 15896 3961
rect 19432 3952 19484 4004
rect 21456 3952 21508 4004
rect 11796 3884 11848 3936
rect 16304 3884 16356 3936
rect 17316 3884 17368 3936
rect 18788 3884 18840 3936
rect 19708 3884 19760 3936
rect 20352 3884 20404 3936
rect 22008 3884 22060 3936
rect 22468 3884 22520 3936
rect 24032 4020 24084 4072
rect 51816 4020 51868 4072
rect 54024 4020 54076 4072
rect 23940 3884 23992 3936
rect 24768 3952 24820 4004
rect 36176 3952 36228 4004
rect 52828 3952 52880 4004
rect 25688 3927 25740 3936
rect 25688 3893 25697 3927
rect 25697 3893 25731 3927
rect 25731 3893 25740 3927
rect 25688 3884 25740 3893
rect 26240 3927 26292 3936
rect 26240 3893 26249 3927
rect 26249 3893 26283 3927
rect 26283 3893 26292 3927
rect 26240 3884 26292 3893
rect 51080 3884 51132 3936
rect 51356 3884 51408 3936
rect 52460 3884 52512 3936
rect 55312 3927 55364 3936
rect 55312 3893 55321 3927
rect 55321 3893 55355 3927
rect 55355 3893 55364 3927
rect 55312 3884 55364 3893
rect 58440 3884 58492 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 3700 3680 3752 3732
rect 4896 3680 4948 3732
rect 4988 3680 5040 3732
rect 6276 3680 6328 3732
rect 6368 3680 6420 3732
rect 7472 3680 7524 3732
rect 9864 3680 9916 3732
rect 17684 3680 17736 3732
rect 20260 3723 20312 3732
rect 20260 3689 20269 3723
rect 20269 3689 20303 3723
rect 20303 3689 20312 3723
rect 20260 3680 20312 3689
rect 20996 3723 21048 3732
rect 20996 3689 21005 3723
rect 21005 3689 21039 3723
rect 21039 3689 21048 3723
rect 20996 3680 21048 3689
rect 21088 3680 21140 3732
rect 25688 3680 25740 3732
rect 32128 3723 32180 3732
rect 32128 3689 32137 3723
rect 32137 3689 32171 3723
rect 32171 3689 32180 3723
rect 32128 3680 32180 3689
rect 52736 3680 52788 3732
rect 8208 3655 8260 3664
rect 2412 3476 2464 3528
rect 6092 3544 6144 3596
rect 6368 3544 6420 3596
rect 8208 3621 8217 3655
rect 8217 3621 8251 3655
rect 8251 3621 8260 3655
rect 8208 3612 8260 3621
rect 9404 3655 9456 3664
rect 9404 3621 9413 3655
rect 9413 3621 9447 3655
rect 9447 3621 9456 3655
rect 9404 3612 9456 3621
rect 9680 3612 9732 3664
rect 11060 3544 11112 3596
rect 5356 3476 5408 3528
rect 9036 3476 9088 3528
rect 9496 3476 9548 3528
rect 9772 3476 9824 3528
rect 10692 3476 10744 3528
rect 11244 3476 11296 3528
rect 14188 3544 14240 3596
rect 12072 3519 12124 3528
rect 12072 3485 12081 3519
rect 12081 3485 12115 3519
rect 12115 3485 12124 3519
rect 12072 3476 12124 3485
rect 13268 3476 13320 3528
rect 13360 3519 13412 3528
rect 13360 3485 13369 3519
rect 13369 3485 13403 3519
rect 13403 3485 13412 3519
rect 13360 3476 13412 3485
rect 13636 3476 13688 3528
rect 19156 3612 19208 3664
rect 19248 3612 19300 3664
rect 26240 3612 26292 3664
rect 46296 3612 46348 3664
rect 51448 3612 51500 3664
rect 16028 3587 16080 3596
rect 16028 3553 16037 3587
rect 16037 3553 16071 3587
rect 16071 3553 16080 3587
rect 16028 3544 16080 3553
rect 21180 3544 21232 3596
rect 21548 3544 21600 3596
rect 50804 3544 50856 3596
rect 51632 3544 51684 3596
rect 53840 3544 53892 3596
rect 2596 3408 2648 3460
rect 4712 3408 4764 3460
rect 5172 3408 5224 3460
rect 6092 3408 6144 3460
rect 9128 3408 9180 3460
rect 4068 3340 4120 3392
rect 14832 3451 14884 3460
rect 14832 3417 14841 3451
rect 14841 3417 14875 3451
rect 14875 3417 14884 3451
rect 14832 3408 14884 3417
rect 16120 3476 16172 3528
rect 17408 3476 17460 3528
rect 18328 3476 18380 3528
rect 20168 3519 20220 3528
rect 20168 3485 20177 3519
rect 20177 3485 20211 3519
rect 20211 3485 20220 3519
rect 20168 3476 20220 3485
rect 21640 3476 21692 3528
rect 21824 3476 21876 3528
rect 23664 3476 23716 3528
rect 24216 3476 24268 3528
rect 24768 3476 24820 3528
rect 25596 3476 25648 3528
rect 26700 3476 26752 3528
rect 27528 3476 27580 3528
rect 28632 3476 28684 3528
rect 34704 3476 34756 3528
rect 35348 3476 35400 3528
rect 35808 3476 35860 3528
rect 36636 3476 36688 3528
rect 37464 3476 37516 3528
rect 38568 3476 38620 3528
rect 39948 3476 40000 3528
rect 40500 3476 40552 3528
rect 41052 3476 41104 3528
rect 42432 3476 42484 3528
rect 42708 3476 42760 3528
rect 44364 3476 44416 3528
rect 45192 3476 45244 3528
rect 46020 3476 46072 3528
rect 47676 3476 47728 3528
rect 48228 3476 48280 3528
rect 50160 3476 50212 3528
rect 50620 3476 50672 3528
rect 51172 3476 51224 3528
rect 52276 3476 52328 3528
rect 14096 3383 14148 3392
rect 14096 3349 14105 3383
rect 14105 3349 14139 3383
rect 14139 3349 14148 3383
rect 14096 3340 14148 3349
rect 15752 3340 15804 3392
rect 16028 3340 16080 3392
rect 20812 3408 20864 3460
rect 30840 3408 30892 3460
rect 31208 3408 31260 3460
rect 53288 3408 53340 3460
rect 57520 3519 57572 3528
rect 57520 3485 57529 3519
rect 57529 3485 57563 3519
rect 57563 3485 57572 3519
rect 57520 3476 57572 3485
rect 58164 3519 58216 3528
rect 58164 3485 58173 3519
rect 58173 3485 58207 3519
rect 58207 3485 58216 3519
rect 58164 3476 58216 3485
rect 18880 3340 18932 3392
rect 19708 3340 19760 3392
rect 20168 3340 20220 3392
rect 22836 3340 22888 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 3424 3136 3476 3188
rect 3792 3179 3844 3188
rect 3792 3145 3801 3179
rect 3801 3145 3835 3179
rect 3835 3145 3844 3179
rect 3792 3136 3844 3145
rect 3884 3136 3936 3188
rect 5356 3136 5408 3188
rect 8208 3136 8260 3188
rect 1952 3068 2004 3120
rect 4620 3068 4672 3120
rect 1492 3000 1544 3052
rect 2412 3043 2464 3052
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2412 3000 2464 3009
rect 5080 3000 5132 3052
rect 5264 2932 5316 2984
rect 6828 3000 6880 3052
rect 7288 3000 7340 3052
rect 7932 3000 7984 3052
rect 8208 3000 8260 3052
rect 9772 3136 9824 3188
rect 13636 3136 13688 3188
rect 14556 3179 14608 3188
rect 14556 3145 14565 3179
rect 14565 3145 14599 3179
rect 14599 3145 14608 3179
rect 14556 3136 14608 3145
rect 15200 3179 15252 3188
rect 15200 3145 15209 3179
rect 15209 3145 15243 3179
rect 15243 3145 15252 3179
rect 15200 3136 15252 3145
rect 16120 3136 16172 3188
rect 17408 3179 17460 3188
rect 17408 3145 17417 3179
rect 17417 3145 17451 3179
rect 17451 3145 17460 3179
rect 17408 3136 17460 3145
rect 8576 3068 8628 3120
rect 8852 3068 8904 3120
rect 10416 3111 10468 3120
rect 5816 2907 5868 2916
rect 2688 2796 2740 2848
rect 5816 2873 5825 2907
rect 5825 2873 5859 2907
rect 5859 2873 5868 2907
rect 5816 2864 5868 2873
rect 7656 2932 7708 2984
rect 7748 2932 7800 2984
rect 7840 2864 7892 2916
rect 8484 2932 8536 2984
rect 8668 3000 8720 3052
rect 8944 3043 8996 3052
rect 8944 3009 8953 3043
rect 8953 3009 8987 3043
rect 8987 3009 8996 3043
rect 8944 3000 8996 3009
rect 10416 3077 10425 3111
rect 10425 3077 10459 3111
rect 10459 3077 10468 3111
rect 10416 3068 10468 3077
rect 9864 3043 9916 3052
rect 9864 3009 9873 3043
rect 9873 3009 9907 3043
rect 9907 3009 9916 3043
rect 9864 3000 9916 3009
rect 10968 3000 11020 3052
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 17040 3068 17092 3120
rect 13084 3000 13136 3052
rect 14464 3000 14516 3052
rect 4896 2796 4948 2848
rect 5632 2839 5684 2848
rect 5632 2805 5641 2839
rect 5641 2805 5675 2839
rect 5675 2805 5684 2839
rect 5632 2796 5684 2805
rect 7472 2796 7524 2848
rect 7932 2796 7984 2848
rect 9036 2864 9088 2916
rect 9220 2796 9272 2848
rect 9404 2864 9456 2916
rect 11060 2864 11112 2916
rect 15016 2932 15068 2984
rect 15660 3000 15712 3052
rect 16396 3000 16448 3052
rect 16948 3000 17000 3052
rect 17776 3136 17828 3188
rect 21088 3136 21140 3188
rect 23020 3179 23072 3188
rect 23020 3145 23029 3179
rect 23029 3145 23063 3179
rect 23063 3145 23072 3179
rect 23020 3136 23072 3145
rect 18052 3111 18104 3120
rect 18052 3077 18061 3111
rect 18061 3077 18095 3111
rect 18095 3077 18104 3111
rect 18052 3068 18104 3077
rect 18788 3111 18840 3120
rect 18788 3077 18797 3111
rect 18797 3077 18831 3111
rect 18831 3077 18840 3111
rect 18788 3068 18840 3077
rect 19064 3068 19116 3120
rect 20628 3068 20680 3120
rect 20996 3111 21048 3120
rect 18512 3000 18564 3052
rect 18696 3000 18748 3052
rect 19984 3000 20036 3052
rect 15568 2932 15620 2984
rect 12072 2864 12124 2916
rect 14464 2864 14516 2916
rect 19064 2932 19116 2984
rect 19248 2932 19300 2984
rect 19616 2932 19668 2984
rect 20352 2932 20404 2984
rect 20628 2932 20680 2984
rect 16396 2864 16448 2916
rect 19432 2864 19484 2916
rect 19892 2864 19944 2916
rect 10416 2796 10468 2848
rect 15108 2796 15160 2848
rect 16672 2796 16724 2848
rect 18420 2796 18472 2848
rect 19800 2796 19852 2848
rect 20536 2796 20588 2848
rect 20996 3077 21005 3111
rect 21005 3077 21039 3111
rect 21039 3077 21048 3111
rect 20996 3068 21048 3077
rect 21364 3068 21416 3120
rect 22192 3111 22244 3120
rect 22192 3077 22201 3111
rect 22201 3077 22235 3111
rect 22235 3077 22244 3111
rect 22192 3068 22244 3077
rect 22376 3111 22428 3120
rect 22376 3077 22385 3111
rect 22385 3077 22419 3111
rect 22419 3077 22428 3111
rect 22376 3068 22428 3077
rect 51908 3068 51960 3120
rect 22836 3043 22888 3052
rect 22836 3009 22845 3043
rect 22845 3009 22879 3043
rect 22879 3009 22888 3043
rect 22836 3000 22888 3009
rect 51724 3000 51776 3052
rect 54760 3000 54812 3052
rect 24492 2932 24544 2984
rect 32772 2932 32824 2984
rect 38292 2932 38344 2984
rect 42156 2932 42208 2984
rect 53104 2932 53156 2984
rect 56600 2975 56652 2984
rect 56600 2941 56609 2975
rect 56609 2941 56643 2975
rect 56643 2941 56652 2975
rect 56600 2932 56652 2941
rect 33876 2864 33928 2916
rect 37188 2864 37240 2916
rect 39120 2864 39172 2916
rect 40224 2864 40276 2916
rect 42984 2864 43036 2916
rect 44088 2864 44140 2916
rect 22468 2796 22520 2848
rect 22836 2796 22888 2848
rect 25044 2796 25096 2848
rect 25320 2796 25372 2848
rect 26148 2796 26200 2848
rect 26976 2796 27028 2848
rect 27804 2796 27856 2848
rect 28080 2839 28132 2848
rect 28080 2805 28089 2839
rect 28089 2805 28123 2839
rect 28123 2805 28132 2839
rect 28080 2796 28132 2805
rect 29184 2796 29236 2848
rect 29736 2796 29788 2848
rect 30012 2839 30064 2848
rect 30012 2805 30021 2839
rect 30021 2805 30055 2839
rect 30055 2805 30064 2839
rect 30012 2796 30064 2805
rect 30564 2796 30616 2848
rect 31668 2796 31720 2848
rect 32220 2796 32272 2848
rect 33324 2796 33376 2848
rect 34428 2796 34480 2848
rect 35440 2796 35492 2848
rect 36360 2796 36412 2848
rect 37740 2796 37792 2848
rect 39672 2796 39724 2848
rect 41604 2796 41656 2848
rect 43536 2796 43588 2848
rect 44916 2796 44968 2848
rect 47400 2864 47452 2916
rect 48780 2864 48832 2916
rect 49884 2864 49936 2916
rect 50988 2864 51040 2916
rect 54208 2864 54260 2916
rect 45468 2796 45520 2848
rect 46848 2796 46900 2848
rect 47952 2796 48004 2848
rect 49332 2796 49384 2848
rect 50712 2796 50764 2848
rect 51540 2796 51592 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 5172 2592 5224 2644
rect 5356 2592 5408 2644
rect 5632 2592 5684 2644
rect 6552 2592 6604 2644
rect 10416 2635 10468 2644
rect 10416 2601 10425 2635
rect 10425 2601 10459 2635
rect 10459 2601 10468 2635
rect 10416 2592 10468 2601
rect 11060 2592 11112 2644
rect 13452 2635 13504 2644
rect 13452 2601 13461 2635
rect 13461 2601 13495 2635
rect 13495 2601 13504 2635
rect 13452 2592 13504 2601
rect 14556 2635 14608 2644
rect 14556 2601 14565 2635
rect 14565 2601 14599 2635
rect 14599 2601 14608 2635
rect 14556 2592 14608 2601
rect 20352 2635 20404 2644
rect 20352 2601 20361 2635
rect 20361 2601 20395 2635
rect 20395 2601 20404 2635
rect 20352 2592 20404 2601
rect 22928 2592 22980 2644
rect 2044 2524 2096 2576
rect 7380 2524 7432 2576
rect 8576 2524 8628 2576
rect 16212 2524 16264 2576
rect 17500 2524 17552 2576
rect 17684 2567 17736 2576
rect 17684 2533 17693 2567
rect 17693 2533 17727 2567
rect 17727 2533 17736 2567
rect 17684 2524 17736 2533
rect 18788 2524 18840 2576
rect 21272 2567 21324 2576
rect 21272 2533 21281 2567
rect 21281 2533 21315 2567
rect 21315 2533 21324 2567
rect 21272 2524 21324 2533
rect 5264 2456 5316 2508
rect 6552 2456 6604 2508
rect 7932 2456 7984 2508
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 2596 2388 2648 2440
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 4804 2388 4856 2440
rect 5448 2388 5500 2440
rect 6184 2388 6236 2440
rect 7196 2388 7248 2440
rect 10968 2456 11020 2508
rect 9588 2388 9640 2440
rect 11520 2431 11572 2440
rect 11520 2397 11529 2431
rect 11529 2397 11563 2431
rect 11563 2397 11572 2431
rect 11520 2388 11572 2397
rect 13636 2456 13688 2508
rect 13176 2388 13228 2440
rect 13912 2388 13964 2440
rect 14556 2388 14608 2440
rect 15108 2431 15160 2440
rect 15108 2397 15117 2431
rect 15117 2397 15151 2431
rect 15151 2397 15160 2431
rect 15108 2388 15160 2397
rect 8116 2320 8168 2372
rect 8484 2320 8536 2372
rect 10416 2320 10468 2372
rect 22376 2456 22428 2508
rect 52000 2592 52052 2644
rect 26424 2524 26476 2576
rect 28356 2524 28408 2576
rect 34152 2524 34204 2576
rect 38016 2524 38068 2576
rect 41880 2524 41932 2576
rect 45744 2524 45796 2576
rect 49608 2524 49660 2576
rect 31944 2456 31996 2508
rect 33048 2456 33100 2508
rect 35532 2456 35584 2508
rect 38844 2456 38896 2508
rect 40776 2456 40828 2508
rect 43260 2456 43312 2508
rect 46572 2456 46624 2508
rect 48504 2456 48556 2508
rect 16856 2388 16908 2440
rect 17500 2388 17552 2440
rect 19064 2388 19116 2440
rect 19432 2388 19484 2440
rect 22100 2388 22152 2440
rect 22652 2388 22704 2440
rect 23020 2388 23072 2440
rect 23296 2388 23348 2440
rect 25872 2388 25924 2440
rect 27252 2388 27304 2440
rect 17960 2320 18012 2372
rect 20352 2320 20404 2372
rect 20720 2320 20772 2372
rect 21916 2320 21968 2372
rect 28908 2388 28960 2440
rect 29460 2388 29512 2440
rect 30288 2388 30340 2440
rect 30840 2388 30892 2440
rect 31116 2388 31168 2440
rect 31392 2388 31444 2440
rect 32496 2388 32548 2440
rect 33600 2388 33652 2440
rect 36084 2388 36136 2440
rect 7748 2252 7800 2304
rect 8852 2252 8904 2304
rect 15292 2295 15344 2304
rect 15292 2261 15301 2295
rect 15301 2261 15335 2295
rect 15335 2261 15344 2295
rect 15292 2252 15344 2261
rect 17408 2252 17460 2304
rect 35716 2252 35768 2304
rect 36912 2320 36964 2372
rect 39396 2388 39448 2440
rect 41328 2388 41380 2440
rect 43812 2388 43864 2440
rect 44640 2320 44692 2372
rect 47124 2388 47176 2440
rect 49056 2388 49108 2440
rect 50896 2388 50948 2440
rect 57888 2499 57940 2508
rect 52552 2388 52604 2440
rect 46756 2252 46808 2304
rect 51264 2252 51316 2304
rect 57888 2465 57897 2499
rect 57897 2465 57931 2499
rect 57931 2465 57940 2499
rect 57888 2456 57940 2465
rect 55956 2431 56008 2440
rect 55956 2397 55965 2431
rect 55965 2397 55999 2431
rect 55999 2397 56008 2431
rect 55956 2388 56008 2397
rect 56600 2431 56652 2440
rect 56600 2397 56609 2431
rect 56609 2397 56643 2431
rect 56643 2397 56652 2431
rect 56600 2388 56652 2397
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 14556 2048 14608 2100
rect 16120 2048 16172 2100
rect 18880 2048 18932 2100
rect 19616 2048 19668 2100
rect 5448 1980 5500 2032
rect 10048 1980 10100 2032
rect 15292 1980 15344 2032
rect 25136 2048 25188 2100
rect 52368 2048 52420 2100
rect 55956 2048 56008 2100
rect 22468 1980 22520 2032
rect 22652 1980 22704 2032
rect 53564 1980 53616 2032
rect 57888 1980 57940 2032
rect 4068 1912 4120 1964
rect 11520 1912 11572 1964
rect 22376 1912 22428 1964
rect 29552 1912 29604 1964
rect 7932 1844 7984 1896
rect 8116 1844 8168 1896
rect 13176 1844 13228 1896
rect 15292 1844 15344 1896
rect 18880 1708 18932 1760
rect 19064 1708 19116 1760
rect 20720 1708 20772 1760
rect 21088 1708 21140 1760
rect 20260 1504 20312 1556
rect 1584 1436 1636 1488
rect 8116 1436 8168 1488
rect 15568 1300 15620 1352
rect 16028 1300 16080 1352
rect 19524 1300 19576 1352
rect 19800 1300 19852 1352
rect 19984 1300 20036 1352
rect 52736 1368 52788 1420
rect 53012 1368 53064 1420
rect 19432 1164 19484 1216
rect 20168 1028 20220 1080
rect 20352 1028 20404 1080
rect 52552 1096 52604 1148
rect 6184 892 6236 944
rect 6736 892 6788 944
rect 19432 892 19484 944
rect 50988 892 51040 944
rect 52552 892 52604 944
rect 52920 892 52972 944
rect 56600 1368 56652 1420
rect 54760 824 54812 876
<< metal2 >>
rect 1766 59200 1822 60000
rect 3330 59200 3386 60000
rect 4894 59200 4950 60000
rect 6458 59200 6514 60000
rect 8022 59200 8078 60000
rect 9586 59200 9642 60000
rect 11150 59200 11206 60000
rect 12714 59200 12770 60000
rect 14278 59200 14334 60000
rect 15842 59200 15898 60000
rect 17406 59200 17462 60000
rect 18970 59200 19026 60000
rect 19076 59214 19288 59242
rect 1780 57594 1808 59200
rect 3344 57594 3372 59200
rect 4908 57594 4936 59200
rect 6472 57594 6500 59200
rect 8036 57594 8064 59200
rect 1768 57588 1820 57594
rect 1768 57530 1820 57536
rect 3332 57588 3384 57594
rect 3332 57530 3384 57536
rect 4896 57588 4948 57594
rect 4896 57530 4948 57536
rect 6460 57588 6512 57594
rect 6460 57530 6512 57536
rect 8024 57588 8076 57594
rect 9600 57576 9628 59200
rect 11164 57594 11192 59200
rect 12728 57594 12756 59200
rect 14292 57594 14320 59200
rect 15856 57594 15884 59200
rect 17420 57594 17448 59200
rect 18984 59106 19012 59200
rect 19076 59106 19104 59214
rect 18984 59078 19104 59106
rect 19260 57610 19288 59214
rect 20534 59200 20590 60000
rect 22098 59200 22154 60000
rect 23662 59200 23718 60000
rect 25226 59200 25282 60000
rect 26790 59200 26846 60000
rect 28354 59200 28410 60000
rect 29918 59200 29974 60000
rect 31482 59200 31538 60000
rect 33046 59200 33102 60000
rect 34610 59200 34666 60000
rect 36174 59200 36230 60000
rect 37738 59200 37794 60000
rect 39302 59200 39358 60000
rect 40866 59200 40922 60000
rect 42430 59200 42486 60000
rect 43994 59200 44050 60000
rect 45558 59200 45614 60000
rect 47122 59200 47178 60000
rect 48686 59200 48742 60000
rect 50250 59200 50306 60000
rect 51814 59200 51870 60000
rect 53378 59200 53434 60000
rect 54942 59200 54998 60000
rect 56506 59200 56562 60000
rect 58070 59200 58126 60000
rect 58438 59256 58494 59265
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 20548 57610 20576 59200
rect 19260 57594 19380 57610
rect 20548 57594 20760 57610
rect 22112 57594 22140 59200
rect 23676 57594 23704 59200
rect 25240 57594 25268 59200
rect 26804 57594 26832 59200
rect 28368 57594 28396 59200
rect 29932 57594 29960 59200
rect 31496 57594 31524 59200
rect 9680 57588 9732 57594
rect 9600 57548 9680 57576
rect 8024 57530 8076 57536
rect 9680 57530 9732 57536
rect 11152 57588 11204 57594
rect 11152 57530 11204 57536
rect 12716 57588 12768 57594
rect 12716 57530 12768 57536
rect 14280 57588 14332 57594
rect 14280 57530 14332 57536
rect 15844 57588 15896 57594
rect 15844 57530 15896 57536
rect 17408 57588 17460 57594
rect 19260 57588 19392 57594
rect 19260 57582 19340 57588
rect 17408 57530 17460 57536
rect 20548 57588 20772 57594
rect 20548 57582 20720 57588
rect 19340 57530 19392 57536
rect 20720 57530 20772 57536
rect 22100 57588 22152 57594
rect 22100 57530 22152 57536
rect 23664 57588 23716 57594
rect 23664 57530 23716 57536
rect 25228 57588 25280 57594
rect 25228 57530 25280 57536
rect 26792 57588 26844 57594
rect 26792 57530 26844 57536
rect 28356 57588 28408 57594
rect 28356 57530 28408 57536
rect 29920 57588 29972 57594
rect 29920 57530 29972 57536
rect 31484 57588 31536 57594
rect 33060 57576 33088 59200
rect 34624 57594 34652 59200
rect 36188 57594 36216 59200
rect 37752 57594 37780 59200
rect 39316 57594 39344 59200
rect 40880 57594 40908 59200
rect 42444 57594 42472 59200
rect 33140 57588 33192 57594
rect 33060 57548 33140 57576
rect 31484 57530 31536 57536
rect 33140 57530 33192 57536
rect 34612 57588 34664 57594
rect 34612 57530 34664 57536
rect 36176 57588 36228 57594
rect 36176 57530 36228 57536
rect 37740 57588 37792 57594
rect 37740 57530 37792 57536
rect 39304 57588 39356 57594
rect 39304 57530 39356 57536
rect 40868 57588 40920 57594
rect 40868 57530 40920 57536
rect 42432 57588 42484 57594
rect 44008 57576 44036 59200
rect 45572 57594 45600 59200
rect 47136 57594 47164 59200
rect 44180 57588 44232 57594
rect 44008 57548 44180 57576
rect 42432 57530 42484 57536
rect 44180 57530 44232 57536
rect 45560 57588 45612 57594
rect 45560 57530 45612 57536
rect 47124 57588 47176 57594
rect 47124 57530 47176 57536
rect 26332 57520 26384 57526
rect 26332 57462 26384 57468
rect 30380 57520 30432 57526
rect 30380 57462 30432 57468
rect 2688 57452 2740 57458
rect 2688 57394 2740 57400
rect 4068 57452 4120 57458
rect 4068 57394 4120 57400
rect 5264 57452 5316 57458
rect 5264 57394 5316 57400
rect 6828 57452 6880 57458
rect 6828 57394 6880 57400
rect 11796 57452 11848 57458
rect 11796 57394 11848 57400
rect 13084 57452 13136 57458
rect 13084 57394 13136 57400
rect 15752 57452 15804 57458
rect 15752 57394 15804 57400
rect 16948 57452 17000 57458
rect 16948 57394 17000 57400
rect 17500 57452 17552 57458
rect 17500 57394 17552 57400
rect 18696 57452 18748 57458
rect 18696 57394 18748 57400
rect 19524 57452 19576 57458
rect 19524 57394 19576 57400
rect 22192 57452 22244 57458
rect 22192 57394 22244 57400
rect 24400 57452 24452 57458
rect 24400 57394 24452 57400
rect 25320 57452 25372 57458
rect 25320 57394 25372 57400
rect 2700 57254 2728 57394
rect 2688 57248 2740 57254
rect 2688 57190 2740 57196
rect 1400 56840 1452 56846
rect 1400 56782 1452 56788
rect 1412 56681 1440 56782
rect 1398 56672 1454 56681
rect 1398 56607 1454 56616
rect 2700 55962 2728 57190
rect 4080 56234 4108 57394
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 5276 56302 5304 57394
rect 6840 56982 6868 57394
rect 6828 56976 6880 56982
rect 6828 56918 6880 56924
rect 11808 56914 11836 57394
rect 11796 56908 11848 56914
rect 11796 56850 11848 56856
rect 13096 56506 13124 57394
rect 15764 56506 15792 57394
rect 13084 56500 13136 56506
rect 13084 56442 13136 56448
rect 15752 56500 15804 56506
rect 15752 56442 15804 56448
rect 14188 56364 14240 56370
rect 14188 56306 14240 56312
rect 15936 56364 15988 56370
rect 15936 56306 15988 56312
rect 5264 56296 5316 56302
rect 5264 56238 5316 56244
rect 4068 56228 4120 56234
rect 4068 56170 4120 56176
rect 14200 56166 14228 56306
rect 14188 56160 14240 56166
rect 14186 56128 14188 56137
rect 14240 56128 14242 56137
rect 4214 56060 4522 56069
rect 14186 56063 14242 56072
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 2688 55956 2740 55962
rect 2688 55898 2740 55904
rect 1400 55752 1452 55758
rect 1400 55694 1452 55700
rect 1412 55593 1440 55694
rect 15948 55622 15976 56306
rect 16960 55894 16988 57394
rect 17512 56506 17540 57394
rect 18512 57316 18564 57322
rect 18512 57258 18564 57264
rect 18144 56840 18196 56846
rect 18144 56782 18196 56788
rect 17500 56500 17552 56506
rect 17500 56442 17552 56448
rect 17684 56364 17736 56370
rect 17684 56306 17736 56312
rect 16948 55888 17000 55894
rect 16948 55830 17000 55836
rect 15936 55616 15988 55622
rect 1398 55584 1454 55593
rect 15936 55558 15988 55564
rect 16488 55616 16540 55622
rect 17040 55616 17092 55622
rect 16488 55558 16540 55564
rect 17038 55584 17040 55593
rect 17696 55593 17724 56306
rect 17776 55752 17828 55758
rect 17776 55694 17828 55700
rect 17092 55584 17094 55593
rect 1398 55519 1454 55528
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 1400 54664 1452 54670
rect 1400 54606 1452 54612
rect 1412 54505 1440 54606
rect 1398 54496 1454 54505
rect 1398 54431 1454 54440
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 1400 53576 1452 53582
rect 1400 53518 1452 53524
rect 1412 53417 1440 53518
rect 1398 53408 1454 53417
rect 1398 53343 1454 53352
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 1400 52488 1452 52494
rect 1400 52430 1452 52436
rect 1412 52329 1440 52430
rect 1398 52320 1454 52329
rect 1398 52255 1454 52264
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 1400 51400 1452 51406
rect 1400 51342 1452 51348
rect 1412 51241 1440 51342
rect 1398 51232 1454 51241
rect 1398 51167 1454 51176
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 16212 50380 16264 50386
rect 16212 50322 16264 50328
rect 1400 50312 1452 50318
rect 1400 50254 1452 50260
rect 1412 50153 1440 50254
rect 1398 50144 1454 50153
rect 1398 50079 1454 50088
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 1400 49224 1452 49230
rect 1400 49166 1452 49172
rect 1412 49065 1440 49166
rect 1398 49056 1454 49065
rect 1398 48991 1454 49000
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 1400 48136 1452 48142
rect 1400 48078 1452 48084
rect 1412 47977 1440 48078
rect 1398 47968 1454 47977
rect 1398 47903 1454 47912
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 13636 44872 13688 44878
rect 13636 44814 13688 44820
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 12440 41540 12492 41546
rect 12440 41482 12492 41488
rect 12992 41540 13044 41546
rect 12992 41482 13044 41488
rect 9864 41472 9916 41478
rect 9864 41414 9916 41420
rect 6552 41200 6604 41206
rect 6552 41142 6604 41148
rect 6368 40928 6420 40934
rect 6368 40870 6420 40876
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 6380 40526 6408 40870
rect 6092 40520 6144 40526
rect 6092 40462 6144 40468
rect 6368 40520 6420 40526
rect 6368 40462 6420 40468
rect 3976 40452 4028 40458
rect 3976 40394 4028 40400
rect 3988 40186 4016 40394
rect 4620 40384 4672 40390
rect 4620 40326 4672 40332
rect 3516 40180 3568 40186
rect 3516 40122 3568 40128
rect 3976 40180 4028 40186
rect 3976 40122 4028 40128
rect 2596 39976 2648 39982
rect 2596 39918 2648 39924
rect 2608 39506 2636 39918
rect 2596 39500 2648 39506
rect 2596 39442 2648 39448
rect 2608 38978 2636 39442
rect 2516 38962 2636 38978
rect 2504 38956 2636 38962
rect 2556 38950 2636 38956
rect 2504 38898 2556 38904
rect 2136 38208 2188 38214
rect 2136 38150 2188 38156
rect 2148 37194 2176 38150
rect 2608 37262 2636 38950
rect 2872 38344 2924 38350
rect 2872 38286 2924 38292
rect 3056 38344 3108 38350
rect 3056 38286 3108 38292
rect 2884 37670 2912 38286
rect 3068 38010 3096 38286
rect 3424 38208 3476 38214
rect 3424 38150 3476 38156
rect 3056 38004 3108 38010
rect 3056 37946 3108 37952
rect 3436 37942 3464 38150
rect 3424 37936 3476 37942
rect 3424 37878 3476 37884
rect 3240 37868 3292 37874
rect 3240 37810 3292 37816
rect 2872 37664 2924 37670
rect 2872 37606 2924 37612
rect 2596 37256 2648 37262
rect 2596 37198 2648 37204
rect 2136 37188 2188 37194
rect 2136 37130 2188 37136
rect 2608 36854 2636 37198
rect 3252 37126 3280 37810
rect 3240 37120 3292 37126
rect 3240 37062 3292 37068
rect 2596 36848 2648 36854
rect 2596 36790 2648 36796
rect 2608 36242 2636 36790
rect 2596 36236 2648 36242
rect 2596 36178 2648 36184
rect 2608 34610 2636 36178
rect 2872 35692 2924 35698
rect 2872 35634 2924 35640
rect 2688 35012 2740 35018
rect 2688 34954 2740 34960
rect 2596 34604 2648 34610
rect 2596 34546 2648 34552
rect 2608 33522 2636 34546
rect 2596 33516 2648 33522
rect 2596 33458 2648 33464
rect 2136 32428 2188 32434
rect 2136 32370 2188 32376
rect 1860 32360 1912 32366
rect 1860 32302 1912 32308
rect 1872 30802 1900 32302
rect 2148 32026 2176 32370
rect 2136 32020 2188 32026
rect 2136 31962 2188 31968
rect 2320 31816 2372 31822
rect 2320 31758 2372 31764
rect 2596 31816 2648 31822
rect 2596 31758 2648 31764
rect 2332 31142 2360 31758
rect 2608 31482 2636 31758
rect 2700 31754 2728 34954
rect 2780 31816 2832 31822
rect 2780 31758 2832 31764
rect 2688 31748 2740 31754
rect 2688 31690 2740 31696
rect 2596 31476 2648 31482
rect 2596 31418 2648 31424
rect 2320 31136 2372 31142
rect 2320 31078 2372 31084
rect 1860 30796 1912 30802
rect 1860 30738 1912 30744
rect 2136 30660 2188 30666
rect 2136 30602 2188 30608
rect 2148 30394 2176 30602
rect 2136 30388 2188 30394
rect 2136 30330 2188 30336
rect 2700 30122 2728 31690
rect 2792 30258 2820 31758
rect 2884 31346 2912 35634
rect 2872 31340 2924 31346
rect 2872 31282 2924 31288
rect 2872 30320 2924 30326
rect 2872 30262 2924 30268
rect 2780 30252 2832 30258
rect 2780 30194 2832 30200
rect 2688 30116 2740 30122
rect 2688 30058 2740 30064
rect 2700 29102 2728 30058
rect 2884 29850 2912 30262
rect 3148 30252 3200 30258
rect 3148 30194 3200 30200
rect 2872 29844 2924 29850
rect 2872 29786 2924 29792
rect 2688 29096 2740 29102
rect 2688 29038 2740 29044
rect 2504 28960 2556 28966
rect 2504 28902 2556 28908
rect 2516 28150 2544 28902
rect 2504 28144 2556 28150
rect 2504 28086 2556 28092
rect 2412 28008 2464 28014
rect 2412 27950 2464 27956
rect 2424 25906 2452 27950
rect 2412 25900 2464 25906
rect 2412 25842 2464 25848
rect 2424 24818 2452 25842
rect 2884 25294 2912 29786
rect 3160 29170 3188 30194
rect 3252 29714 3280 37062
rect 3332 31340 3384 31346
rect 3332 31282 3384 31288
rect 3344 30326 3372 31282
rect 3424 30592 3476 30598
rect 3424 30534 3476 30540
rect 3332 30320 3384 30326
rect 3332 30262 3384 30268
rect 3240 29708 3292 29714
rect 3240 29650 3292 29656
rect 2964 29164 3016 29170
rect 2964 29106 3016 29112
rect 3148 29164 3200 29170
rect 3148 29106 3200 29112
rect 2976 28762 3004 29106
rect 2964 28756 3016 28762
rect 2964 28698 3016 28704
rect 3344 28558 3372 30262
rect 3436 30258 3464 30534
rect 3424 30252 3476 30258
rect 3424 30194 3476 30200
rect 3436 29170 3464 30194
rect 3424 29164 3476 29170
rect 3424 29106 3476 29112
rect 3528 29034 3556 40122
rect 3792 40044 3844 40050
rect 3792 39986 3844 39992
rect 3804 39642 3832 39986
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 3792 39636 3844 39642
rect 3792 39578 3844 39584
rect 4632 39506 4660 40326
rect 6104 40118 6132 40462
rect 6368 40384 6420 40390
rect 6368 40326 6420 40332
rect 6092 40112 6144 40118
rect 6092 40054 6144 40060
rect 6380 40050 6408 40326
rect 6368 40044 6420 40050
rect 6368 39986 6420 39992
rect 5264 39568 5316 39574
rect 5264 39510 5316 39516
rect 4620 39500 4672 39506
rect 4620 39442 4672 39448
rect 4896 39432 4948 39438
rect 4896 39374 4948 39380
rect 4620 39364 4672 39370
rect 4620 39306 4672 39312
rect 4632 38962 4660 39306
rect 4908 38962 4936 39374
rect 5080 39024 5132 39030
rect 5080 38966 5132 38972
rect 4620 38956 4672 38962
rect 4620 38898 4672 38904
rect 4896 38956 4948 38962
rect 4896 38898 4948 38904
rect 4632 38758 4660 38898
rect 4712 38820 4764 38826
rect 4712 38762 4764 38768
rect 3976 38752 4028 38758
rect 3976 38694 4028 38700
rect 4620 38752 4672 38758
rect 4620 38694 4672 38700
rect 3988 38282 4016 38694
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4632 38418 4660 38694
rect 4724 38554 4752 38762
rect 4712 38548 4764 38554
rect 4712 38490 4764 38496
rect 4620 38412 4672 38418
rect 4620 38354 4672 38360
rect 4908 38350 4936 38898
rect 4896 38344 4948 38350
rect 4894 38312 4896 38321
rect 4948 38312 4950 38321
rect 3976 38276 4028 38282
rect 4894 38247 4950 38256
rect 3976 38218 4028 38224
rect 3792 33856 3844 33862
rect 3792 33798 3844 33804
rect 3804 33590 3832 33798
rect 3792 33584 3844 33590
rect 3792 33526 3844 33532
rect 3608 32224 3660 32230
rect 3608 32166 3660 32172
rect 3620 31278 3648 32166
rect 3608 31272 3660 31278
rect 3608 31214 3660 31220
rect 3620 29646 3648 31214
rect 3608 29640 3660 29646
rect 3608 29582 3660 29588
rect 3988 29238 4016 38218
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4620 36100 4672 36106
rect 4620 36042 4672 36048
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4632 35290 4660 36042
rect 4712 35488 4764 35494
rect 4712 35430 4764 35436
rect 4620 35284 4672 35290
rect 4620 35226 4672 35232
rect 4724 35086 4752 35430
rect 4988 35216 5040 35222
rect 4988 35158 5040 35164
rect 4712 35080 4764 35086
rect 4712 35022 4764 35028
rect 4620 34740 4672 34746
rect 4620 34682 4672 34688
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4632 33590 4660 34682
rect 4712 34468 4764 34474
rect 4712 34410 4764 34416
rect 4724 33658 4752 34410
rect 4896 34400 4948 34406
rect 4896 34342 4948 34348
rect 4908 34066 4936 34342
rect 4896 34060 4948 34066
rect 4896 34002 4948 34008
rect 4712 33652 4764 33658
rect 4712 33594 4764 33600
rect 4620 33584 4672 33590
rect 4620 33526 4672 33532
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4908 31754 4936 34002
rect 5000 33046 5028 35158
rect 5092 34134 5120 38966
rect 5172 36848 5224 36854
rect 5172 36790 5224 36796
rect 5184 36378 5212 36790
rect 5172 36372 5224 36378
rect 5172 36314 5224 36320
rect 5184 35766 5212 36314
rect 5172 35760 5224 35766
rect 5172 35702 5224 35708
rect 5080 34128 5132 34134
rect 5132 34076 5212 34082
rect 5080 34070 5212 34076
rect 5092 34054 5212 34070
rect 5080 33924 5132 33930
rect 5080 33866 5132 33872
rect 5092 33318 5120 33866
rect 5184 33658 5212 34054
rect 5172 33652 5224 33658
rect 5172 33594 5224 33600
rect 5080 33312 5132 33318
rect 5080 33254 5132 33260
rect 4988 33040 5040 33046
rect 4988 32982 5040 32988
rect 5000 31822 5028 32982
rect 4988 31816 5040 31822
rect 4988 31758 5040 31764
rect 4896 31748 4948 31754
rect 4896 31690 4948 31696
rect 4804 31680 4856 31686
rect 4804 31622 4856 31628
rect 4068 31136 4120 31142
rect 4068 31078 4120 31084
rect 3976 29232 4028 29238
rect 3976 29174 4028 29180
rect 3516 29028 3568 29034
rect 3516 28970 3568 28976
rect 3332 28552 3384 28558
rect 3332 28494 3384 28500
rect 3792 28484 3844 28490
rect 3792 28426 3844 28432
rect 3804 28218 3832 28426
rect 3792 28212 3844 28218
rect 3792 28154 3844 28160
rect 3608 28008 3660 28014
rect 3608 27950 3660 27956
rect 3056 27396 3108 27402
rect 3056 27338 3108 27344
rect 3068 26382 3096 27338
rect 3620 27062 3648 27950
rect 3608 27056 3660 27062
rect 3608 26998 3660 27004
rect 3240 26988 3292 26994
rect 3240 26930 3292 26936
rect 3252 26382 3280 26930
rect 3056 26376 3108 26382
rect 2976 26336 3056 26364
rect 2872 25288 2924 25294
rect 2872 25230 2924 25236
rect 2412 24812 2464 24818
rect 2412 24754 2464 24760
rect 1952 23724 2004 23730
rect 1952 23666 2004 23672
rect 1964 22710 1992 23666
rect 2320 22976 2372 22982
rect 2320 22918 2372 22924
rect 2332 22710 2360 22918
rect 1952 22704 2004 22710
rect 1952 22646 2004 22652
rect 2320 22704 2372 22710
rect 2320 22646 2372 22652
rect 2424 22642 2452 24754
rect 2976 24614 3004 26336
rect 3056 26318 3108 26324
rect 3240 26376 3292 26382
rect 3240 26318 3292 26324
rect 3620 26042 3648 26998
rect 3976 26784 4028 26790
rect 3976 26726 4028 26732
rect 3884 26444 3936 26450
rect 3884 26386 3936 26392
rect 3792 26240 3844 26246
rect 3792 26182 3844 26188
rect 3608 26036 3660 26042
rect 3608 25978 3660 25984
rect 3804 25974 3832 26182
rect 3792 25968 3844 25974
rect 3792 25910 3844 25916
rect 3896 25362 3924 26386
rect 3988 26314 4016 26726
rect 4080 26382 4108 31078
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4816 30666 4844 31622
rect 4804 30660 4856 30666
rect 4804 30602 4856 30608
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4712 29640 4764 29646
rect 4712 29582 4764 29588
rect 4620 29300 4672 29306
rect 4620 29242 4672 29248
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4632 26602 4660 29242
rect 4724 29238 4752 29582
rect 4804 29572 4856 29578
rect 4804 29514 4856 29520
rect 4712 29232 4764 29238
rect 4712 29174 4764 29180
rect 4816 29170 4844 29514
rect 4988 29504 5040 29510
rect 4988 29446 5040 29452
rect 4804 29164 4856 29170
rect 4804 29106 4856 29112
rect 4712 29028 4764 29034
rect 4712 28970 4764 28976
rect 4724 28558 4752 28970
rect 4712 28552 4764 28558
rect 4712 28494 4764 28500
rect 4816 28490 4844 29106
rect 4896 29028 4948 29034
rect 4896 28970 4948 28976
rect 4804 28484 4856 28490
rect 4804 28426 4856 28432
rect 4908 27470 4936 28970
rect 5000 28082 5028 29446
rect 4988 28076 5040 28082
rect 4988 28018 5040 28024
rect 5092 27606 5120 33254
rect 5184 29288 5212 33594
rect 5276 33114 5304 39510
rect 6092 39364 6144 39370
rect 6092 39306 6144 39312
rect 6104 38554 6132 39306
rect 6380 38962 6408 39986
rect 6368 38956 6420 38962
rect 6368 38898 6420 38904
rect 6092 38548 6144 38554
rect 6092 38490 6144 38496
rect 6380 38214 6408 38898
rect 6564 38758 6592 41142
rect 7656 41132 7708 41138
rect 7656 41074 7708 41080
rect 7104 41064 7156 41070
rect 7104 41006 7156 41012
rect 7116 40118 7144 41006
rect 7564 40928 7616 40934
rect 7564 40870 7616 40876
rect 7104 40112 7156 40118
rect 7104 40054 7156 40060
rect 7288 39432 7340 39438
rect 7288 39374 7340 39380
rect 6828 39296 6880 39302
rect 6828 39238 6880 39244
rect 6840 38962 6868 39238
rect 6828 38956 6880 38962
rect 6828 38898 6880 38904
rect 6552 38752 6604 38758
rect 6552 38694 6604 38700
rect 6644 38752 6696 38758
rect 6644 38694 6696 38700
rect 6460 38480 6512 38486
rect 6460 38422 6512 38428
rect 6472 38214 6500 38422
rect 6564 38264 6592 38694
rect 6656 38418 6684 38694
rect 6644 38412 6696 38418
rect 6644 38354 6696 38360
rect 6736 38344 6788 38350
rect 6734 38312 6736 38321
rect 6788 38312 6790 38321
rect 6644 38276 6696 38282
rect 6564 38236 6644 38264
rect 6734 38247 6790 38256
rect 6644 38218 6696 38224
rect 6368 38208 6420 38214
rect 6368 38150 6420 38156
rect 6460 38208 6512 38214
rect 6460 38150 6512 38156
rect 6380 38010 6408 38150
rect 6368 38004 6420 38010
rect 6368 37946 6420 37952
rect 5632 37664 5684 37670
rect 5632 37606 5684 37612
rect 5356 36236 5408 36242
rect 5356 36178 5408 36184
rect 5368 35018 5396 36178
rect 5356 35012 5408 35018
rect 5356 34954 5408 34960
rect 5644 34950 5672 37606
rect 6840 36854 6868 38898
rect 7300 38758 7328 39374
rect 7288 38752 7340 38758
rect 7288 38694 7340 38700
rect 7012 37188 7064 37194
rect 7012 37130 7064 37136
rect 6828 36848 6880 36854
rect 6828 36790 6880 36796
rect 7024 36378 7052 37130
rect 7104 36576 7156 36582
rect 7104 36518 7156 36524
rect 7012 36372 7064 36378
rect 7012 36314 7064 36320
rect 6644 36032 6696 36038
rect 6644 35974 6696 35980
rect 6092 35488 6144 35494
rect 6092 35430 6144 35436
rect 6552 35488 6604 35494
rect 6552 35430 6604 35436
rect 6104 35290 6132 35430
rect 6092 35284 6144 35290
rect 6092 35226 6144 35232
rect 5632 34944 5684 34950
rect 5632 34886 5684 34892
rect 5644 34746 5672 34886
rect 5632 34740 5684 34746
rect 5632 34682 5684 34688
rect 5448 34604 5500 34610
rect 5448 34546 5500 34552
rect 5460 34406 5488 34546
rect 5448 34400 5500 34406
rect 5448 34342 5500 34348
rect 5460 34202 5488 34342
rect 5448 34196 5500 34202
rect 5448 34138 5500 34144
rect 5460 33998 5488 34138
rect 5448 33992 5500 33998
rect 5448 33934 5500 33940
rect 5356 33584 5408 33590
rect 5356 33526 5408 33532
rect 5264 33108 5316 33114
rect 5264 33050 5316 33056
rect 5276 31958 5304 33050
rect 5264 31952 5316 31958
rect 5264 31894 5316 31900
rect 5264 31816 5316 31822
rect 5264 31758 5316 31764
rect 5276 31482 5304 31758
rect 5264 31476 5316 31482
rect 5264 31418 5316 31424
rect 5184 29260 5304 29288
rect 5172 29164 5224 29170
rect 5172 29106 5224 29112
rect 5184 28558 5212 29106
rect 5172 28552 5224 28558
rect 5172 28494 5224 28500
rect 5172 28008 5224 28014
rect 5172 27950 5224 27956
rect 5080 27600 5132 27606
rect 5080 27542 5132 27548
rect 5184 27470 5212 27950
rect 4896 27464 4948 27470
rect 4896 27406 4948 27412
rect 5172 27464 5224 27470
rect 5172 27406 5224 27412
rect 4632 26586 4752 26602
rect 4632 26580 4764 26586
rect 4632 26574 4712 26580
rect 4712 26522 4764 26528
rect 4620 26512 4672 26518
rect 4620 26454 4672 26460
rect 4724 26466 4752 26522
rect 4068 26376 4120 26382
rect 4120 26336 4200 26364
rect 4068 26318 4120 26324
rect 3976 26308 4028 26314
rect 3976 26250 4028 26256
rect 4172 25702 4200 26336
rect 4160 25696 4212 25702
rect 4160 25638 4212 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4632 25362 4660 26454
rect 4724 26438 4844 26466
rect 4712 26376 4764 26382
rect 4712 26318 4764 26324
rect 3884 25356 3936 25362
rect 3884 25298 3936 25304
rect 4620 25356 4672 25362
rect 4620 25298 4672 25304
rect 4724 25294 4752 26318
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 3608 25152 3660 25158
rect 3608 25094 3660 25100
rect 3620 24818 3648 25094
rect 4080 24818 4108 25230
rect 4724 24954 4752 25230
rect 4712 24948 4764 24954
rect 4712 24890 4764 24896
rect 3608 24812 3660 24818
rect 3608 24754 3660 24760
rect 4068 24812 4120 24818
rect 4068 24754 4120 24760
rect 3884 24744 3936 24750
rect 3884 24686 3936 24692
rect 2964 24608 3016 24614
rect 2964 24550 3016 24556
rect 3896 24410 3924 24686
rect 3884 24404 3936 24410
rect 3884 24346 3936 24352
rect 3240 23724 3292 23730
rect 3240 23666 3292 23672
rect 2688 23520 2740 23526
rect 2688 23462 2740 23468
rect 2596 22976 2648 22982
rect 2596 22918 2648 22924
rect 2412 22636 2464 22642
rect 2412 22578 2464 22584
rect 2608 22234 2636 22918
rect 2596 22228 2648 22234
rect 2596 22170 2648 22176
rect 2228 21956 2280 21962
rect 2228 21898 2280 21904
rect 2240 21690 2268 21898
rect 2608 21690 2636 22170
rect 2228 21684 2280 21690
rect 2228 21626 2280 21632
rect 2596 21684 2648 21690
rect 2596 21626 2648 21632
rect 2700 21554 2728 23462
rect 2780 23112 2832 23118
rect 2780 23054 2832 23060
rect 2964 23112 3016 23118
rect 2964 23054 3016 23060
rect 2792 22778 2820 23054
rect 2780 22772 2832 22778
rect 2780 22714 2832 22720
rect 2976 21554 3004 23054
rect 3252 21894 3280 23666
rect 3792 23656 3844 23662
rect 3792 23598 3844 23604
rect 3804 22710 3832 23598
rect 3792 22704 3844 22710
rect 3792 22646 3844 22652
rect 3240 21888 3292 21894
rect 3240 21830 3292 21836
rect 2504 21548 2556 21554
rect 2504 21490 2556 21496
rect 2688 21548 2740 21554
rect 2688 21490 2740 21496
rect 2964 21548 3016 21554
rect 2964 21490 3016 21496
rect 2516 20806 2544 21490
rect 3252 21486 3280 21830
rect 3804 21554 3832 22646
rect 3896 22030 3924 24346
rect 4080 23322 4108 24754
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4160 24132 4212 24138
rect 4160 24074 4212 24080
rect 4172 23866 4200 24074
rect 4160 23860 4212 23866
rect 4160 23802 4212 23808
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4816 23322 4844 26438
rect 4988 25696 5040 25702
rect 4988 25638 5040 25644
rect 4068 23316 4120 23322
rect 4068 23258 4120 23264
rect 4528 23316 4580 23322
rect 4528 23258 4580 23264
rect 4804 23316 4856 23322
rect 4804 23258 4856 23264
rect 3884 22024 3936 22030
rect 3884 21966 3936 21972
rect 3976 21888 4028 21894
rect 3976 21830 4028 21836
rect 3988 21622 4016 21830
rect 3976 21616 4028 21622
rect 3976 21558 4028 21564
rect 3792 21548 3844 21554
rect 3792 21490 3844 21496
rect 3240 21480 3292 21486
rect 3240 21422 3292 21428
rect 2504 20800 2556 20806
rect 2504 20742 2556 20748
rect 2412 19372 2464 19378
rect 2412 19314 2464 19320
rect 2136 19168 2188 19174
rect 2136 19110 2188 19116
rect 2148 18766 2176 19110
rect 1860 18760 1912 18766
rect 1860 18702 1912 18708
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 1676 18284 1728 18290
rect 1676 18226 1728 18232
rect 1688 17882 1716 18226
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1872 17270 1900 18702
rect 2424 18426 2452 19314
rect 4080 18698 4108 23258
rect 4540 22642 4568 23258
rect 4896 22976 4948 22982
rect 4896 22918 4948 22924
rect 4908 22642 4936 22918
rect 4528 22636 4580 22642
rect 4528 22578 4580 22584
rect 4712 22636 4764 22642
rect 4712 22578 4764 22584
rect 4896 22636 4948 22642
rect 4896 22578 4948 22584
rect 4620 22432 4672 22438
rect 4620 22374 4672 22380
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 21962 4660 22374
rect 4620 21956 4672 21962
rect 4620 21898 4672 21904
rect 4724 21690 4752 22578
rect 4712 21684 4764 21690
rect 4712 21626 4764 21632
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 5000 20806 5028 25638
rect 5276 24682 5304 29260
rect 5368 28150 5396 33526
rect 5460 32570 5488 33934
rect 5540 33924 5592 33930
rect 5540 33866 5592 33872
rect 5552 33522 5580 33866
rect 5540 33516 5592 33522
rect 5540 33458 5592 33464
rect 5552 32570 5580 33458
rect 5448 32564 5500 32570
rect 5448 32506 5500 32512
rect 5540 32564 5592 32570
rect 5540 32506 5592 32512
rect 5460 31958 5488 32506
rect 5448 31952 5500 31958
rect 5448 31894 5500 31900
rect 5552 31414 5580 32506
rect 5644 31657 5672 34682
rect 5724 32768 5776 32774
rect 5724 32710 5776 32716
rect 5630 31648 5686 31657
rect 5630 31583 5686 31592
rect 5540 31408 5592 31414
rect 5540 31350 5592 31356
rect 5632 31340 5684 31346
rect 5632 31282 5684 31288
rect 5644 30598 5672 31282
rect 5632 30592 5684 30598
rect 5632 30534 5684 30540
rect 5356 28144 5408 28150
rect 5356 28086 5408 28092
rect 5448 28076 5500 28082
rect 5448 28018 5500 28024
rect 5460 27470 5488 28018
rect 5448 27464 5500 27470
rect 5448 27406 5500 27412
rect 5632 27396 5684 27402
rect 5632 27338 5684 27344
rect 5448 26988 5500 26994
rect 5448 26930 5500 26936
rect 5460 26314 5488 26930
rect 5448 26308 5500 26314
rect 5448 26250 5500 26256
rect 5460 25974 5488 26250
rect 5644 25974 5672 27338
rect 5448 25968 5500 25974
rect 5448 25910 5500 25916
rect 5632 25968 5684 25974
rect 5632 25910 5684 25916
rect 5644 25498 5672 25910
rect 5632 25492 5684 25498
rect 5632 25434 5684 25440
rect 5264 24676 5316 24682
rect 5264 24618 5316 24624
rect 5080 23316 5132 23322
rect 5080 23258 5132 23264
rect 4988 20800 5040 20806
rect 4988 20742 5040 20748
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4804 19780 4856 19786
rect 4804 19722 4856 19728
rect 4620 19712 4672 19718
rect 4620 19654 4672 19660
rect 4632 19281 4660 19654
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4618 19272 4674 19281
rect 4618 19207 4674 19216
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 4068 18692 4120 18698
rect 4068 18634 4120 18640
rect 3332 18624 3384 18630
rect 4160 18624 4212 18630
rect 3332 18566 3384 18572
rect 4158 18592 4160 18601
rect 4212 18592 4214 18601
rect 2412 18420 2464 18426
rect 2412 18362 2464 18368
rect 3344 18290 3372 18566
rect 4158 18527 4214 18536
rect 4068 18352 4120 18358
rect 4068 18294 4120 18300
rect 3332 18284 3384 18290
rect 3332 18226 3384 18232
rect 2412 18216 2464 18222
rect 2412 18158 2464 18164
rect 3240 18216 3292 18222
rect 3240 18158 3292 18164
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1860 17264 1912 17270
rect 1860 17206 1912 17212
rect 1872 16658 1900 17206
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1964 16590 1992 18022
rect 2424 17678 2452 18158
rect 2412 17672 2464 17678
rect 2412 17614 2464 17620
rect 1952 16584 2004 16590
rect 1952 16526 2004 16532
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 2148 15706 2176 16050
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 2424 15502 2452 17614
rect 2780 17264 2832 17270
rect 2780 17206 2832 17212
rect 2504 15904 2556 15910
rect 2504 15846 2556 15852
rect 2596 15904 2648 15910
rect 2596 15846 2648 15852
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2424 14822 2452 15438
rect 2516 15026 2544 15846
rect 2608 15570 2636 15846
rect 2792 15570 2820 17206
rect 3252 16794 3280 18158
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 3344 17746 3372 18022
rect 4080 17882 4108 18294
rect 4632 18222 4660 18770
rect 4620 18216 4672 18222
rect 4620 18158 4672 18164
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 3332 17740 3384 17746
rect 3332 17682 3384 17688
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 3792 16176 3844 16182
rect 3792 16118 3844 16124
rect 2596 15564 2648 15570
rect 2596 15506 2648 15512
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 2792 15094 2820 15506
rect 3804 15366 3832 16118
rect 4632 16046 4660 18158
rect 4724 17678 4752 19314
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4252 15428 4304 15434
rect 4252 15370 4304 15376
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3804 15162 3832 15302
rect 4264 15162 4292 15370
rect 4724 15178 4752 17614
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4632 15150 4752 15178
rect 2780 15088 2832 15094
rect 2780 15030 2832 15036
rect 3240 15088 3292 15094
rect 3240 15030 3292 15036
rect 2504 15020 2556 15026
rect 2504 14962 2556 14968
rect 2412 14816 2464 14822
rect 2412 14758 2464 14764
rect 2424 13530 2452 14758
rect 2412 13524 2464 13530
rect 2412 13466 2464 13472
rect 2424 12782 2452 13466
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 2516 12238 2544 12582
rect 2792 12442 2820 12718
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2700 11830 2728 12038
rect 2688 11824 2740 11830
rect 2688 11766 2740 11772
rect 2792 11762 2820 12378
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 2056 10266 2084 10610
rect 2700 10606 2728 11086
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 2228 9988 2280 9994
rect 2228 9930 2280 9936
rect 2042 8664 2098 8673
rect 2042 8599 2098 8608
rect 1584 8356 1636 8362
rect 1584 8298 1636 8304
rect 1492 7744 1544 7750
rect 1492 7686 1544 7692
rect 1504 3058 1532 7686
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 1596 2446 1624 8298
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1872 5681 1900 6054
rect 1858 5672 1914 5681
rect 1858 5607 1914 5616
rect 1768 5568 1820 5574
rect 1768 5510 1820 5516
rect 1780 4690 1808 5510
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1964 3126 1992 3878
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 2056 2582 2084 8599
rect 2136 8356 2188 8362
rect 2136 8298 2188 8304
rect 2148 3097 2176 8298
rect 2240 7410 2268 9930
rect 2424 9654 2452 10406
rect 2700 9994 2728 10542
rect 2688 9988 2740 9994
rect 2688 9930 2740 9936
rect 2412 9648 2464 9654
rect 2412 9590 2464 9596
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2240 6798 2268 7346
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2240 5710 2268 6598
rect 2332 6254 2360 9318
rect 3252 8838 3280 15030
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 13530 4660 15150
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4724 14618 4752 14962
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4816 14498 4844 19722
rect 4896 19236 4948 19242
rect 4896 19178 4948 19184
rect 4908 18698 4936 19178
rect 4896 18692 4948 18698
rect 4896 18634 4948 18640
rect 4908 17814 4936 18634
rect 4896 17808 4948 17814
rect 4896 17750 4948 17756
rect 4896 17604 4948 17610
rect 5000 17592 5028 20742
rect 5092 17814 5120 23258
rect 5276 22094 5304 24618
rect 5736 23254 5764 32710
rect 5816 27872 5868 27878
rect 5816 27814 5868 27820
rect 5540 23248 5592 23254
rect 5540 23190 5592 23196
rect 5724 23248 5776 23254
rect 5724 23190 5776 23196
rect 5552 22574 5580 23190
rect 5736 22778 5764 23190
rect 5724 22772 5776 22778
rect 5724 22714 5776 22720
rect 5540 22568 5592 22574
rect 5540 22510 5592 22516
rect 5552 22234 5580 22510
rect 5540 22228 5592 22234
rect 5540 22170 5592 22176
rect 5276 22066 5488 22094
rect 5356 20528 5408 20534
rect 5356 20470 5408 20476
rect 5368 19718 5396 20470
rect 5356 19712 5408 19718
rect 5356 19654 5408 19660
rect 5368 19446 5396 19654
rect 5356 19440 5408 19446
rect 5356 19382 5408 19388
rect 5460 19174 5488 22066
rect 5632 21956 5684 21962
rect 5632 21898 5684 21904
rect 5644 21622 5672 21898
rect 5632 21616 5684 21622
rect 5632 21558 5684 21564
rect 5736 20058 5764 22714
rect 5828 22094 5856 27814
rect 6104 25906 6132 35226
rect 6564 35018 6592 35430
rect 6368 35012 6420 35018
rect 6368 34954 6420 34960
rect 6552 35012 6604 35018
rect 6552 34954 6604 34960
rect 6380 33930 6408 34954
rect 6564 34678 6592 34954
rect 6552 34672 6604 34678
rect 6552 34614 6604 34620
rect 6368 33924 6420 33930
rect 6368 33866 6420 33872
rect 6460 33652 6512 33658
rect 6460 33594 6512 33600
rect 6184 32020 6236 32026
rect 6184 31962 6236 31968
rect 6092 25900 6144 25906
rect 6092 25842 6144 25848
rect 6092 23112 6144 23118
rect 6092 23054 6144 23060
rect 5908 23044 5960 23050
rect 5908 22986 5960 22992
rect 5920 22778 5948 22986
rect 5908 22772 5960 22778
rect 5908 22714 5960 22720
rect 6000 22094 6052 22098
rect 6104 22094 6132 23054
rect 5828 22066 5948 22094
rect 5724 20052 5776 20058
rect 5724 19994 5776 20000
rect 5736 19514 5764 19994
rect 5724 19508 5776 19514
rect 5724 19450 5776 19456
rect 5632 19304 5684 19310
rect 5632 19246 5684 19252
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 5644 18970 5672 19246
rect 5632 18964 5684 18970
rect 5632 18906 5684 18912
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5552 18222 5580 18702
rect 5632 18624 5684 18630
rect 5632 18566 5684 18572
rect 5644 18358 5672 18566
rect 5632 18352 5684 18358
rect 5632 18294 5684 18300
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 5080 17808 5132 17814
rect 5080 17750 5132 17756
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 4948 17564 5028 17592
rect 4896 17546 4948 17552
rect 4908 16726 4936 17546
rect 4988 17196 5040 17202
rect 4988 17138 5040 17144
rect 5000 16794 5028 17138
rect 5184 16998 5212 17614
rect 5172 16992 5224 16998
rect 5172 16934 5224 16940
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 4896 16720 4948 16726
rect 4896 16662 4948 16668
rect 5080 15360 5132 15366
rect 5080 15302 5132 15308
rect 4724 14470 4844 14498
rect 4988 14544 5040 14550
rect 4988 14486 5040 14492
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3804 11354 3832 12786
rect 3896 12714 3924 13262
rect 4632 12850 4660 13466
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3896 11218 3924 12650
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 4632 10742 4660 12038
rect 4724 11694 4752 14470
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4816 11642 4844 12786
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4908 11762 4936 12038
rect 5000 11778 5028 14486
rect 5092 14482 5120 15302
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 5092 12986 5120 13262
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 5092 11898 5120 12922
rect 5184 12170 5212 16934
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5368 12782 5396 15982
rect 5644 15366 5672 18294
rect 5816 18148 5868 18154
rect 5816 18090 5868 18096
rect 5828 17882 5856 18090
rect 5816 17876 5868 17882
rect 5816 17818 5868 17824
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5644 14278 5672 15302
rect 5920 14822 5948 22066
rect 6000 22092 6132 22094
rect 6052 22066 6132 22092
rect 6000 22034 6052 22040
rect 6092 18216 6144 18222
rect 6092 18158 6144 18164
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 6012 16998 6040 17138
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 6012 16590 6040 16934
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 6012 15910 6040 16526
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5552 13870 5580 14214
rect 5540 13864 5592 13870
rect 5538 13832 5540 13841
rect 5592 13832 5594 13841
rect 5538 13767 5594 13776
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 5172 12164 5224 12170
rect 5172 12106 5224 12112
rect 5276 12102 5304 12582
rect 5368 12306 5396 12718
rect 5644 12434 5672 14214
rect 5552 12406 5672 12434
rect 6012 12434 6040 15846
rect 6104 15502 6132 18158
rect 6196 17882 6224 31962
rect 6368 28416 6420 28422
rect 6368 28358 6420 28364
rect 6380 28082 6408 28358
rect 6368 28076 6420 28082
rect 6368 28018 6420 28024
rect 6472 27470 6500 33594
rect 6656 32910 6684 35974
rect 6736 35012 6788 35018
rect 6736 34954 6788 34960
rect 6748 34066 6776 34954
rect 6736 34060 6788 34066
rect 6736 34002 6788 34008
rect 7116 33658 7144 36518
rect 7196 35692 7248 35698
rect 7196 35634 7248 35640
rect 7208 35290 7236 35634
rect 7196 35284 7248 35290
rect 7196 35226 7248 35232
rect 7104 33652 7156 33658
rect 7104 33594 7156 33600
rect 6920 33516 6972 33522
rect 6920 33458 6972 33464
rect 6932 33114 6960 33458
rect 7012 33312 7064 33318
rect 7012 33254 7064 33260
rect 6920 33108 6972 33114
rect 6920 33050 6972 33056
rect 6644 32904 6696 32910
rect 6644 32846 6696 32852
rect 6552 32360 6604 32366
rect 6552 32302 6604 32308
rect 6564 31686 6592 32302
rect 6828 32224 6880 32230
rect 6828 32166 6880 32172
rect 6552 31680 6604 31686
rect 6552 31622 6604 31628
rect 6564 31414 6592 31622
rect 6552 31408 6604 31414
rect 6552 31350 6604 31356
rect 6840 31346 6868 32166
rect 7024 32026 7052 33254
rect 7104 32428 7156 32434
rect 7104 32370 7156 32376
rect 7012 32020 7064 32026
rect 7012 31962 7064 31968
rect 7116 31754 7144 32370
rect 7024 31726 7144 31754
rect 6828 31340 6880 31346
rect 6828 31282 6880 31288
rect 6644 31136 6696 31142
rect 6644 31078 6696 31084
rect 6656 30666 6684 31078
rect 6644 30660 6696 30666
rect 6644 30602 6696 30608
rect 7024 30598 7052 31726
rect 6736 30592 6788 30598
rect 6736 30534 6788 30540
rect 7012 30592 7064 30598
rect 7012 30534 7064 30540
rect 6748 28150 6776 30534
rect 6736 28144 6788 28150
rect 6736 28086 6788 28092
rect 6552 28076 6604 28082
rect 6552 28018 6604 28024
rect 6564 27538 6592 28018
rect 6828 27940 6880 27946
rect 6828 27882 6880 27888
rect 6552 27532 6604 27538
rect 6552 27474 6604 27480
rect 6460 27464 6512 27470
rect 6460 27406 6512 27412
rect 6564 27130 6592 27474
rect 6840 27402 6868 27882
rect 7024 27470 7052 30534
rect 7104 28076 7156 28082
rect 7104 28018 7156 28024
rect 7116 27470 7144 28018
rect 7012 27464 7064 27470
rect 7012 27406 7064 27412
rect 7104 27464 7156 27470
rect 7104 27406 7156 27412
rect 6828 27396 6880 27402
rect 6828 27338 6880 27344
rect 6552 27124 6604 27130
rect 6552 27066 6604 27072
rect 6736 26376 6788 26382
rect 6736 26318 6788 26324
rect 6748 25909 6776 26318
rect 7012 26240 7064 26246
rect 7012 26182 7064 26188
rect 6552 25900 6604 25906
rect 6552 25842 6604 25848
rect 6705 25903 6776 25909
rect 7024 25906 7052 26182
rect 6757 25860 6776 25903
rect 7012 25900 7064 25906
rect 6705 25845 6757 25851
rect 7012 25842 7064 25848
rect 6460 25696 6512 25702
rect 6460 25638 6512 25644
rect 6472 25294 6500 25638
rect 6564 25498 6592 25842
rect 6552 25492 6604 25498
rect 6552 25434 6604 25440
rect 6460 25288 6512 25294
rect 6460 25230 6512 25236
rect 6564 24154 6592 25434
rect 7196 24608 7248 24614
rect 7196 24550 7248 24556
rect 7208 24206 7236 24550
rect 6472 24126 6592 24154
rect 6920 24200 6972 24206
rect 6920 24142 6972 24148
rect 7196 24200 7248 24206
rect 7196 24142 7248 24148
rect 6368 21956 6420 21962
rect 6368 21898 6420 21904
rect 6380 21690 6408 21898
rect 6472 21690 6500 24126
rect 6552 24064 6604 24070
rect 6552 24006 6604 24012
rect 6368 21684 6420 21690
rect 6368 21626 6420 21632
rect 6460 21684 6512 21690
rect 6460 21626 6512 21632
rect 6472 21554 6500 21626
rect 6460 21548 6512 21554
rect 6460 21490 6512 21496
rect 6184 17876 6236 17882
rect 6184 17818 6236 17824
rect 6564 17270 6592 24006
rect 6736 23656 6788 23662
rect 6736 23598 6788 23604
rect 6644 22568 6696 22574
rect 6748 22522 6776 23598
rect 6932 22982 6960 24142
rect 6920 22976 6972 22982
rect 6920 22918 6972 22924
rect 6696 22516 6776 22522
rect 6644 22510 6776 22516
rect 6656 22494 6776 22510
rect 6748 21554 6776 22494
rect 6932 22094 6960 22918
rect 7300 22094 7328 38694
rect 7472 37256 7524 37262
rect 7472 37198 7524 37204
rect 7484 36854 7512 37198
rect 7472 36848 7524 36854
rect 7472 36790 7524 36796
rect 7472 36576 7524 36582
rect 7472 36518 7524 36524
rect 7484 36174 7512 36518
rect 7472 36168 7524 36174
rect 7472 36110 7524 36116
rect 7576 35222 7604 40870
rect 7668 39438 7696 41074
rect 9876 40730 9904 41414
rect 11060 41200 11112 41206
rect 11060 41142 11112 41148
rect 10600 41132 10652 41138
rect 10600 41074 10652 41080
rect 10416 40928 10468 40934
rect 10416 40870 10468 40876
rect 9864 40724 9916 40730
rect 9864 40666 9916 40672
rect 9220 40588 9272 40594
rect 9220 40530 9272 40536
rect 7748 40384 7800 40390
rect 7748 40326 7800 40332
rect 7760 40186 7788 40326
rect 7748 40180 7800 40186
rect 7748 40122 7800 40128
rect 7656 39432 7708 39438
rect 7656 39374 7708 39380
rect 7668 38350 7696 39374
rect 7656 38344 7708 38350
rect 7656 38286 7708 38292
rect 7760 37262 7788 40122
rect 9232 40118 9260 40530
rect 9876 40526 9904 40666
rect 9864 40520 9916 40526
rect 9864 40462 9916 40468
rect 10048 40520 10100 40526
rect 10048 40462 10100 40468
rect 9588 40384 9640 40390
rect 9588 40326 9640 40332
rect 9600 40118 9628 40326
rect 9220 40112 9272 40118
rect 9220 40054 9272 40060
rect 9588 40112 9640 40118
rect 9588 40054 9640 40060
rect 9232 39982 9260 40054
rect 9220 39976 9272 39982
rect 9220 39918 9272 39924
rect 9232 39438 9260 39918
rect 9220 39432 9272 39438
rect 9220 39374 9272 39380
rect 8208 39296 8260 39302
rect 8208 39238 8260 39244
rect 8220 38894 8248 39238
rect 8208 38888 8260 38894
rect 8208 38830 8260 38836
rect 8024 38208 8076 38214
rect 8024 38150 8076 38156
rect 7748 37256 7800 37262
rect 7748 37198 7800 37204
rect 7840 37256 7892 37262
rect 7840 37198 7892 37204
rect 7656 37188 7708 37194
rect 7656 37130 7708 37136
rect 7668 36922 7696 37130
rect 7656 36916 7708 36922
rect 7656 36858 7708 36864
rect 7852 36786 7880 37198
rect 7840 36780 7892 36786
rect 7840 36722 7892 36728
rect 7932 36780 7984 36786
rect 7932 36722 7984 36728
rect 7944 35630 7972 36722
rect 7932 35624 7984 35630
rect 7932 35566 7984 35572
rect 7564 35216 7616 35222
rect 7564 35158 7616 35164
rect 7576 34610 7604 35158
rect 8036 34626 8064 38150
rect 7564 34604 7616 34610
rect 7564 34546 7616 34552
rect 7944 34598 8064 34626
rect 7576 34406 7604 34546
rect 7564 34400 7616 34406
rect 7564 34342 7616 34348
rect 7380 33856 7432 33862
rect 7380 33798 7432 33804
rect 7392 32910 7420 33798
rect 7380 32904 7432 32910
rect 7432 32852 7512 32858
rect 7380 32846 7512 32852
rect 7392 32830 7512 32846
rect 7380 31748 7432 31754
rect 7380 31690 7432 31696
rect 7392 31346 7420 31690
rect 7380 31340 7432 31346
rect 7380 31282 7432 31288
rect 7392 30394 7420 31282
rect 7380 30388 7432 30394
rect 7380 30330 7432 30336
rect 7484 26042 7512 32830
rect 7564 32836 7616 32842
rect 7564 32778 7616 32784
rect 7748 32836 7800 32842
rect 7748 32778 7800 32784
rect 7576 30326 7604 32778
rect 7760 32434 7788 32778
rect 7748 32428 7800 32434
rect 7748 32370 7800 32376
rect 7564 30320 7616 30326
rect 7564 30262 7616 30268
rect 7576 26382 7604 30262
rect 7760 27402 7788 32370
rect 7944 31278 7972 34598
rect 8024 34536 8076 34542
rect 8024 34478 8076 34484
rect 8036 33658 8064 34478
rect 8116 33856 8168 33862
rect 8116 33798 8168 33804
rect 8128 33658 8156 33798
rect 8024 33652 8076 33658
rect 8024 33594 8076 33600
rect 8116 33652 8168 33658
rect 8116 33594 8168 33600
rect 8036 32910 8064 33594
rect 8220 33538 8248 38830
rect 9232 38214 9260 39374
rect 9956 39364 10008 39370
rect 9956 39306 10008 39312
rect 9968 39098 9996 39306
rect 9956 39092 10008 39098
rect 9956 39034 10008 39040
rect 9312 38276 9364 38282
rect 9312 38218 9364 38224
rect 9220 38208 9272 38214
rect 9220 38150 9272 38156
rect 9324 37670 9352 38218
rect 10060 38010 10088 40462
rect 10140 40452 10192 40458
rect 10140 40394 10192 40400
rect 10152 39846 10180 40394
rect 10140 39840 10192 39846
rect 10140 39782 10192 39788
rect 10152 38826 10180 39782
rect 10428 38826 10456 40870
rect 10508 40520 10560 40526
rect 10508 40462 10560 40468
rect 10520 40050 10548 40462
rect 10508 40044 10560 40050
rect 10508 39986 10560 39992
rect 10508 39840 10560 39846
rect 10508 39782 10560 39788
rect 10140 38820 10192 38826
rect 10140 38762 10192 38768
rect 10416 38820 10468 38826
rect 10416 38762 10468 38768
rect 10048 38004 10100 38010
rect 10048 37946 10100 37952
rect 8300 37664 8352 37670
rect 8300 37606 8352 37612
rect 9312 37664 9364 37670
rect 9312 37606 9364 37612
rect 8312 36650 8340 37606
rect 10152 37274 10180 38762
rect 10232 38208 10284 38214
rect 10232 38150 10284 38156
rect 10060 37246 10180 37274
rect 8392 37120 8444 37126
rect 8392 37062 8444 37068
rect 8300 36644 8352 36650
rect 8300 36586 8352 36592
rect 8128 33510 8248 33538
rect 8024 32904 8076 32910
rect 8024 32846 8076 32852
rect 7932 31272 7984 31278
rect 7932 31214 7984 31220
rect 7944 30938 7972 31214
rect 7932 30932 7984 30938
rect 7932 30874 7984 30880
rect 8128 29850 8156 33510
rect 8208 32020 8260 32026
rect 8208 31962 8260 31968
rect 8220 31890 8248 31962
rect 8312 31958 8340 36586
rect 8404 34610 8432 37062
rect 9772 36780 9824 36786
rect 9772 36722 9824 36728
rect 9312 36168 9364 36174
rect 9312 36110 9364 36116
rect 9324 35630 9352 36110
rect 9496 36032 9548 36038
rect 9496 35974 9548 35980
rect 9312 35624 9364 35630
rect 9312 35566 9364 35572
rect 9128 34740 9180 34746
rect 9128 34682 9180 34688
rect 8392 34604 8444 34610
rect 8392 34546 8444 34552
rect 8668 34604 8720 34610
rect 8668 34546 8720 34552
rect 8392 33856 8444 33862
rect 8392 33798 8444 33804
rect 8300 31952 8352 31958
rect 8300 31894 8352 31900
rect 8208 31884 8260 31890
rect 8208 31826 8260 31832
rect 8220 30734 8248 31826
rect 8312 31521 8340 31894
rect 8298 31512 8354 31521
rect 8298 31447 8300 31456
rect 8352 31447 8354 31456
rect 8300 31418 8352 31424
rect 8208 30728 8260 30734
rect 8208 30670 8260 30676
rect 7932 29844 7984 29850
rect 7932 29786 7984 29792
rect 8116 29844 8168 29850
rect 8116 29786 8168 29792
rect 7944 29238 7972 29786
rect 8220 29714 8248 30670
rect 8208 29708 8260 29714
rect 8208 29650 8260 29656
rect 7932 29232 7984 29238
rect 7932 29174 7984 29180
rect 8208 29164 8260 29170
rect 8208 29106 8260 29112
rect 8220 28966 8248 29106
rect 8208 28960 8260 28966
rect 8208 28902 8260 28908
rect 8220 28014 8248 28902
rect 8208 28008 8260 28014
rect 8208 27950 8260 27956
rect 7840 27872 7892 27878
rect 7840 27814 7892 27820
rect 7748 27396 7800 27402
rect 7748 27338 7800 27344
rect 7564 26376 7616 26382
rect 7564 26318 7616 26324
rect 7760 26314 7788 27338
rect 7748 26308 7800 26314
rect 7748 26250 7800 26256
rect 7472 26036 7524 26042
rect 7472 25978 7524 25984
rect 7852 24954 7880 27814
rect 8208 27532 8260 27538
rect 8208 27474 8260 27480
rect 7932 27328 7984 27334
rect 7932 27270 7984 27276
rect 8116 27328 8168 27334
rect 8116 27270 8168 27276
rect 7944 27146 7972 27270
rect 7944 27118 8064 27146
rect 7932 26988 7984 26994
rect 7932 26930 7984 26936
rect 7944 26586 7972 26930
rect 7932 26580 7984 26586
rect 7932 26522 7984 26528
rect 7840 24948 7892 24954
rect 7840 24890 7892 24896
rect 7840 24404 7892 24410
rect 7840 24346 7892 24352
rect 7852 23730 7880 24346
rect 7840 23724 7892 23730
rect 7840 23666 7892 23672
rect 7840 23248 7892 23254
rect 7840 23190 7892 23196
rect 7852 22710 7880 23190
rect 7840 22704 7892 22710
rect 7840 22646 7892 22652
rect 6932 22066 7052 22094
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 6736 21548 6788 21554
rect 6736 21490 6788 21496
rect 6840 18970 6868 21626
rect 7024 21554 7052 22066
rect 7116 22066 7328 22094
rect 8036 22094 8064 27118
rect 8128 26518 8156 27270
rect 8220 26994 8248 27474
rect 8208 26988 8260 26994
rect 8208 26930 8260 26936
rect 8116 26512 8168 26518
rect 8116 26454 8168 26460
rect 8220 25362 8248 26930
rect 8312 26858 8340 31418
rect 8404 30326 8432 33798
rect 8680 33386 8708 34546
rect 8668 33380 8720 33386
rect 8668 33322 8720 33328
rect 8576 32360 8628 32366
rect 8576 32302 8628 32308
rect 8392 30320 8444 30326
rect 8392 30262 8444 30268
rect 8404 27334 8432 30262
rect 8588 28762 8616 32302
rect 8576 28756 8628 28762
rect 8576 28698 8628 28704
rect 8588 28218 8616 28698
rect 8576 28212 8628 28218
rect 8576 28154 8628 28160
rect 8484 27600 8536 27606
rect 8484 27542 8536 27548
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8300 26852 8352 26858
rect 8300 26794 8352 26800
rect 8392 26376 8444 26382
rect 8392 26318 8444 26324
rect 8404 26042 8432 26318
rect 8392 26036 8444 26042
rect 8392 25978 8444 25984
rect 8404 25430 8432 25978
rect 8392 25424 8444 25430
rect 8392 25366 8444 25372
rect 8208 25356 8260 25362
rect 8208 25298 8260 25304
rect 8220 24274 8248 25298
rect 8208 24268 8260 24274
rect 8208 24210 8260 24216
rect 8220 23730 8248 24210
rect 8208 23724 8260 23730
rect 8208 23666 8260 23672
rect 8392 22432 8444 22438
rect 8392 22374 8444 22380
rect 8036 22066 8248 22094
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 6736 18896 6788 18902
rect 6736 18838 6788 18844
rect 6748 18086 6776 18838
rect 6932 18766 6960 19314
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 7012 18760 7064 18766
rect 7012 18702 7064 18708
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6932 18086 6960 18566
rect 7024 18358 7052 18702
rect 7012 18352 7064 18358
rect 7012 18294 7064 18300
rect 6736 18080 6788 18086
rect 6736 18022 6788 18028
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6552 17264 6604 17270
rect 6552 17206 6604 17212
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6564 15434 6592 15846
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6552 15428 6604 15434
rect 6552 15370 6604 15376
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6380 12434 6408 13126
rect 6564 12918 6592 15370
rect 6656 14414 6684 15438
rect 6748 15094 6776 18022
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6736 15088 6788 15094
rect 6736 15030 6788 15036
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6656 13394 6684 14350
rect 6644 13388 6696 13394
rect 6644 13330 6696 13336
rect 6552 12912 6604 12918
rect 6552 12854 6604 12860
rect 6012 12406 6132 12434
rect 6380 12406 6592 12434
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 4896 11756 4948 11762
rect 5000 11750 5212 11778
rect 4896 11698 4948 11704
rect 5080 11688 5132 11694
rect 4816 11614 5028 11642
rect 5080 11630 5132 11636
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4724 11150 4752 11494
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3436 9382 3464 9862
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3436 9042 3464 9318
rect 3424 9036 3476 9042
rect 3424 8978 3476 8984
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 2596 8356 2648 8362
rect 2596 8298 2648 8304
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2516 6798 2544 7686
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2320 6248 2372 6254
rect 2320 6190 2372 6196
rect 2332 5914 2360 6190
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2332 5234 2360 5850
rect 2504 5568 2556 5574
rect 2504 5510 2556 5516
rect 2516 5234 2544 5510
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2332 3516 2360 5170
rect 2504 4616 2556 4622
rect 2608 4604 2636 8298
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 2556 4576 2636 4604
rect 2504 4558 2556 4564
rect 2412 3528 2464 3534
rect 2332 3488 2412 3516
rect 2412 3470 2464 3476
rect 2134 3088 2190 3097
rect 2424 3058 2452 3470
rect 2134 3023 2190 3032
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2516 2961 2544 4558
rect 2700 4146 2728 7754
rect 3148 7268 3200 7274
rect 3148 7210 3200 7216
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2976 6798 3004 7142
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2976 6390 3004 6598
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 3068 4282 3096 4558
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 3160 4146 3188 7210
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 2594 4040 2650 4049
rect 2594 3975 2650 3984
rect 2608 3466 2636 3975
rect 2596 3460 2648 3466
rect 2596 3402 2648 3408
rect 2594 3088 2650 3097
rect 2594 3023 2650 3032
rect 2502 2952 2558 2961
rect 2502 2887 2558 2896
rect 2044 2576 2096 2582
rect 2044 2518 2096 2524
rect 2608 2446 2636 3023
rect 2700 2854 2728 4082
rect 2688 2848 2740 2854
rect 2688 2790 2740 2796
rect 3252 2446 3280 8774
rect 3424 8016 3476 8022
rect 3424 7958 3476 7964
rect 3514 7984 3570 7993
rect 3436 6186 3464 7958
rect 3514 7919 3570 7928
rect 3528 7546 3556 7919
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3528 6458 3556 7482
rect 3620 7154 3648 9998
rect 3712 7342 3740 10066
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3896 9625 3924 9862
rect 3882 9616 3938 9625
rect 3882 9551 3938 9560
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4620 8356 4672 8362
rect 4620 8298 4672 8304
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3896 7886 3924 8230
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3804 7410 3832 7686
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3620 7126 3740 7154
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3436 3194 3464 6122
rect 3620 4214 3648 6938
rect 3712 4486 3740 7126
rect 3804 5370 3832 7346
rect 3896 7342 3924 7822
rect 3976 7744 4028 7750
rect 3974 7712 3976 7721
rect 4028 7712 4030 7721
rect 3974 7647 4030 7656
rect 3988 7478 4016 7647
rect 3976 7472 4028 7478
rect 3976 7414 4028 7420
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3700 4480 3752 4486
rect 3700 4422 3752 4428
rect 3712 4282 3740 4422
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3608 4208 3660 4214
rect 3608 4150 3660 4156
rect 3700 4004 3752 4010
rect 3700 3946 3752 3952
rect 3712 3738 3740 3946
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 3804 3194 3832 5102
rect 3988 4758 4016 6870
rect 3976 4752 4028 4758
rect 3976 4694 4028 4700
rect 3976 4548 4028 4554
rect 3976 4490 4028 4496
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3896 3194 3924 4082
rect 3988 4010 4016 4490
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 4080 3398 4108 7822
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4172 4554 4200 4626
rect 4632 4622 4660 8298
rect 4724 8022 4752 10950
rect 4816 8838 4844 11494
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4712 8016 4764 8022
rect 4712 7958 4764 7964
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4160 4548 4212 4554
rect 4160 4490 4212 4496
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 1596 1494 1624 2382
rect 4080 1970 4108 3334
rect 4632 3126 4660 4422
rect 4724 3466 4752 7686
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4816 2446 4844 8774
rect 4908 5234 4936 11086
rect 5000 11014 5028 11614
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 5000 9994 5028 10610
rect 5092 10266 5120 11630
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 5184 10130 5212 11750
rect 5276 11218 5304 12038
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5368 10810 5396 12242
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5264 10736 5316 10742
rect 5460 10690 5488 11494
rect 5264 10678 5316 10684
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 5000 8634 5028 9930
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 5000 7954 5028 8570
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 5092 7410 5120 8910
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5184 7546 5212 7686
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 5276 6934 5304 10678
rect 5368 10662 5488 10690
rect 5368 7002 5396 10662
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5460 7886 5488 10202
rect 5552 9586 5580 12406
rect 5816 12164 5868 12170
rect 5816 12106 5868 12112
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5552 8906 5580 9522
rect 5644 9518 5672 11018
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5552 7478 5580 8230
rect 5644 8022 5672 8434
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5736 7954 5764 8978
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5264 6928 5316 6934
rect 5264 6870 5316 6876
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 5000 5846 5028 6598
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 4988 5840 5040 5846
rect 4988 5782 5040 5788
rect 5092 5370 5120 6054
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 4908 4214 4936 4966
rect 4896 4208 4948 4214
rect 4896 4150 4948 4156
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 4908 3913 4936 4014
rect 4894 3904 4950 3913
rect 4894 3839 4950 3848
rect 4894 3768 4950 3777
rect 5000 3738 5028 4966
rect 5092 4690 5120 5306
rect 5172 5296 5224 5302
rect 5172 5238 5224 5244
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 5078 4584 5134 4593
rect 5078 4519 5134 4528
rect 4894 3703 4896 3712
rect 4948 3703 4950 3712
rect 4988 3732 5040 3738
rect 4896 3674 4948 3680
rect 4988 3674 5040 3680
rect 4894 3224 4950 3233
rect 4894 3159 4950 3168
rect 4908 2854 4936 3159
rect 5092 3058 5120 4519
rect 5184 3466 5212 5238
rect 5276 4729 5304 6734
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5262 4720 5318 4729
rect 5262 4655 5318 4664
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5276 3913 5304 4558
rect 5262 3904 5318 3913
rect 5262 3839 5318 3848
rect 5368 3534 5396 5170
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5172 3460 5224 3466
rect 5172 3402 5224 3408
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 4896 2848 4948 2854
rect 4896 2790 4948 2796
rect 5170 2816 5226 2825
rect 5170 2751 5226 2760
rect 5184 2650 5212 2751
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5276 2514 5304 2926
rect 5368 2650 5396 3130
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 5460 2446 5488 6258
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5538 5536 5594 5545
rect 5538 5471 5594 5480
rect 5552 4622 5580 5471
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5538 4312 5594 4321
rect 5538 4247 5540 4256
rect 5592 4247 5594 4256
rect 5540 4218 5592 4224
rect 5538 4040 5594 4049
rect 5538 3975 5594 3984
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5460 2038 5488 2382
rect 5448 2032 5500 2038
rect 5448 1974 5500 1980
rect 4068 1964 4120 1970
rect 4068 1906 4120 1912
rect 1584 1488 1636 1494
rect 1584 1430 1636 1436
rect 5552 800 5580 3975
rect 5644 2854 5672 6054
rect 5736 5556 5764 7142
rect 5828 6730 5856 12106
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 5920 8430 5948 9454
rect 6104 8673 6132 12406
rect 6564 11234 6592 12406
rect 6656 11762 6684 13330
rect 6840 12850 6868 15302
rect 7024 15162 7052 15438
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 7116 15042 7144 22066
rect 7748 20460 7800 20466
rect 7748 20402 7800 20408
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7668 19378 7696 19654
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7288 19236 7340 19242
rect 7288 19178 7340 19184
rect 7300 18766 7328 19178
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 7288 18760 7340 18766
rect 7288 18702 7340 18708
rect 7196 18624 7248 18630
rect 7196 18566 7248 18572
rect 7208 18426 7236 18566
rect 7196 18420 7248 18426
rect 7196 18362 7248 18368
rect 7300 15570 7328 18702
rect 7392 18290 7420 18770
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7668 18358 7696 18566
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7760 18086 7788 20402
rect 7840 19780 7892 19786
rect 7840 19722 7892 19728
rect 7852 19514 7880 19722
rect 7840 19508 7892 19514
rect 7840 19450 7892 19456
rect 8220 19242 8248 22066
rect 8404 22030 8432 22374
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8208 19236 8260 19242
rect 8208 19178 8260 19184
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8312 18426 8340 19110
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7564 16516 7616 16522
rect 7564 16458 7616 16464
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7024 15014 7144 15042
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6932 12850 6960 13126
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6932 11354 6960 11630
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6644 11280 6696 11286
rect 6564 11228 6644 11234
rect 6564 11222 6696 11228
rect 6734 11248 6790 11257
rect 6564 11206 6684 11222
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6090 8664 6146 8673
rect 6090 8599 6146 8608
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 6000 7812 6052 7818
rect 6000 7754 6052 7760
rect 6012 7002 6040 7754
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5828 5710 5856 6666
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 6012 5794 6040 6258
rect 5920 5766 6040 5794
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5736 5528 5856 5556
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5644 800 5672 2586
rect 5736 800 5764 4966
rect 5828 4185 5856 5528
rect 5814 4176 5870 4185
rect 5814 4111 5870 4120
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5828 2922 5856 4014
rect 5816 2916 5868 2922
rect 5816 2858 5868 2864
rect 5920 2774 5948 5766
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 6012 4826 6040 5170
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 5998 3904 6054 3913
rect 5998 3839 6054 3848
rect 5828 2746 5948 2774
rect 5828 800 5856 2746
rect 6012 1442 6040 3839
rect 6104 3602 6132 6802
rect 6196 6798 6224 7142
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6288 6066 6316 9318
rect 6380 8809 6408 10950
rect 6366 8800 6422 8809
rect 6366 8735 6422 8744
rect 6656 8498 6684 11206
rect 6734 11183 6736 11192
rect 6788 11183 6790 11192
rect 6736 11154 6788 11160
rect 6932 8906 6960 11290
rect 7024 11234 7052 15014
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7116 12442 7144 13806
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7208 11558 7236 12786
rect 7300 12782 7328 15506
rect 7392 15502 7420 16390
rect 7576 15706 7604 16458
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7392 15201 7420 15438
rect 7378 15192 7434 15201
rect 7378 15127 7434 15136
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7300 11257 7328 12718
rect 7286 11248 7342 11257
rect 7024 11206 7144 11234
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 6920 8900 6972 8906
rect 6920 8842 6972 8848
rect 7024 8566 7052 10202
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6196 6038 6316 6066
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6092 3460 6144 3466
rect 6092 3402 6144 3408
rect 5920 1414 6040 1442
rect 5920 800 5948 1414
rect 6104 1170 6132 3402
rect 6196 2446 6224 6038
rect 6380 5302 6408 8366
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6748 6390 6776 7822
rect 7116 7342 7144 11206
rect 7196 11212 7248 11218
rect 7286 11183 7288 11192
rect 7196 11154 7248 11160
rect 7340 11183 7342 11192
rect 7288 11154 7340 11160
rect 7208 11064 7236 11154
rect 7300 11123 7328 11154
rect 7392 11064 7420 14554
rect 7656 14408 7708 14414
rect 7656 14350 7708 14356
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7484 14006 7512 14214
rect 7668 14074 7696 14350
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7472 14000 7524 14006
rect 7472 13942 7524 13948
rect 7564 14000 7616 14006
rect 7564 13942 7616 13948
rect 7472 13184 7524 13190
rect 7576 13172 7604 13942
rect 7524 13144 7604 13172
rect 7472 13126 7524 13132
rect 7484 12918 7512 13126
rect 7472 12912 7524 12918
rect 7472 12854 7524 12860
rect 7484 11150 7512 12854
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7208 11036 7420 11064
rect 7484 10810 7512 11086
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7668 10266 7696 10610
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7472 8900 7524 8906
rect 7472 8842 7524 8848
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 6368 5296 6420 5302
rect 6368 5238 6420 5244
rect 6276 5092 6328 5098
rect 6276 5034 6328 5040
rect 6288 4622 6316 5034
rect 6472 5030 6500 6326
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6288 4282 6316 4558
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 6472 4026 6500 4966
rect 6564 4282 6592 5102
rect 6656 4622 6684 6054
rect 6748 5914 6776 6326
rect 6828 6248 6880 6254
rect 6880 6208 6960 6236
rect 6828 6190 6880 6196
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6932 5710 6960 6208
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 7024 5710 7052 6122
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6828 5636 6880 5642
rect 6828 5578 6880 5584
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6748 5302 6776 5510
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 6748 4826 6776 5238
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6736 4548 6788 4554
rect 6736 4490 6788 4496
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6564 4078 6592 4218
rect 6380 3998 6500 4026
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6380 3738 6408 3998
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 6012 1142 6132 1170
rect 6012 800 6040 1142
rect 6196 1034 6224 2382
rect 6104 1006 6224 1034
rect 6104 800 6132 1006
rect 6184 944 6236 950
rect 6184 886 6236 892
rect 6196 800 6224 886
rect 6288 800 6316 3674
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6380 3210 6408 3538
rect 6472 3346 6500 3878
rect 6472 3318 6684 3346
rect 6380 3182 6500 3210
rect 6366 2952 6422 2961
rect 6366 2887 6422 2896
rect 6380 800 6408 2887
rect 6472 800 6500 3182
rect 6550 2680 6606 2689
rect 6550 2615 6552 2624
rect 6604 2615 6606 2624
rect 6552 2586 6604 2592
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 6564 800 6592 2450
rect 6656 800 6684 3318
rect 6748 950 6776 4490
rect 6840 3058 6868 5578
rect 6932 4010 6960 5646
rect 7024 5234 7052 5646
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7012 4752 7064 4758
rect 7012 4694 7064 4700
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 6918 3088 6974 3097
rect 6828 3052 6880 3058
rect 6918 3023 6974 3032
rect 6828 2994 6880 3000
rect 6736 944 6788 950
rect 6736 886 6788 892
rect 6840 800 6868 2994
rect 6932 800 6960 3023
rect 7024 800 7052 4694
rect 7116 4622 7144 6598
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 7116 4282 7144 4422
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7102 4176 7158 4185
rect 7102 4111 7158 4120
rect 7116 3942 7144 4111
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7208 2446 7236 8774
rect 7484 7886 7512 8842
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7300 4486 7328 6190
rect 7392 5710 7420 6802
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7300 3058 7328 4422
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7392 2774 7420 5646
rect 7484 4282 7512 7822
rect 7576 6798 7604 8298
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7484 3738 7512 4014
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7484 2854 7512 3674
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7300 2746 7420 2774
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7208 800 7236 2382
rect 7300 800 7328 2746
rect 7380 2576 7432 2582
rect 7380 2518 7432 2524
rect 7392 800 7420 2518
rect 7576 800 7604 6734
rect 7760 5914 7788 18022
rect 8220 14414 8248 18226
rect 8496 15706 8524 27542
rect 9036 25696 9088 25702
rect 9036 25638 9088 25644
rect 9048 22094 9076 25638
rect 8956 22066 9076 22094
rect 8956 21962 8984 22066
rect 8944 21956 8996 21962
rect 8944 21898 8996 21904
rect 8956 21350 8984 21898
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 8668 15904 8720 15910
rect 8668 15846 8720 15852
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8312 15162 8340 15438
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8220 13326 8248 14350
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8220 12850 8248 13262
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 7944 12238 7972 12378
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 7944 11830 7972 12174
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 7944 10674 7972 11766
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 7944 7546 7972 7958
rect 8036 7818 8064 8230
rect 8024 7812 8076 7818
rect 8024 7754 8076 7760
rect 8036 7546 8064 7754
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7668 4826 7696 5170
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7760 4758 7788 4966
rect 7748 4752 7800 4758
rect 7748 4694 7800 4700
rect 7852 4554 7880 5170
rect 8036 5030 8064 6598
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 7932 4616 7984 4622
rect 8036 4604 8064 4966
rect 7984 4576 8064 4604
rect 7932 4558 7984 4564
rect 7840 4548 7892 4554
rect 7840 4490 7892 4496
rect 7654 4312 7710 4321
rect 7654 4247 7656 4256
rect 7708 4247 7710 4256
rect 7656 4218 7708 4224
rect 7852 4078 7880 4490
rect 7944 4146 7972 4558
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7944 3058 7972 4082
rect 8022 3088 8078 3097
rect 7932 3052 7984 3058
rect 8022 3023 8078 3032
rect 7932 2994 7984 3000
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7668 800 7696 2926
rect 7760 2825 7788 2926
rect 7840 2916 7892 2922
rect 7840 2858 7892 2864
rect 7746 2816 7802 2825
rect 7746 2751 7802 2760
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7760 800 7788 2246
rect 7852 800 7880 2858
rect 7932 2848 7984 2854
rect 7932 2790 7984 2796
rect 7944 2514 7972 2790
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 7932 1896 7984 1902
rect 7932 1838 7984 1844
rect 7944 800 7972 1838
rect 8036 800 8064 3023
rect 8128 2378 8156 8774
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8220 7342 8248 8570
rect 8576 8424 8628 8430
rect 8574 8392 8576 8401
rect 8628 8392 8630 8401
rect 8574 8327 8630 8336
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8220 3670 8248 7142
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8206 3224 8262 3233
rect 8206 3159 8208 3168
rect 8260 3159 8262 3168
rect 8208 3130 8260 3136
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8116 2372 8168 2378
rect 8116 2314 8168 2320
rect 8128 1902 8156 2314
rect 8116 1896 8168 1902
rect 8116 1838 8168 1844
rect 8116 1488 8168 1494
rect 8116 1430 8168 1436
rect 8128 800 8156 1430
rect 8220 800 8248 2994
rect 8312 800 8340 4422
rect 8404 800 8432 6734
rect 8576 6724 8628 6730
rect 8576 6666 8628 6672
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8496 4078 8524 6258
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8496 2990 8524 4014
rect 8588 3126 8616 6666
rect 8680 4826 8708 15846
rect 8760 14816 8812 14822
rect 8852 14816 8904 14822
rect 8760 14758 8812 14764
rect 8850 14784 8852 14793
rect 8904 14784 8906 14793
rect 8772 13802 8800 14758
rect 8850 14719 8906 14728
rect 8760 13796 8812 13802
rect 8760 13738 8812 13744
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8772 11762 8800 12582
rect 8956 12434 8984 21286
rect 9140 20330 9168 34682
rect 9324 32910 9352 35566
rect 9508 34678 9536 35974
rect 9784 35630 9812 36722
rect 9772 35624 9824 35630
rect 9772 35566 9824 35572
rect 9496 34672 9548 34678
rect 9496 34614 9548 34620
rect 9588 34604 9640 34610
rect 9588 34546 9640 34552
rect 9600 34241 9628 34546
rect 9586 34232 9642 34241
rect 9586 34167 9642 34176
rect 9312 32904 9364 32910
rect 9312 32846 9364 32852
rect 9784 32842 9812 35566
rect 10060 35154 10088 37246
rect 10244 37194 10272 38150
rect 10414 38040 10470 38049
rect 10520 38026 10548 39782
rect 10612 39302 10640 41074
rect 10692 40044 10744 40050
rect 10692 39986 10744 39992
rect 10600 39296 10652 39302
rect 10600 39238 10652 39244
rect 10612 38350 10640 39238
rect 10704 38962 10732 39986
rect 11072 39438 11100 41142
rect 12452 40390 12480 41482
rect 13004 41274 13032 41482
rect 13084 41472 13136 41478
rect 13084 41414 13136 41420
rect 13544 41472 13596 41478
rect 13544 41414 13596 41420
rect 12992 41268 13044 41274
rect 12992 41210 13044 41216
rect 12624 40928 12676 40934
rect 12624 40870 12676 40876
rect 12636 40526 12664 40870
rect 12624 40520 12676 40526
rect 12624 40462 12676 40468
rect 12808 40520 12860 40526
rect 12808 40462 12860 40468
rect 12440 40384 12492 40390
rect 12440 40326 12492 40332
rect 12624 40384 12676 40390
rect 12624 40326 12676 40332
rect 11244 40180 11296 40186
rect 11244 40122 11296 40128
rect 11256 39438 11284 40122
rect 11704 40044 11756 40050
rect 11704 39986 11756 39992
rect 11716 39642 11744 39986
rect 11704 39636 11756 39642
rect 11704 39578 11756 39584
rect 11060 39432 11112 39438
rect 11060 39374 11112 39380
rect 11244 39432 11296 39438
rect 11244 39374 11296 39380
rect 10692 38956 10744 38962
rect 10692 38898 10744 38904
rect 10600 38344 10652 38350
rect 10600 38286 10652 38292
rect 10470 37998 10548 38026
rect 10414 37975 10470 37984
rect 10428 37942 10456 37975
rect 10416 37936 10468 37942
rect 10416 37878 10468 37884
rect 10232 37188 10284 37194
rect 10232 37130 10284 37136
rect 10244 36174 10272 37130
rect 10232 36168 10284 36174
rect 10232 36110 10284 36116
rect 10140 36032 10192 36038
rect 10140 35974 10192 35980
rect 10152 35630 10180 35974
rect 10244 35698 10272 36110
rect 10416 36100 10468 36106
rect 10416 36042 10468 36048
rect 10232 35692 10284 35698
rect 10232 35634 10284 35640
rect 10140 35624 10192 35630
rect 10140 35566 10192 35572
rect 10048 35148 10100 35154
rect 10048 35090 10100 35096
rect 9956 35080 10008 35086
rect 9956 35022 10008 35028
rect 9968 34610 9996 35022
rect 9956 34604 10008 34610
rect 9956 34546 10008 34552
rect 9864 32972 9916 32978
rect 9864 32914 9916 32920
rect 9772 32836 9824 32842
rect 9772 32778 9824 32784
rect 9784 32722 9812 32778
rect 9692 32694 9812 32722
rect 9404 32496 9456 32502
rect 9404 32438 9456 32444
rect 9220 30048 9272 30054
rect 9220 29990 9272 29996
rect 9232 29646 9260 29990
rect 9220 29640 9272 29646
rect 9220 29582 9272 29588
rect 9416 29238 9444 32438
rect 9404 29232 9456 29238
rect 9404 29174 9456 29180
rect 9312 28552 9364 28558
rect 9312 28494 9364 28500
rect 9324 27538 9352 28494
rect 9416 28218 9444 29174
rect 9496 28960 9548 28966
rect 9496 28902 9548 28908
rect 9508 28558 9536 28902
rect 9496 28552 9548 28558
rect 9496 28494 9548 28500
rect 9692 28422 9720 32694
rect 9876 30258 9904 32914
rect 9968 32502 9996 34546
rect 10060 34542 10088 35090
rect 10048 34536 10100 34542
rect 10048 34478 10100 34484
rect 10060 34066 10088 34478
rect 10048 34060 10100 34066
rect 10048 34002 10100 34008
rect 10152 33998 10180 35566
rect 10244 35154 10272 35634
rect 10232 35148 10284 35154
rect 10232 35090 10284 35096
rect 10428 34746 10456 36042
rect 10704 35630 10732 38898
rect 11072 37942 11100 39374
rect 11060 37936 11112 37942
rect 11060 37878 11112 37884
rect 11072 36378 11100 37878
rect 11256 37874 11284 39374
rect 12452 37942 12480 40326
rect 12636 40118 12664 40326
rect 12820 40186 12848 40462
rect 13004 40440 13032 41210
rect 13096 41138 13124 41414
rect 13084 41132 13136 41138
rect 13084 41074 13136 41080
rect 13556 41002 13584 41414
rect 13544 40996 13596 41002
rect 13544 40938 13596 40944
rect 13084 40452 13136 40458
rect 13004 40412 13084 40440
rect 13084 40394 13136 40400
rect 12808 40180 12860 40186
rect 12808 40122 12860 40128
rect 12624 40112 12676 40118
rect 12624 40054 12676 40060
rect 12532 38004 12584 38010
rect 12532 37946 12584 37952
rect 12440 37936 12492 37942
rect 12440 37878 12492 37884
rect 11244 37868 11296 37874
rect 11244 37810 11296 37816
rect 11888 37868 11940 37874
rect 11888 37810 11940 37816
rect 11900 37262 11928 37810
rect 11888 37256 11940 37262
rect 11888 37198 11940 37204
rect 12544 36922 12572 37946
rect 12532 36916 12584 36922
rect 12532 36858 12584 36864
rect 12544 36378 12572 36858
rect 11060 36372 11112 36378
rect 11060 36314 11112 36320
rect 12532 36372 12584 36378
rect 12532 36314 12584 36320
rect 11072 35766 11100 36314
rect 11704 36032 11756 36038
rect 11704 35974 11756 35980
rect 11060 35760 11112 35766
rect 11060 35702 11112 35708
rect 11520 35760 11572 35766
rect 11520 35702 11572 35708
rect 10692 35624 10744 35630
rect 10692 35566 10744 35572
rect 10600 35488 10652 35494
rect 10600 35430 10652 35436
rect 10416 34740 10468 34746
rect 10416 34682 10468 34688
rect 10612 33998 10640 35430
rect 11060 35012 11112 35018
rect 11060 34954 11112 34960
rect 10968 34604 11020 34610
rect 10968 34546 11020 34552
rect 10140 33992 10192 33998
rect 10140 33934 10192 33940
rect 10600 33992 10652 33998
rect 10600 33934 10652 33940
rect 10980 33318 11008 34546
rect 11072 34202 11100 34954
rect 11532 34610 11560 35702
rect 11716 34610 11744 35974
rect 11980 35692 12032 35698
rect 11980 35634 12032 35640
rect 11992 35290 12020 35634
rect 11980 35284 12032 35290
rect 11980 35226 12032 35232
rect 11992 35086 12020 35226
rect 11980 35080 12032 35086
rect 11980 35022 12032 35028
rect 12820 34678 12848 40122
rect 13096 39098 13124 40394
rect 13084 39092 13136 39098
rect 13084 39034 13136 39040
rect 12900 38956 12952 38962
rect 12900 38898 12952 38904
rect 12912 37806 12940 38898
rect 12900 37800 12952 37806
rect 12900 37742 12952 37748
rect 12808 34672 12860 34678
rect 12808 34614 12860 34620
rect 11520 34604 11572 34610
rect 11520 34546 11572 34552
rect 11704 34604 11756 34610
rect 11704 34546 11756 34552
rect 11520 34468 11572 34474
rect 11520 34410 11572 34416
rect 11060 34196 11112 34202
rect 11060 34138 11112 34144
rect 11532 33998 11560 34410
rect 11796 34400 11848 34406
rect 11796 34342 11848 34348
rect 11520 33992 11572 33998
rect 11520 33934 11572 33940
rect 11704 33516 11756 33522
rect 11704 33458 11756 33464
rect 10968 33312 11020 33318
rect 10968 33254 11020 33260
rect 10140 32836 10192 32842
rect 10140 32778 10192 32784
rect 10692 32836 10744 32842
rect 10692 32778 10744 32784
rect 9956 32496 10008 32502
rect 9956 32438 10008 32444
rect 10152 31754 10180 32778
rect 10416 32360 10468 32366
rect 10416 32302 10468 32308
rect 10428 32230 10456 32302
rect 10704 32230 10732 32778
rect 10980 32774 11008 33254
rect 11060 32904 11112 32910
rect 11060 32846 11112 32852
rect 10784 32768 10836 32774
rect 10784 32710 10836 32716
rect 10968 32768 11020 32774
rect 10968 32710 11020 32716
rect 10796 32434 10824 32710
rect 10980 32434 11008 32710
rect 10784 32428 10836 32434
rect 10784 32370 10836 32376
rect 10968 32428 11020 32434
rect 10968 32370 11020 32376
rect 10980 32314 11008 32370
rect 10888 32286 11008 32314
rect 10324 32224 10376 32230
rect 10324 32166 10376 32172
rect 10416 32224 10468 32230
rect 10416 32166 10468 32172
rect 10692 32224 10744 32230
rect 10692 32166 10744 32172
rect 10336 31822 10364 32166
rect 10324 31816 10376 31822
rect 10324 31758 10376 31764
rect 10152 31726 10272 31754
rect 10140 31340 10192 31346
rect 10140 31282 10192 31288
rect 10152 31142 10180 31282
rect 10140 31136 10192 31142
rect 10140 31078 10192 31084
rect 10048 30592 10100 30598
rect 10048 30534 10100 30540
rect 9864 30252 9916 30258
rect 9864 30194 9916 30200
rect 10060 30190 10088 30534
rect 10048 30184 10100 30190
rect 10048 30126 10100 30132
rect 10060 29578 10088 30126
rect 10048 29572 10100 29578
rect 10048 29514 10100 29520
rect 9956 29504 10008 29510
rect 9956 29446 10008 29452
rect 9968 29034 9996 29446
rect 9956 29028 10008 29034
rect 9956 28970 10008 28976
rect 9772 28484 9824 28490
rect 9772 28426 9824 28432
rect 9680 28416 9732 28422
rect 9680 28358 9732 28364
rect 9404 28212 9456 28218
rect 9404 28154 9456 28160
rect 9680 28144 9732 28150
rect 9680 28086 9732 28092
rect 9496 28076 9548 28082
rect 9496 28018 9548 28024
rect 9508 27878 9536 28018
rect 9496 27872 9548 27878
rect 9496 27814 9548 27820
rect 9312 27532 9364 27538
rect 9312 27474 9364 27480
rect 9508 27470 9536 27814
rect 9220 27464 9272 27470
rect 9220 27406 9272 27412
rect 9496 27464 9548 27470
rect 9496 27406 9548 27412
rect 9232 26994 9260 27406
rect 9220 26988 9272 26994
rect 9220 26930 9272 26936
rect 9312 26852 9364 26858
rect 9312 26794 9364 26800
rect 9220 26784 9272 26790
rect 9220 26726 9272 26732
rect 9232 23118 9260 26726
rect 9324 26314 9352 26794
rect 9508 26790 9536 27406
rect 9496 26784 9548 26790
rect 9496 26726 9548 26732
rect 9312 26308 9364 26314
rect 9312 26250 9364 26256
rect 9324 23866 9352 26250
rect 9692 25906 9720 28086
rect 9784 28014 9812 28426
rect 9968 28098 9996 28970
rect 10048 28416 10100 28422
rect 10048 28358 10100 28364
rect 9876 28070 9996 28098
rect 9772 28008 9824 28014
rect 9772 27950 9824 27956
rect 9772 25968 9824 25974
rect 9772 25910 9824 25916
rect 9680 25900 9732 25906
rect 9680 25842 9732 25848
rect 9496 25832 9548 25838
rect 9496 25774 9548 25780
rect 9312 23860 9364 23866
rect 9312 23802 9364 23808
rect 9324 23186 9352 23802
rect 9312 23180 9364 23186
rect 9312 23122 9364 23128
rect 9220 23112 9272 23118
rect 9220 23054 9272 23060
rect 9128 20324 9180 20330
rect 9128 20266 9180 20272
rect 9220 20256 9272 20262
rect 9220 20198 9272 20204
rect 9232 19446 9260 20198
rect 9220 19440 9272 19446
rect 9220 19382 9272 19388
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 9232 18086 9260 18226
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9232 17814 9260 18022
rect 9220 17808 9272 17814
rect 9220 17750 9272 17756
rect 9404 16584 9456 16590
rect 9404 16526 9456 16532
rect 9416 14550 9444 16526
rect 9508 15094 9536 25774
rect 9784 25294 9812 25910
rect 9772 25288 9824 25294
rect 9772 25230 9824 25236
rect 9876 25140 9904 28070
rect 9956 26920 10008 26926
rect 9956 26862 10008 26868
rect 9968 25158 9996 26862
rect 10060 25974 10088 28358
rect 10048 25968 10100 25974
rect 10048 25910 10100 25916
rect 10048 25220 10100 25226
rect 10048 25162 10100 25168
rect 9692 25112 9904 25140
rect 9956 25152 10008 25158
rect 9692 22234 9720 25112
rect 9956 25094 10008 25100
rect 9772 24608 9824 24614
rect 9772 24550 9824 24556
rect 9784 24206 9812 24550
rect 9772 24200 9824 24206
rect 9772 24142 9824 24148
rect 9862 24168 9918 24177
rect 9862 24103 9864 24112
rect 9916 24103 9918 24112
rect 9864 24074 9916 24080
rect 9772 23860 9824 23866
rect 9772 23802 9824 23808
rect 9680 22228 9732 22234
rect 9680 22170 9732 22176
rect 9784 21622 9812 23802
rect 9864 22772 9916 22778
rect 9864 22714 9916 22720
rect 9772 21616 9824 21622
rect 9772 21558 9824 21564
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 9600 18766 9628 19790
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9600 18222 9628 18702
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 9600 17202 9628 18158
rect 9876 17882 9904 22714
rect 9968 22094 9996 25094
rect 10060 23866 10088 25162
rect 10152 24410 10180 31078
rect 10244 29850 10272 31726
rect 10232 29844 10284 29850
rect 10232 29786 10284 29792
rect 10784 29640 10836 29646
rect 10784 29582 10836 29588
rect 10600 29232 10652 29238
rect 10600 29174 10652 29180
rect 10612 28422 10640 29174
rect 10600 28416 10652 28422
rect 10600 28358 10652 28364
rect 10612 28150 10640 28358
rect 10600 28144 10652 28150
rect 10600 28086 10652 28092
rect 10796 27996 10824 29582
rect 10888 29170 10916 32286
rect 10968 32224 11020 32230
rect 10968 32166 11020 32172
rect 10980 30326 11008 32166
rect 11072 32026 11100 32846
rect 11060 32020 11112 32026
rect 11060 31962 11112 31968
rect 11072 30734 11100 31962
rect 11336 31952 11388 31958
rect 11336 31894 11388 31900
rect 11348 31657 11376 31894
rect 11334 31648 11390 31657
rect 11334 31583 11390 31592
rect 11060 30728 11112 30734
rect 11060 30670 11112 30676
rect 10968 30320 11020 30326
rect 10968 30262 11020 30268
rect 11060 30252 11112 30258
rect 11060 30194 11112 30200
rect 10968 29844 11020 29850
rect 10968 29786 11020 29792
rect 10980 29238 11008 29786
rect 11072 29510 11100 30194
rect 11060 29504 11112 29510
rect 11060 29446 11112 29452
rect 11072 29238 11100 29446
rect 10968 29232 11020 29238
rect 10968 29174 11020 29180
rect 11060 29232 11112 29238
rect 11060 29174 11112 29180
rect 10876 29164 10928 29170
rect 10876 29106 10928 29112
rect 10968 29028 11020 29034
rect 10968 28970 11020 28976
rect 10876 28008 10928 28014
rect 10796 27968 10876 27996
rect 10876 27950 10928 27956
rect 10888 27470 10916 27950
rect 10876 27464 10928 27470
rect 10876 27406 10928 27412
rect 10508 27124 10560 27130
rect 10508 27066 10560 27072
rect 10416 24948 10468 24954
rect 10416 24890 10468 24896
rect 10232 24812 10284 24818
rect 10232 24754 10284 24760
rect 10140 24404 10192 24410
rect 10140 24346 10192 24352
rect 10048 23860 10100 23866
rect 10048 23802 10100 23808
rect 10244 23322 10272 24754
rect 10324 24064 10376 24070
rect 10324 24006 10376 24012
rect 10232 23316 10284 23322
rect 10232 23258 10284 23264
rect 10336 23118 10364 24006
rect 10324 23112 10376 23118
rect 10324 23054 10376 23060
rect 9968 22066 10180 22094
rect 10048 21956 10100 21962
rect 10048 21898 10100 21904
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9968 21554 9996 21830
rect 10060 21690 10088 21898
rect 10048 21684 10100 21690
rect 10048 21626 10100 21632
rect 10060 21554 10088 21626
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 10048 21548 10100 21554
rect 10048 21490 10100 21496
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9600 16658 9628 17138
rect 9692 16794 9720 17614
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9496 15088 9548 15094
rect 9496 15030 9548 15036
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9600 14822 9628 14962
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9600 14550 9628 14758
rect 9404 14544 9456 14550
rect 9404 14486 9456 14492
rect 9588 14544 9640 14550
rect 9588 14486 9640 14492
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9404 13456 9456 13462
rect 9404 13398 9456 13404
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 8864 12406 8984 12434
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 8772 8498 8800 8842
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8864 8378 8892 12406
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8956 10742 8984 10950
rect 8944 10736 8996 10742
rect 8944 10678 8996 10684
rect 9048 8514 9076 13126
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9140 10810 9168 11086
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 9416 9178 9444 13398
rect 9508 13190 9536 13670
rect 9600 13530 9628 14282
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9600 12714 9628 13466
rect 9588 12708 9640 12714
rect 9588 12650 9640 12656
rect 9496 12368 9548 12374
rect 9496 12310 9548 12316
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9220 8900 9272 8906
rect 9220 8842 9272 8848
rect 9048 8486 9168 8514
rect 8772 8362 8892 8378
rect 8760 8356 8892 8362
rect 8812 8350 8892 8356
rect 8760 8298 8812 8304
rect 8772 7206 8800 8298
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8760 7200 8812 7206
rect 8760 7142 8812 7148
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8668 4072 8720 4078
rect 8666 4040 8668 4049
rect 8720 4040 8722 4049
rect 8772 4010 8800 6802
rect 8864 5710 8892 8230
rect 8944 7744 8996 7750
rect 8996 7704 9076 7732
rect 8944 7686 8996 7692
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8666 3975 8722 3984
rect 8760 4004 8812 4010
rect 8760 3946 8812 3952
rect 8772 3777 8800 3946
rect 8758 3768 8814 3777
rect 8758 3703 8814 3712
rect 8864 3126 8892 5306
rect 8956 3942 8984 6598
rect 9048 6322 9076 7704
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9036 5840 9088 5846
rect 9036 5782 9088 5788
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 9048 3534 9076 5782
rect 9140 4622 9168 8486
rect 9232 7886 9260 8842
rect 9324 8430 9352 8978
rect 9508 8786 9536 12310
rect 9600 9110 9628 12650
rect 9692 12170 9720 16730
rect 9864 16720 9916 16726
rect 9864 16662 9916 16668
rect 9876 15502 9904 16662
rect 10152 16250 10180 22066
rect 10336 21962 10364 23054
rect 10428 22094 10456 24890
rect 10520 23730 10548 27066
rect 10692 25152 10744 25158
rect 10692 25094 10744 25100
rect 10704 23730 10732 25094
rect 10784 24948 10836 24954
rect 10784 24890 10836 24896
rect 10796 24138 10824 24890
rect 10876 24880 10928 24886
rect 10876 24822 10928 24828
rect 10784 24132 10836 24138
rect 10784 24074 10836 24080
rect 10888 23730 10916 24822
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 10692 23724 10744 23730
rect 10692 23666 10744 23672
rect 10876 23724 10928 23730
rect 10876 23666 10928 23672
rect 10520 22778 10548 23666
rect 10508 22772 10560 22778
rect 10508 22714 10560 22720
rect 10980 22094 11008 28970
rect 11152 27464 11204 27470
rect 11152 27406 11204 27412
rect 11164 26926 11192 27406
rect 11152 26920 11204 26926
rect 11152 26862 11204 26868
rect 11060 24064 11112 24070
rect 11060 24006 11112 24012
rect 11072 23798 11100 24006
rect 11060 23792 11112 23798
rect 11060 23734 11112 23740
rect 10428 22066 10548 22094
rect 10416 22024 10468 22030
rect 10416 21966 10468 21972
rect 10324 21956 10376 21962
rect 10324 21898 10376 21904
rect 10428 21554 10456 21966
rect 10416 21548 10468 21554
rect 10416 21490 10468 21496
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 10336 17202 10364 18022
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10244 16114 10272 16594
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10428 16182 10456 16390
rect 10416 16176 10468 16182
rect 10416 16118 10468 16124
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10244 15706 10272 16050
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9784 14346 9812 14894
rect 10520 14822 10548 22066
rect 10888 22066 11008 22094
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 10796 20942 10824 21286
rect 10888 21146 10916 22066
rect 10968 21888 11020 21894
rect 10968 21830 11020 21836
rect 10876 21140 10928 21146
rect 10876 21082 10928 21088
rect 10784 20936 10836 20942
rect 10784 20878 10836 20884
rect 10888 19258 10916 21082
rect 10796 19242 10916 19258
rect 10784 19236 10916 19242
rect 10836 19230 10916 19236
rect 10784 19178 10836 19184
rect 10692 19168 10744 19174
rect 10690 19136 10692 19145
rect 10744 19136 10746 19145
rect 10690 19071 10746 19080
rect 10888 18902 10916 19230
rect 10876 18896 10928 18902
rect 10876 18838 10928 18844
rect 10600 18692 10652 18698
rect 10600 18634 10652 18640
rect 10612 17678 10640 18634
rect 10888 18290 10916 18838
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 10888 18154 10916 18226
rect 10876 18148 10928 18154
rect 10876 18090 10928 18096
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10060 14618 10088 14758
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 9772 14340 9824 14346
rect 9772 14282 9824 14288
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9692 10130 9720 12106
rect 9784 11121 9812 14010
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9864 13796 9916 13802
rect 9864 13738 9916 13744
rect 9876 13462 9904 13738
rect 10060 13530 10088 13874
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9876 13190 9904 13262
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9770 11112 9826 11121
rect 9770 11047 9826 11056
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9680 9920 9732 9926
rect 9784 9908 9812 10406
rect 9732 9880 9812 9908
rect 9680 9862 9732 9868
rect 9692 9586 9720 9862
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9416 8758 9536 8786
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9416 8294 9444 8758
rect 9600 8537 9628 8774
rect 9692 8634 9720 9114
rect 10152 8634 10180 14282
rect 10612 13530 10640 16934
rect 10980 16590 11008 21830
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 11072 19242 11100 20198
rect 11060 19236 11112 19242
rect 11060 19178 11112 19184
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 11072 18358 11100 18566
rect 11060 18352 11112 18358
rect 11060 18294 11112 18300
rect 11072 16590 11100 18294
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 11164 16250 11192 26862
rect 11348 24954 11376 31583
rect 11716 30258 11744 33458
rect 11808 31754 11836 34342
rect 12808 32564 12860 32570
rect 12808 32506 12860 32512
rect 11808 31726 12112 31754
rect 11704 30252 11756 30258
rect 11704 30194 11756 30200
rect 11612 29300 11664 29306
rect 11612 29242 11664 29248
rect 11624 28082 11652 29242
rect 11716 29102 11744 30194
rect 11888 30184 11940 30190
rect 11888 30126 11940 30132
rect 11900 29850 11928 30126
rect 11888 29844 11940 29850
rect 11888 29786 11940 29792
rect 11900 29714 11928 29786
rect 11888 29708 11940 29714
rect 11888 29650 11940 29656
rect 11704 29096 11756 29102
rect 11704 29038 11756 29044
rect 11612 28076 11664 28082
rect 11612 28018 11664 28024
rect 11624 26586 11652 28018
rect 11612 26580 11664 26586
rect 11612 26522 11664 26528
rect 11716 25430 11744 29038
rect 11796 28076 11848 28082
rect 11796 28018 11848 28024
rect 11808 27674 11836 28018
rect 11796 27668 11848 27674
rect 11796 27610 11848 27616
rect 11704 25424 11756 25430
rect 11704 25366 11756 25372
rect 11336 24948 11388 24954
rect 11336 24890 11388 24896
rect 11704 24812 11756 24818
rect 11704 24754 11756 24760
rect 11428 24744 11480 24750
rect 11428 24686 11480 24692
rect 11336 24336 11388 24342
rect 11336 24278 11388 24284
rect 11244 23724 11296 23730
rect 11244 23666 11296 23672
rect 11256 23254 11284 23666
rect 11348 23254 11376 24278
rect 11440 24206 11468 24686
rect 11716 24206 11744 24754
rect 11980 24608 12032 24614
rect 12084 24596 12112 31726
rect 12348 31136 12400 31142
rect 12348 31078 12400 31084
rect 12360 30938 12388 31078
rect 12348 30932 12400 30938
rect 12348 30874 12400 30880
rect 12256 29640 12308 29646
rect 12256 29582 12308 29588
rect 12164 27464 12216 27470
rect 12164 27406 12216 27412
rect 12176 26450 12204 27406
rect 12164 26444 12216 26450
rect 12164 26386 12216 26392
rect 12164 24608 12216 24614
rect 12084 24568 12164 24596
rect 11980 24550 12032 24556
rect 12164 24550 12216 24556
rect 11428 24200 11480 24206
rect 11428 24142 11480 24148
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 11440 23662 11468 24142
rect 11796 24132 11848 24138
rect 11796 24074 11848 24080
rect 11428 23656 11480 23662
rect 11428 23598 11480 23604
rect 11612 23520 11664 23526
rect 11612 23462 11664 23468
rect 11244 23248 11296 23254
rect 11244 23190 11296 23196
rect 11336 23248 11388 23254
rect 11336 23190 11388 23196
rect 11244 23112 11296 23118
rect 11244 23054 11296 23060
rect 11428 23112 11480 23118
rect 11428 23054 11480 23060
rect 11256 22778 11284 23054
rect 11244 22772 11296 22778
rect 11244 22714 11296 22720
rect 11244 22024 11296 22030
rect 11244 21966 11296 21972
rect 11256 21486 11284 21966
rect 11440 21962 11468 23054
rect 11624 23050 11652 23462
rect 11808 23322 11836 24074
rect 11796 23316 11848 23322
rect 11796 23258 11848 23264
rect 11612 23044 11664 23050
rect 11612 22986 11664 22992
rect 11624 22094 11652 22986
rect 11532 22066 11652 22094
rect 11704 22092 11756 22098
rect 11532 22030 11560 22066
rect 11704 22034 11756 22040
rect 11520 22024 11572 22030
rect 11520 21966 11572 21972
rect 11716 21962 11744 22034
rect 11428 21956 11480 21962
rect 11428 21898 11480 21904
rect 11704 21956 11756 21962
rect 11704 21898 11756 21904
rect 11440 21690 11468 21898
rect 11428 21684 11480 21690
rect 11428 21626 11480 21632
rect 11244 21480 11296 21486
rect 11244 21422 11296 21428
rect 11520 21412 11572 21418
rect 11520 21354 11572 21360
rect 11428 20936 11480 20942
rect 11428 20878 11480 20884
rect 11440 20262 11468 20878
rect 11428 20256 11480 20262
rect 11428 20198 11480 20204
rect 11428 18216 11480 18222
rect 11428 18158 11480 18164
rect 11440 17338 11468 18158
rect 11428 17332 11480 17338
rect 11428 17274 11480 17280
rect 11244 16516 11296 16522
rect 11244 16458 11296 16464
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11256 16182 11284 16458
rect 11244 16176 11296 16182
rect 11244 16118 11296 16124
rect 11532 16114 11560 21354
rect 11992 20602 12020 24550
rect 12176 21690 12204 24550
rect 12268 23254 12296 29582
rect 12360 24682 12388 30874
rect 12820 29306 12848 32506
rect 12912 31890 12940 37742
rect 13176 37256 13228 37262
rect 13176 37198 13228 37204
rect 13084 36100 13136 36106
rect 13084 36042 13136 36048
rect 13096 35578 13124 36042
rect 13188 35766 13216 37198
rect 13556 37097 13584 40938
rect 13542 37088 13598 37097
rect 13542 37023 13598 37032
rect 13360 36100 13412 36106
rect 13360 36042 13412 36048
rect 13372 35834 13400 36042
rect 13360 35828 13412 35834
rect 13360 35770 13412 35776
rect 13176 35760 13228 35766
rect 13176 35702 13228 35708
rect 13452 35692 13504 35698
rect 13452 35634 13504 35640
rect 13096 35550 13216 35578
rect 13188 35018 13216 35550
rect 13464 35086 13492 35634
rect 13452 35080 13504 35086
rect 13452 35022 13504 35028
rect 13176 35012 13228 35018
rect 13176 34954 13228 34960
rect 13188 34626 13216 34954
rect 13188 34610 13308 34626
rect 13464 34610 13492 35022
rect 13188 34604 13320 34610
rect 13188 34598 13268 34604
rect 13268 34546 13320 34552
rect 13452 34604 13504 34610
rect 13452 34546 13504 34552
rect 13176 34536 13228 34542
rect 13176 34478 13228 34484
rect 12992 33312 13044 33318
rect 12992 33254 13044 33260
rect 13004 32842 13032 33254
rect 12992 32836 13044 32842
rect 12992 32778 13044 32784
rect 12900 31884 12952 31890
rect 12952 31844 13032 31872
rect 12900 31826 12952 31832
rect 12808 29300 12860 29306
rect 12808 29242 12860 29248
rect 12820 28694 12848 29242
rect 12808 28688 12860 28694
rect 12808 28630 12860 28636
rect 13004 28558 13032 31844
rect 13084 31748 13136 31754
rect 13084 31690 13136 31696
rect 13096 31482 13124 31690
rect 13084 31476 13136 31482
rect 13084 31418 13136 31424
rect 13096 30734 13124 31418
rect 13188 30734 13216 34478
rect 13084 30728 13136 30734
rect 13084 30670 13136 30676
rect 13176 30728 13228 30734
rect 13176 30670 13228 30676
rect 12532 28552 12584 28558
rect 12532 28494 12584 28500
rect 12992 28552 13044 28558
rect 12992 28494 13044 28500
rect 12440 28484 12492 28490
rect 12440 28426 12492 28432
rect 12452 28098 12480 28426
rect 12544 28218 12572 28494
rect 12900 28416 12952 28422
rect 12900 28358 12952 28364
rect 12532 28212 12584 28218
rect 12532 28154 12584 28160
rect 12716 28144 12768 28150
rect 12452 28082 12664 28098
rect 12716 28086 12768 28092
rect 12452 28076 12676 28082
rect 12452 28070 12624 28076
rect 12452 27674 12480 28070
rect 12624 28018 12676 28024
rect 12440 27668 12492 27674
rect 12440 27610 12492 27616
rect 12728 26994 12756 28086
rect 12912 27470 12940 28358
rect 13188 28082 13216 30670
rect 13280 30666 13308 34546
rect 13544 32836 13596 32842
rect 13544 32778 13596 32784
rect 13452 31884 13504 31890
rect 13452 31826 13504 31832
rect 13268 30660 13320 30666
rect 13268 30602 13320 30608
rect 13280 28150 13308 30602
rect 13464 29782 13492 31826
rect 13556 31482 13584 32778
rect 13544 31476 13596 31482
rect 13544 31418 13596 31424
rect 13452 29776 13504 29782
rect 13452 29718 13504 29724
rect 13360 29164 13412 29170
rect 13360 29106 13412 29112
rect 13372 28218 13400 29106
rect 13464 28490 13492 29718
rect 13452 28484 13504 28490
rect 13452 28426 13504 28432
rect 13360 28212 13412 28218
rect 13360 28154 13412 28160
rect 13268 28144 13320 28150
rect 13268 28086 13320 28092
rect 13176 28076 13228 28082
rect 13176 28018 13228 28024
rect 12900 27464 12952 27470
rect 12900 27406 12952 27412
rect 13188 26994 13216 28018
rect 12716 26988 12768 26994
rect 12716 26930 12768 26936
rect 13176 26988 13228 26994
rect 13176 26930 13228 26936
rect 12440 26920 12492 26926
rect 12440 26862 12492 26868
rect 12452 26382 12480 26862
rect 12440 26376 12492 26382
rect 12440 26318 12492 26324
rect 12348 24676 12400 24682
rect 12348 24618 12400 24624
rect 12256 23248 12308 23254
rect 12256 23190 12308 23196
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 12176 20806 12204 21490
rect 12348 20868 12400 20874
rect 12348 20810 12400 20816
rect 12164 20800 12216 20806
rect 12164 20742 12216 20748
rect 11980 20596 12032 20602
rect 11980 20538 12032 20544
rect 12176 20534 12204 20742
rect 12164 20528 12216 20534
rect 12164 20470 12216 20476
rect 12256 20392 12308 20398
rect 12256 20334 12308 20340
rect 11980 19372 12032 19378
rect 11980 19314 12032 19320
rect 11612 19168 11664 19174
rect 11612 19110 11664 19116
rect 11702 19136 11758 19145
rect 11624 18834 11652 19110
rect 11702 19071 11758 19080
rect 11612 18828 11664 18834
rect 11612 18770 11664 18776
rect 11624 18426 11652 18770
rect 11716 18766 11744 19071
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11612 18420 11664 18426
rect 11612 18362 11664 18368
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11624 16114 11652 17138
rect 11716 17066 11744 18702
rect 11900 18426 11928 18702
rect 11992 18426 12020 19314
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11980 18420 12032 18426
rect 11980 18362 12032 18368
rect 12072 17536 12124 17542
rect 12268 17524 12296 20334
rect 12360 18290 12388 20810
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 12124 17496 12296 17524
rect 12072 17478 12124 17484
rect 12084 17270 12112 17478
rect 12360 17270 12388 18226
rect 12072 17264 12124 17270
rect 12072 17206 12124 17212
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 11704 17060 11756 17066
rect 11704 17002 11756 17008
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11716 16096 11744 16526
rect 11980 16108 12032 16114
rect 11716 16068 11980 16096
rect 10876 15496 10928 15502
rect 10980 15473 11008 16050
rect 10876 15438 10928 15444
rect 10966 15464 11022 15473
rect 10888 13938 10916 15438
rect 10966 15399 11022 15408
rect 10980 15366 11008 15399
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10600 13524 10652 13530
rect 10600 13466 10652 13472
rect 10612 13258 10640 13466
rect 10600 13252 10652 13258
rect 10600 13194 10652 13200
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 10232 10464 10284 10470
rect 10230 10432 10232 10441
rect 10284 10432 10286 10441
rect 10230 10367 10286 10376
rect 10244 10062 10272 10367
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10520 9654 10548 12718
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10612 10062 10640 10134
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10508 9648 10560 9654
rect 10508 9590 10560 9596
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10600 9444 10652 9450
rect 10600 9386 10652 9392
rect 10612 8974 10640 9386
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 9586 8528 9642 8537
rect 9586 8463 9642 8472
rect 9692 8294 9720 8570
rect 9772 8560 9824 8566
rect 9770 8528 9772 8537
rect 9824 8528 9826 8537
rect 9770 8463 9826 8472
rect 9416 8266 9536 8294
rect 9508 7886 9536 8266
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9586 8120 9642 8129
rect 9586 8055 9588 8064
rect 9640 8055 9642 8064
rect 9588 8026 9640 8032
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9680 7880 9732 7886
rect 9784 7868 9812 8463
rect 9732 7840 9812 7868
rect 9680 7822 9732 7828
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9508 7546 9536 7686
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9232 6798 9260 7142
rect 9508 7041 9536 7346
rect 9772 7200 9824 7206
rect 9586 7168 9642 7177
rect 9772 7142 9824 7148
rect 9586 7103 9642 7112
rect 9494 7032 9550 7041
rect 9494 6967 9550 6976
rect 9496 6928 9548 6934
rect 9496 6870 9548 6876
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9232 5846 9260 6394
rect 9508 6322 9536 6870
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9232 5370 9260 5646
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9402 5128 9458 5137
rect 9402 5063 9458 5072
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 9128 3460 9180 3466
rect 9128 3402 9180 3408
rect 8576 3120 8628 3126
rect 8852 3120 8904 3126
rect 8576 3062 8628 3068
rect 8666 3088 8722 3097
rect 8852 3062 8904 3068
rect 8942 3088 8998 3097
rect 8666 3023 8668 3032
rect 8720 3023 8722 3032
rect 8668 2994 8720 3000
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8864 2774 8892 3062
rect 8942 3023 8944 3032
rect 8996 3023 8998 3032
rect 8944 2994 8996 3000
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 8772 2746 8892 2774
rect 8576 2576 8628 2582
rect 8576 2518 8628 2524
rect 8484 2372 8536 2378
rect 8484 2314 8536 2320
rect 8496 800 8524 2314
rect 8588 800 8616 2518
rect 8772 800 8800 2746
rect 8852 2304 8904 2310
rect 8852 2246 8904 2252
rect 8864 800 8892 2246
rect 9048 800 9076 2858
rect 9140 800 9168 3402
rect 9232 2854 9260 3878
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 9324 800 9352 4082
rect 9416 3670 9444 5063
rect 9494 4040 9550 4049
rect 9494 3975 9496 3984
rect 9548 3975 9550 3984
rect 9496 3946 9548 3952
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9404 2916 9456 2922
rect 9404 2858 9456 2864
rect 9416 800 9444 2858
rect 9508 1442 9536 3470
rect 9600 2446 9628 7103
rect 9784 4146 9812 7142
rect 10060 6186 10088 7754
rect 10152 7546 10180 8570
rect 10612 7954 10640 8910
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9876 4010 9904 4626
rect 9864 4004 9916 4010
rect 9864 3946 9916 3952
rect 9876 3738 9904 3946
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 9508 1414 9628 1442
rect 9600 800 9628 1414
rect 9692 800 9720 3606
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9784 3194 9812 3470
rect 9862 3360 9918 3369
rect 9862 3295 9918 3304
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9876 3058 9904 3295
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9968 800 9996 6054
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10140 5092 10192 5098
rect 10140 5034 10192 5040
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 10060 4486 10088 4762
rect 10152 4554 10180 5034
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 10060 2038 10088 4422
rect 10048 2032 10100 2038
rect 10048 1974 10100 1980
rect 10244 800 10272 5646
rect 10336 4826 10364 7482
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10324 4820 10376 4826
rect 10324 4762 10376 4768
rect 10336 4729 10364 4762
rect 10322 4720 10378 4729
rect 10322 4655 10378 4664
rect 10428 3126 10456 7142
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 10428 2854 10456 3062
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 10414 2680 10470 2689
rect 10414 2615 10416 2624
rect 10468 2615 10470 2624
rect 10416 2586 10468 2592
rect 10428 2378 10456 2586
rect 10416 2372 10468 2378
rect 10416 2314 10468 2320
rect 10520 800 10548 6054
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 3641 10640 3878
rect 10598 3632 10654 3641
rect 10598 3567 10654 3576
rect 10704 3534 10732 8298
rect 10796 7750 10824 9454
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10888 6662 10916 8434
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10796 800 10824 5646
rect 10888 2774 10916 6598
rect 10980 4826 11008 15302
rect 11716 14958 11744 16068
rect 11980 16050 12032 16056
rect 12084 15502 12112 17206
rect 12452 16250 12480 26318
rect 12624 26308 12676 26314
rect 12624 26250 12676 26256
rect 12636 25770 12664 26250
rect 12992 25900 13044 25906
rect 12992 25842 13044 25848
rect 12624 25764 12676 25770
rect 12624 25706 12676 25712
rect 13004 25702 13032 25842
rect 12992 25696 13044 25702
rect 12992 25638 13044 25644
rect 12716 25152 12768 25158
rect 12716 25094 12768 25100
rect 13452 25152 13504 25158
rect 13452 25094 13504 25100
rect 12624 24948 12676 24954
rect 12624 24890 12676 24896
rect 12636 24138 12664 24890
rect 12728 24818 12756 25094
rect 13464 24818 13492 25094
rect 12716 24812 12768 24818
rect 12716 24754 12768 24760
rect 12808 24812 12860 24818
rect 12808 24754 12860 24760
rect 13084 24812 13136 24818
rect 13084 24754 13136 24760
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 12820 24682 12848 24754
rect 12808 24676 12860 24682
rect 12808 24618 12860 24624
rect 12900 24200 12952 24206
rect 12900 24142 12952 24148
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 12912 23662 12940 24142
rect 13096 23866 13124 24754
rect 13464 23866 13492 24754
rect 13544 24064 13596 24070
rect 13544 24006 13596 24012
rect 13084 23860 13136 23866
rect 13084 23802 13136 23808
rect 13452 23860 13504 23866
rect 13452 23802 13504 23808
rect 13556 23730 13584 24006
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 12900 23656 12952 23662
rect 13648 23610 13676 44814
rect 16028 42016 16080 42022
rect 16028 41958 16080 41964
rect 14740 41744 14792 41750
rect 14740 41686 14792 41692
rect 13912 41676 13964 41682
rect 13912 41618 13964 41624
rect 13924 41070 13952 41618
rect 14752 41614 14780 41686
rect 16040 41614 16068 41958
rect 14556 41608 14608 41614
rect 14556 41550 14608 41556
rect 14740 41608 14792 41614
rect 14740 41550 14792 41556
rect 16028 41608 16080 41614
rect 16028 41550 16080 41556
rect 14096 41472 14148 41478
rect 14096 41414 14148 41420
rect 13912 41064 13964 41070
rect 13912 41006 13964 41012
rect 13728 40928 13780 40934
rect 13728 40870 13780 40876
rect 13740 39370 13768 40870
rect 13924 40594 13952 41006
rect 13912 40588 13964 40594
rect 13912 40530 13964 40536
rect 13820 40520 13872 40526
rect 13820 40462 13872 40468
rect 13832 39846 13860 40462
rect 14108 40050 14136 41414
rect 14372 41132 14424 41138
rect 14372 41074 14424 41080
rect 14188 40996 14240 41002
rect 14188 40938 14240 40944
rect 14200 40594 14228 40938
rect 14384 40594 14412 41074
rect 14568 40730 14596 41550
rect 14752 41138 14780 41550
rect 15292 41472 15344 41478
rect 15292 41414 15344 41420
rect 14740 41132 14792 41138
rect 14740 41074 14792 41080
rect 15016 41132 15068 41138
rect 15016 41074 15068 41080
rect 14556 40724 14608 40730
rect 14556 40666 14608 40672
rect 14188 40588 14240 40594
rect 14188 40530 14240 40536
rect 14372 40588 14424 40594
rect 14372 40530 14424 40536
rect 14096 40044 14148 40050
rect 14096 39986 14148 39992
rect 13820 39840 13872 39846
rect 13820 39782 13872 39788
rect 13728 39364 13780 39370
rect 13728 39306 13780 39312
rect 13832 38758 13860 39782
rect 14096 39636 14148 39642
rect 14096 39578 14148 39584
rect 13820 38752 13872 38758
rect 13820 38694 13872 38700
rect 13832 36106 13860 38694
rect 14004 36780 14056 36786
rect 14004 36722 14056 36728
rect 14016 36378 14044 36722
rect 14004 36372 14056 36378
rect 14004 36314 14056 36320
rect 13820 36100 13872 36106
rect 13820 36042 13872 36048
rect 14004 36032 14056 36038
rect 14004 35974 14056 35980
rect 14016 35562 14044 35974
rect 14004 35556 14056 35562
rect 14004 35498 14056 35504
rect 13912 35488 13964 35494
rect 13912 35430 13964 35436
rect 13924 33590 13952 35430
rect 13912 33584 13964 33590
rect 13912 33526 13964 33532
rect 14016 32570 14044 35498
rect 14108 35018 14136 39578
rect 14200 39438 14228 40530
rect 15028 39642 15056 41074
rect 15200 40656 15252 40662
rect 15200 40598 15252 40604
rect 15108 40384 15160 40390
rect 15108 40326 15160 40332
rect 15016 39636 15068 39642
rect 15016 39578 15068 39584
rect 14188 39432 14240 39438
rect 14188 39374 14240 39380
rect 14648 37188 14700 37194
rect 14648 37130 14700 37136
rect 14556 37120 14608 37126
rect 14556 37062 14608 37068
rect 14372 36372 14424 36378
rect 14372 36314 14424 36320
rect 14384 36174 14412 36314
rect 14568 36174 14596 37062
rect 14660 36922 14688 37130
rect 14648 36916 14700 36922
rect 14648 36858 14700 36864
rect 15120 36378 15148 40326
rect 15212 39642 15240 40598
rect 15200 39636 15252 39642
rect 15200 39578 15252 39584
rect 15108 36372 15160 36378
rect 15108 36314 15160 36320
rect 14372 36168 14424 36174
rect 14372 36110 14424 36116
rect 14556 36168 14608 36174
rect 14556 36110 14608 36116
rect 14740 36168 14792 36174
rect 14740 36110 14792 36116
rect 14280 36100 14332 36106
rect 14280 36042 14332 36048
rect 14096 35012 14148 35018
rect 14096 34954 14148 34960
rect 14292 34134 14320 36042
rect 14752 35494 14780 36110
rect 14740 35488 14792 35494
rect 14740 35430 14792 35436
rect 15108 34944 15160 34950
rect 15108 34886 15160 34892
rect 14556 34400 14608 34406
rect 14556 34342 14608 34348
rect 14568 34241 14596 34342
rect 14554 34232 14610 34241
rect 15120 34202 15148 34886
rect 14554 34167 14556 34176
rect 14608 34167 14610 34176
rect 15108 34196 15160 34202
rect 14556 34138 14608 34144
rect 15108 34138 15160 34144
rect 14280 34128 14332 34134
rect 14280 34070 14332 34076
rect 14924 33992 14976 33998
rect 14924 33934 14976 33940
rect 14648 33924 14700 33930
rect 14648 33866 14700 33872
rect 14004 32564 14056 32570
rect 14004 32506 14056 32512
rect 13820 32224 13872 32230
rect 13820 32166 13872 32172
rect 13832 30734 13860 32166
rect 14556 32020 14608 32026
rect 14556 31962 14608 31968
rect 14568 31822 14596 31962
rect 14556 31816 14608 31822
rect 14556 31758 14608 31764
rect 14096 31680 14148 31686
rect 14096 31622 14148 31628
rect 14108 31414 14136 31622
rect 14096 31408 14148 31414
rect 14096 31350 14148 31356
rect 14660 31210 14688 33866
rect 14936 33590 14964 33934
rect 15304 33640 15332 41414
rect 15384 40520 15436 40526
rect 15384 40462 15436 40468
rect 15396 39982 15424 40462
rect 15384 39976 15436 39982
rect 15384 39918 15436 39924
rect 15396 39846 15424 39918
rect 15384 39840 15436 39846
rect 15384 39782 15436 39788
rect 15396 39506 15424 39782
rect 15384 39500 15436 39506
rect 15384 39442 15436 39448
rect 15396 37262 15424 39442
rect 16120 38344 16172 38350
rect 16120 38286 16172 38292
rect 15936 38276 15988 38282
rect 15936 38218 15988 38224
rect 15948 38010 15976 38218
rect 15936 38004 15988 38010
rect 15936 37946 15988 37952
rect 16132 37874 16160 38286
rect 16120 37868 16172 37874
rect 16120 37810 16172 37816
rect 15384 37256 15436 37262
rect 15384 37198 15436 37204
rect 15396 36786 15424 37198
rect 15476 37188 15528 37194
rect 15476 37130 15528 37136
rect 15488 36922 15516 37130
rect 15476 36916 15528 36922
rect 15476 36858 15528 36864
rect 15384 36780 15436 36786
rect 15384 36722 15436 36728
rect 15732 36780 15784 36786
rect 16120 36780 16172 36786
rect 15784 36728 15792 36768
rect 15732 36722 15792 36728
rect 16120 36722 16172 36728
rect 15396 35154 15424 36722
rect 15476 36576 15528 36582
rect 15476 36518 15528 36524
rect 15384 35148 15436 35154
rect 15384 35090 15436 35096
rect 15304 33612 15424 33640
rect 14924 33584 14976 33590
rect 14924 33526 14976 33532
rect 15016 33516 15068 33522
rect 15016 33458 15068 33464
rect 15292 33516 15344 33522
rect 15292 33458 15344 33464
rect 15028 32774 15056 33458
rect 15304 33114 15332 33458
rect 15292 33108 15344 33114
rect 15292 33050 15344 33056
rect 15016 32768 15068 32774
rect 15016 32710 15068 32716
rect 14740 32564 14792 32570
rect 15028 32552 15056 32710
rect 14740 32506 14792 32512
rect 14936 32524 15056 32552
rect 14752 31822 14780 32506
rect 14936 32434 14964 32524
rect 14924 32428 14976 32434
rect 14924 32370 14976 32376
rect 15016 32428 15068 32434
rect 15016 32370 15068 32376
rect 14740 31816 14792 31822
rect 14740 31758 14792 31764
rect 14924 31340 14976 31346
rect 14924 31282 14976 31288
rect 13912 31204 13964 31210
rect 13912 31146 13964 31152
rect 14648 31204 14700 31210
rect 14648 31146 14700 31152
rect 13820 30728 13872 30734
rect 13820 30670 13872 30676
rect 13820 29164 13872 29170
rect 13924 29152 13952 31146
rect 14936 30938 14964 31282
rect 14924 30932 14976 30938
rect 14924 30874 14976 30880
rect 14280 30728 14332 30734
rect 14280 30670 14332 30676
rect 14292 30122 14320 30670
rect 15028 30258 15056 32370
rect 15396 32366 15424 33612
rect 15488 33522 15516 36518
rect 15764 36378 15792 36722
rect 15844 36644 15896 36650
rect 15844 36586 15896 36592
rect 15752 36372 15804 36378
rect 15752 36314 15804 36320
rect 15856 36106 15884 36586
rect 16132 36582 16160 36722
rect 16120 36576 16172 36582
rect 16120 36518 16172 36524
rect 15844 36100 15896 36106
rect 15844 36042 15896 36048
rect 16120 34740 16172 34746
rect 16120 34682 16172 34688
rect 15936 33856 15988 33862
rect 15936 33798 15988 33804
rect 15948 33590 15976 33798
rect 15936 33584 15988 33590
rect 15936 33526 15988 33532
rect 15476 33516 15528 33522
rect 15476 33458 15528 33464
rect 16132 32910 16160 34682
rect 16120 32904 16172 32910
rect 16120 32846 16172 32852
rect 16028 32836 16080 32842
rect 16028 32778 16080 32784
rect 15384 32360 15436 32366
rect 15384 32302 15436 32308
rect 15568 31748 15620 31754
rect 15568 31690 15620 31696
rect 15384 31476 15436 31482
rect 15384 31418 15436 31424
rect 15200 31272 15252 31278
rect 15200 31214 15252 31220
rect 15212 30734 15240 31214
rect 15200 30728 15252 30734
rect 15200 30670 15252 30676
rect 15200 30592 15252 30598
rect 15200 30534 15252 30540
rect 15212 30258 15240 30534
rect 14556 30252 14608 30258
rect 14556 30194 14608 30200
rect 15016 30252 15068 30258
rect 15016 30194 15068 30200
rect 15200 30252 15252 30258
rect 15200 30194 15252 30200
rect 14280 30116 14332 30122
rect 14280 30058 14332 30064
rect 14292 29170 14320 30058
rect 14372 29232 14424 29238
rect 14372 29174 14424 29180
rect 13872 29124 13952 29152
rect 14280 29164 14332 29170
rect 13820 29106 13872 29112
rect 14280 29106 14332 29112
rect 13832 26586 13860 29106
rect 13912 28484 13964 28490
rect 13912 28426 13964 28432
rect 13924 28218 13952 28426
rect 14384 28218 14412 29174
rect 14568 28558 14596 30194
rect 14740 30048 14792 30054
rect 14740 29990 14792 29996
rect 14556 28552 14608 28558
rect 14556 28494 14608 28500
rect 13912 28212 13964 28218
rect 13912 28154 13964 28160
rect 14372 28212 14424 28218
rect 14372 28154 14424 28160
rect 13820 26580 13872 26586
rect 13820 26522 13872 26528
rect 13924 25974 13952 28154
rect 14004 26240 14056 26246
rect 14004 26182 14056 26188
rect 13912 25968 13964 25974
rect 13912 25910 13964 25916
rect 13728 25288 13780 25294
rect 13728 25230 13780 25236
rect 13740 23730 13768 25230
rect 13820 24608 13872 24614
rect 13820 24550 13872 24556
rect 13832 24206 13860 24550
rect 13820 24200 13872 24206
rect 13820 24142 13872 24148
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 12900 23598 12952 23604
rect 13556 23582 13676 23610
rect 12624 21888 12676 21894
rect 12624 21830 12676 21836
rect 12532 20460 12584 20466
rect 12532 20402 12584 20408
rect 12544 20058 12572 20402
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12544 18290 12572 18906
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 12176 15026 12204 16186
rect 12544 15706 12572 17138
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12544 15094 12572 15642
rect 12532 15088 12584 15094
rect 12532 15030 12584 15036
rect 12636 15026 12664 21830
rect 13176 21140 13228 21146
rect 13176 21082 13228 21088
rect 13084 20800 13136 20806
rect 13084 20742 13136 20748
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 12728 19174 12756 19858
rect 13096 19854 13124 20742
rect 13188 19854 13216 21082
rect 13268 21072 13320 21078
rect 13268 21014 13320 21020
rect 13280 20806 13308 21014
rect 13268 20800 13320 20806
rect 13268 20742 13320 20748
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13280 19922 13308 20402
rect 13268 19916 13320 19922
rect 13268 19858 13320 19864
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12728 18358 12756 19110
rect 12716 18352 12768 18358
rect 12716 18294 12768 18300
rect 12728 17882 12756 18294
rect 13188 18290 13216 19790
rect 13176 18284 13228 18290
rect 13228 18244 13492 18272
rect 13176 18226 13228 18232
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 12992 17808 13044 17814
rect 12992 17750 13044 17756
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12728 16658 12756 17546
rect 13004 17542 13032 17750
rect 13464 17678 13492 18244
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 12808 17536 12860 17542
rect 12808 17478 12860 17484
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12728 16114 12756 16390
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12728 15978 12756 16050
rect 12716 15972 12768 15978
rect 12716 15914 12768 15920
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11348 13394 11376 14894
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11992 13938 12020 14350
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 11992 12714 12020 13874
rect 12176 13682 12204 13874
rect 12176 13654 12296 13682
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 11980 12708 12032 12714
rect 11980 12650 12032 12656
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 11072 12238 11100 12582
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11992 11762 12020 12650
rect 12176 12374 12204 12786
rect 12164 12368 12216 12374
rect 12164 12310 12216 12316
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11532 11150 11560 11630
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11532 9994 11560 11086
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11886 9344 11942 9353
rect 11716 9042 11744 9318
rect 11886 9279 11942 9288
rect 11794 9072 11850 9081
rect 11704 9036 11756 9042
rect 11900 9042 11928 9279
rect 12268 9110 12296 13654
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12452 11354 12480 12242
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 9994 12480 10406
rect 12440 9988 12492 9994
rect 12440 9930 12492 9936
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 11794 9007 11850 9016
rect 11888 9036 11940 9042
rect 11704 8978 11756 8984
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11256 7206 11284 8910
rect 11808 8430 11836 9007
rect 11888 8978 11940 8984
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 11888 8900 11940 8906
rect 11888 8842 11940 8848
rect 11900 8498 11928 8842
rect 12268 8537 12296 8910
rect 12254 8528 12310 8537
rect 11888 8492 11940 8498
rect 12254 8463 12256 8472
rect 11888 8434 11940 8440
rect 12308 8463 12310 8472
rect 12256 8434 12308 8440
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 11072 3602 11100 6122
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 11060 3596 11112 3602
rect 11060 3538 11112 3544
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 10980 2961 11008 2994
rect 10966 2952 11022 2961
rect 10966 2887 11022 2896
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 10888 2746 11008 2774
rect 10980 2514 11008 2746
rect 11072 2650 11100 2858
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 11164 1170 11192 5034
rect 11256 3534 11284 7142
rect 11624 6798 11652 8298
rect 11992 8090 12020 8366
rect 12452 8265 12480 9930
rect 12636 9586 12664 10610
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12728 9178 12756 15914
rect 12820 15434 12848 17478
rect 13280 17338 13308 17614
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 12992 16720 13044 16726
rect 12992 16662 13044 16668
rect 13004 16114 13032 16662
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12912 15314 12940 15982
rect 13004 15366 13032 16050
rect 12820 15286 12940 15314
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 12820 15094 12848 15286
rect 12808 15088 12860 15094
rect 12808 15030 12860 15036
rect 13004 12434 13032 15302
rect 12912 12406 13032 12434
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12820 10062 12848 10406
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12820 9586 12848 9862
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12438 8256 12494 8265
rect 12438 8191 12494 8200
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11072 1142 11192 1170
rect 11072 800 11100 1142
rect 11348 800 11376 5646
rect 11428 5228 11480 5234
rect 11428 5170 11480 5176
rect 11440 4758 11468 5170
rect 11796 5160 11848 5166
rect 11796 5102 11848 5108
rect 11704 5092 11756 5098
rect 11704 5034 11756 5040
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11428 4752 11480 4758
rect 11428 4694 11480 4700
rect 11440 4622 11468 4694
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11440 4078 11468 4558
rect 11532 4486 11560 4626
rect 11520 4480 11572 4486
rect 11520 4422 11572 4428
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11518 4040 11574 4049
rect 11518 3975 11574 3984
rect 11532 3058 11560 3975
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 11532 1970 11560 2382
rect 11520 1964 11572 1970
rect 11520 1906 11572 1912
rect 11624 800 11652 4966
rect 11716 4826 11744 5034
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 11716 4078 11744 4762
rect 11808 4622 11836 5102
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11808 3942 11836 4558
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11900 800 11928 5646
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11992 4486 12020 4966
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11992 4010 12020 4422
rect 11980 4004 12032 4010
rect 11980 3946 12032 3952
rect 12084 3534 12112 7686
rect 12728 7478 12756 8774
rect 12808 8560 12860 8566
rect 12808 8502 12860 8508
rect 12820 8430 12848 8502
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 12716 7472 12768 7478
rect 12716 7414 12768 7420
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 12084 2922 12112 3470
rect 12072 2916 12124 2922
rect 12072 2858 12124 2864
rect 12176 800 12204 6054
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12254 4720 12310 4729
rect 12254 4655 12256 4664
rect 12308 4655 12310 4664
rect 12256 4626 12308 4632
rect 12452 800 12480 5646
rect 12728 800 12756 5646
rect 12912 4078 12940 12406
rect 13280 12306 13308 17070
rect 13360 16176 13412 16182
rect 13360 16118 13412 16124
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13372 12170 13400 16118
rect 13556 12434 13584 23582
rect 13636 23520 13688 23526
rect 13636 23462 13688 23468
rect 13648 21146 13676 23462
rect 13740 23118 13768 23666
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 13820 22772 13872 22778
rect 13820 22714 13872 22720
rect 13636 21140 13688 21146
rect 13636 21082 13688 21088
rect 13728 21072 13780 21078
rect 13728 21014 13780 21020
rect 13636 21004 13688 21010
rect 13636 20946 13688 20952
rect 13648 20874 13676 20946
rect 13636 20868 13688 20874
rect 13636 20810 13688 20816
rect 13648 20602 13676 20810
rect 13636 20596 13688 20602
rect 13636 20538 13688 20544
rect 13740 20534 13768 21014
rect 13728 20528 13780 20534
rect 13728 20470 13780 20476
rect 13728 19780 13780 19786
rect 13728 19722 13780 19728
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13648 18290 13676 18906
rect 13740 18834 13768 19722
rect 13832 19446 13860 22714
rect 14016 22094 14044 26182
rect 14188 25696 14240 25702
rect 14188 25638 14240 25644
rect 14200 25158 14228 25638
rect 14188 25152 14240 25158
rect 14188 25094 14240 25100
rect 14016 22066 14136 22094
rect 14108 22030 14136 22066
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 14096 20392 14148 20398
rect 14096 20334 14148 20340
rect 14108 19514 14136 20334
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 13820 19440 13872 19446
rect 13820 19382 13872 19388
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13924 18358 13952 19246
rect 13912 18352 13964 18358
rect 13912 18294 13964 18300
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 13912 18148 13964 18154
rect 13912 18090 13964 18096
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13636 17740 13688 17746
rect 13636 17682 13688 17688
rect 13648 15502 13676 17682
rect 13832 17678 13860 18022
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13924 17338 13952 18090
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 14108 17338 14136 17478
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 14096 17332 14148 17338
rect 14096 17274 14148 17280
rect 13912 16516 13964 16522
rect 13912 16458 13964 16464
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13832 15570 13860 15846
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 13924 15416 13952 16458
rect 14004 15496 14056 15502
rect 14004 15438 14056 15444
rect 13464 12406 13584 12434
rect 13832 15388 13952 15416
rect 13360 12164 13412 12170
rect 13360 12106 13412 12112
rect 13372 11354 13400 12106
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 13280 9450 13308 9862
rect 13268 9444 13320 9450
rect 13268 9386 13320 9392
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 13096 8974 13124 9318
rect 13280 9178 13308 9386
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 13358 8664 13414 8673
rect 13358 8599 13360 8608
rect 13412 8599 13414 8608
rect 13360 8570 13412 8576
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13084 6724 13136 6730
rect 13084 6666 13136 6672
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 13004 800 13032 5714
rect 13096 3058 13124 6666
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 13280 5914 13308 6190
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 13188 2446 13216 5578
rect 13372 3534 13400 7822
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 13188 1902 13216 2382
rect 13176 1896 13228 1902
rect 13176 1838 13228 1844
rect 13280 800 13308 3470
rect 13464 2650 13492 12406
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 13556 800 13584 4966
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13648 3194 13676 3470
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13740 2774 13768 12310
rect 13832 11762 13860 15388
rect 14016 15314 14044 15438
rect 13924 15286 14044 15314
rect 13924 15026 13952 15286
rect 14004 15088 14056 15094
rect 14004 15030 14056 15036
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 13924 14822 13952 14962
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13924 8650 13952 14758
rect 14016 14074 14044 15030
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 14016 13326 14044 14010
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 14096 13252 14148 13258
rect 14096 13194 14148 13200
rect 14108 12238 14136 13194
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 14108 11830 14136 12174
rect 14096 11824 14148 11830
rect 14096 11766 14148 11772
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 14016 10810 14044 11698
rect 14200 11014 14228 25094
rect 14568 24954 14596 28494
rect 14752 28370 14780 29990
rect 15396 29102 15424 31418
rect 15476 31408 15528 31414
rect 15476 31350 15528 31356
rect 15488 30938 15516 31350
rect 15476 30932 15528 30938
rect 15476 30874 15528 30880
rect 15580 30122 15608 31690
rect 15844 31680 15896 31686
rect 15844 31622 15896 31628
rect 15752 30728 15804 30734
rect 15752 30670 15804 30676
rect 15660 30660 15712 30666
rect 15660 30602 15712 30608
rect 15672 30326 15700 30602
rect 15660 30320 15712 30326
rect 15660 30262 15712 30268
rect 15568 30116 15620 30122
rect 15568 30058 15620 30064
rect 15384 29096 15436 29102
rect 15384 29038 15436 29044
rect 14924 29028 14976 29034
rect 14924 28970 14976 28976
rect 14832 28960 14884 28966
rect 14832 28902 14884 28908
rect 14844 28558 14872 28902
rect 14832 28552 14884 28558
rect 14832 28494 14884 28500
rect 14752 28342 14872 28370
rect 14740 27940 14792 27946
rect 14740 27882 14792 27888
rect 14752 27470 14780 27882
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 14740 25152 14792 25158
rect 14740 25094 14792 25100
rect 14556 24948 14608 24954
rect 14556 24890 14608 24896
rect 14280 24812 14332 24818
rect 14280 24754 14332 24760
rect 14292 24342 14320 24754
rect 14280 24336 14332 24342
rect 14280 24278 14332 24284
rect 14752 24206 14780 25094
rect 14740 24200 14792 24206
rect 14740 24142 14792 24148
rect 14556 24064 14608 24070
rect 14556 24006 14608 24012
rect 14568 22710 14596 24006
rect 14844 23746 14872 28342
rect 14936 25514 14964 28970
rect 15580 28762 15608 30058
rect 15568 28756 15620 28762
rect 15568 28698 15620 28704
rect 15200 28484 15252 28490
rect 15200 28426 15252 28432
rect 15212 28082 15240 28426
rect 15292 28416 15344 28422
rect 15292 28358 15344 28364
rect 15304 28150 15332 28358
rect 15292 28144 15344 28150
rect 15292 28086 15344 28092
rect 15764 28082 15792 30670
rect 15856 30258 15884 31622
rect 16040 31482 16068 32778
rect 16120 32768 16172 32774
rect 16120 32710 16172 32716
rect 16028 31476 16080 31482
rect 16028 31418 16080 31424
rect 16028 31136 16080 31142
rect 16028 31078 16080 31084
rect 15844 30252 15896 30258
rect 15844 30194 15896 30200
rect 15856 29782 15884 30194
rect 15844 29776 15896 29782
rect 15844 29718 15896 29724
rect 15844 29300 15896 29306
rect 15844 29242 15896 29248
rect 15856 28558 15884 29242
rect 15844 28552 15896 28558
rect 15844 28494 15896 28500
rect 15200 28076 15252 28082
rect 15200 28018 15252 28024
rect 15752 28076 15804 28082
rect 15752 28018 15804 28024
rect 15108 25832 15160 25838
rect 15108 25774 15160 25780
rect 14936 25486 15056 25514
rect 14924 24880 14976 24886
rect 14924 24822 14976 24828
rect 14936 24206 14964 24822
rect 14924 24200 14976 24206
rect 14924 24142 14976 24148
rect 14936 23866 14964 24142
rect 14924 23860 14976 23866
rect 14924 23802 14976 23808
rect 14844 23718 14964 23746
rect 14556 22704 14608 22710
rect 14556 22646 14608 22652
rect 14832 22636 14884 22642
rect 14832 22578 14884 22584
rect 14280 22432 14332 22438
rect 14280 22374 14332 22380
rect 14292 18290 14320 22374
rect 14844 22166 14872 22578
rect 14832 22160 14884 22166
rect 14832 22102 14884 22108
rect 14936 21894 14964 23718
rect 14924 21888 14976 21894
rect 14924 21830 14976 21836
rect 14936 21486 14964 21830
rect 14924 21480 14976 21486
rect 14924 21422 14976 21428
rect 14464 21344 14516 21350
rect 14464 21286 14516 21292
rect 14648 21344 14700 21350
rect 14648 21286 14700 21292
rect 14476 20874 14504 21286
rect 14660 20942 14688 21286
rect 14648 20936 14700 20942
rect 14648 20878 14700 20884
rect 14464 20868 14516 20874
rect 14464 20810 14516 20816
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14384 17542 14412 18226
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14384 17202 14412 17478
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14476 17134 14504 20810
rect 14832 19848 14884 19854
rect 14830 19816 14832 19825
rect 14884 19816 14886 19825
rect 14830 19751 14886 19760
rect 14556 19304 14608 19310
rect 14556 19246 14608 19252
rect 14568 18290 14596 19246
rect 14556 18284 14608 18290
rect 14740 18284 14792 18290
rect 14556 18226 14608 18232
rect 14660 18244 14740 18272
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14292 15706 14320 16050
rect 14568 16046 14596 18226
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14660 14958 14688 18244
rect 14740 18226 14792 18232
rect 14936 18170 14964 21422
rect 15028 20058 15056 25486
rect 15120 24954 15148 25774
rect 15292 25696 15344 25702
rect 15292 25638 15344 25644
rect 15304 25294 15332 25638
rect 15292 25288 15344 25294
rect 15292 25230 15344 25236
rect 15200 25220 15252 25226
rect 15200 25162 15252 25168
rect 15212 24954 15240 25162
rect 15108 24948 15160 24954
rect 15108 24890 15160 24896
rect 15200 24948 15252 24954
rect 15200 24890 15252 24896
rect 15120 24138 15148 24890
rect 15108 24132 15160 24138
rect 15108 24074 15160 24080
rect 15212 23798 15240 24890
rect 15476 24608 15528 24614
rect 15476 24550 15528 24556
rect 15292 24064 15344 24070
rect 15292 24006 15344 24012
rect 15200 23792 15252 23798
rect 15200 23734 15252 23740
rect 15304 23730 15332 24006
rect 15108 23724 15160 23730
rect 15108 23666 15160 23672
rect 15292 23724 15344 23730
rect 15292 23666 15344 23672
rect 15120 22778 15148 23666
rect 15108 22772 15160 22778
rect 15108 22714 15160 22720
rect 15304 22642 15332 23666
rect 15488 23662 15516 24550
rect 15476 23656 15528 23662
rect 15476 23598 15528 23604
rect 15660 23656 15712 23662
rect 15660 23598 15712 23604
rect 15384 23520 15436 23526
rect 15384 23462 15436 23468
rect 15292 22636 15344 22642
rect 15292 22578 15344 22584
rect 15396 20942 15424 23462
rect 15488 22982 15516 23598
rect 15476 22976 15528 22982
rect 15476 22918 15528 22924
rect 15476 21548 15528 21554
rect 15476 21490 15528 21496
rect 15384 20936 15436 20942
rect 15384 20878 15436 20884
rect 15488 20466 15516 21490
rect 15672 20942 15700 23598
rect 15752 22432 15804 22438
rect 15752 22374 15804 22380
rect 15764 22030 15792 22374
rect 15752 22024 15804 22030
rect 15752 21966 15804 21972
rect 15764 21026 15792 21966
rect 15764 20998 15976 21026
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15672 20602 15700 20878
rect 15752 20868 15804 20874
rect 15752 20810 15804 20816
rect 15660 20596 15712 20602
rect 15660 20538 15712 20544
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 15016 20052 15068 20058
rect 15016 19994 15068 20000
rect 15016 19712 15068 19718
rect 15016 19654 15068 19660
rect 14752 18142 14964 18170
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14292 12986 14320 13874
rect 14660 13870 14688 14894
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14752 13682 14780 18142
rect 14936 18086 14964 18142
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14936 16114 14964 17070
rect 14924 16108 14976 16114
rect 14924 16050 14976 16056
rect 15028 15994 15056 19654
rect 15212 17202 15240 20402
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 14384 13654 14780 13682
rect 14844 15966 15056 15994
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14384 12186 14412 13654
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14660 12850 14688 13126
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 14476 12434 14504 12786
rect 14844 12442 14872 15966
rect 15108 15496 15160 15502
rect 15108 15438 15160 15444
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14936 14006 14964 14554
rect 15120 14414 15148 15438
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 15108 14408 15160 14414
rect 15108 14350 15160 14356
rect 14924 14000 14976 14006
rect 14924 13942 14976 13948
rect 15120 13938 15148 14350
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 14924 12776 14976 12782
rect 14924 12718 14976 12724
rect 14832 12436 14884 12442
rect 14476 12406 14688 12434
rect 14384 12158 14596 12186
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14292 11830 14320 12038
rect 14280 11824 14332 11830
rect 14280 11766 14332 11772
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 14004 10804 14056 10810
rect 14004 10746 14056 10752
rect 14384 10742 14412 12038
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14476 11150 14504 11494
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14372 10736 14424 10742
rect 14372 10678 14424 10684
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 13924 8622 14228 8650
rect 14292 8634 14320 9114
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 14476 8634 14504 9046
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 13912 7812 13964 7818
rect 13912 7754 13964 7760
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13832 6866 13860 7278
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13648 2746 13768 2774
rect 13648 2514 13676 2746
rect 13636 2508 13688 2514
rect 13636 2450 13688 2456
rect 13832 800 13860 6122
rect 13924 2446 13952 7754
rect 14016 6866 14044 8434
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 14016 5234 14044 6802
rect 14200 5370 14228 8622
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14292 7410 14320 7822
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 14292 4622 14320 7142
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14016 2774 14044 4558
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14108 3233 14136 3334
rect 14094 3224 14150 3233
rect 14094 3159 14150 3168
rect 14016 2746 14136 2774
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 14108 800 14136 2746
rect 14200 800 14228 3538
rect 14384 800 14412 4966
rect 14476 3058 14504 7890
rect 14568 7546 14596 12158
rect 14660 9160 14688 12406
rect 14832 12378 14884 12384
rect 14832 12232 14884 12238
rect 14752 12180 14832 12186
rect 14752 12174 14884 12180
rect 14752 12158 14872 12174
rect 14936 12170 14964 12718
rect 15120 12238 15148 12786
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 14924 12164 14976 12170
rect 14752 11898 14780 12158
rect 14976 12124 15056 12152
rect 14924 12106 14976 12112
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14844 11234 14872 12038
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 14936 11762 14964 11834
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 15028 11694 15056 12124
rect 15120 11762 15148 12174
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15016 11688 15068 11694
rect 15016 11630 15068 11636
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 14844 11206 14964 11234
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14740 9172 14792 9178
rect 14660 9132 14740 9160
rect 14740 9114 14792 9120
rect 14844 8650 14872 11018
rect 14752 8622 14872 8650
rect 14752 8401 14780 8622
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 14738 8392 14794 8401
rect 14738 8327 14794 8336
rect 14752 7886 14780 8327
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14568 7206 14596 7482
rect 14844 7342 14872 8434
rect 14936 7750 14964 11206
rect 15028 9722 15056 11494
rect 15212 10198 15240 14758
rect 15304 14278 15332 17138
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15396 15502 15424 16390
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 15764 12986 15792 20810
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15856 18766 15884 18906
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15856 16250 15884 16526
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15948 14346 15976 20998
rect 16040 17746 16068 31078
rect 16132 30326 16160 32710
rect 16120 30320 16172 30326
rect 16120 30262 16172 30268
rect 16120 29028 16172 29034
rect 16120 28970 16172 28976
rect 16132 22506 16160 28970
rect 16120 22500 16172 22506
rect 16120 22442 16172 22448
rect 16132 21962 16160 22442
rect 16120 21956 16172 21962
rect 16120 21898 16172 21904
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 16028 15428 16080 15434
rect 16028 15370 16080 15376
rect 16040 14822 16068 15370
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15488 11150 15516 12174
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15672 11218 15700 11698
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15476 11144 15528 11150
rect 15396 11092 15476 11098
rect 15396 11086 15528 11092
rect 15396 11070 15516 11086
rect 15396 10606 15424 11070
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15200 10192 15252 10198
rect 15200 10134 15252 10140
rect 15016 9716 15068 9722
rect 15016 9658 15068 9664
rect 15212 9450 15240 10134
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15200 9444 15252 9450
rect 15200 9386 15252 9392
rect 15016 8492 15068 8498
rect 15016 8434 15068 8440
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14752 6322 14780 6598
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14844 5710 14872 7278
rect 14936 6934 14964 7686
rect 15028 7546 15056 8434
rect 15108 8016 15160 8022
rect 15108 7958 15160 7964
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 14924 6928 14976 6934
rect 14924 6870 14976 6876
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14556 5636 14608 5642
rect 14556 5578 14608 5584
rect 14568 5370 14596 5578
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 14554 3224 14610 3233
rect 14554 3159 14556 3168
rect 14608 3159 14610 3168
rect 14556 3130 14608 3136
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 14476 800 14504 2858
rect 14554 2680 14610 2689
rect 14554 2615 14556 2624
rect 14608 2615 14610 2624
rect 14556 2586 14608 2592
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14568 2106 14596 2382
rect 14556 2100 14608 2106
rect 14556 2042 14608 2048
rect 14660 800 14688 4014
rect 14752 800 14780 4558
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14844 3466 14872 4422
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14936 800 14964 6734
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 15028 800 15056 2926
rect 15120 2854 15148 7958
rect 15212 6390 15240 9386
rect 15304 7410 15332 9454
rect 15396 8974 15424 10542
rect 15476 10532 15528 10538
rect 15476 10474 15528 10480
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15488 8566 15516 10474
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15580 9353 15608 9998
rect 15660 9376 15712 9382
rect 15566 9344 15622 9353
rect 15660 9318 15712 9324
rect 15566 9279 15622 9288
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15304 6662 15332 7346
rect 15384 7268 15436 7274
rect 15384 7210 15436 7216
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15304 5574 15332 6054
rect 15396 5642 15424 7210
rect 15488 5914 15516 7686
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15384 5636 15436 5642
rect 15384 5578 15436 5584
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15396 5370 15424 5578
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15292 4004 15344 4010
rect 15292 3946 15344 3952
rect 15198 3224 15254 3233
rect 15198 3159 15200 3168
rect 15252 3159 15254 3168
rect 15200 3130 15252 3136
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 15120 2446 15148 2790
rect 15304 2774 15332 3946
rect 15212 2746 15332 2774
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 15212 800 15240 2746
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 15304 2038 15332 2246
rect 15292 2032 15344 2038
rect 15292 1974 15344 1980
rect 15292 1896 15344 1902
rect 15292 1838 15344 1844
rect 15304 800 15332 1838
rect 15396 800 15424 4966
rect 15488 2774 15516 5510
rect 15580 5302 15608 6598
rect 15568 5296 15620 5302
rect 15568 5238 15620 5244
rect 15568 4276 15620 4282
rect 15568 4218 15620 4224
rect 15580 3097 15608 4218
rect 15566 3088 15622 3097
rect 15672 3058 15700 9318
rect 15752 6724 15804 6730
rect 15752 6666 15804 6672
rect 15764 6186 15792 6666
rect 15752 6180 15804 6186
rect 15752 6122 15804 6128
rect 15764 5914 15792 6122
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15856 4282 15884 14214
rect 15948 11286 15976 14282
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 16028 6248 16080 6254
rect 16028 6190 16080 6196
rect 16040 5710 16068 6190
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 16040 4690 16068 5646
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 15764 3398 15792 4082
rect 15842 4040 15898 4049
rect 15842 3975 15844 3984
rect 15896 3975 15898 3984
rect 15844 3946 15896 3952
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 15566 3023 15622 3032
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 15568 2984 15620 2990
rect 15620 2932 15700 2938
rect 15568 2926 15700 2932
rect 15580 2910 15700 2926
rect 15488 2746 15608 2774
rect 15580 1442 15608 2746
rect 15672 1578 15700 2910
rect 15672 1550 15884 1578
rect 15580 1414 15700 1442
rect 15568 1352 15620 1358
rect 15568 1294 15620 1300
rect 15580 800 15608 1294
rect 15672 800 15700 1414
rect 15856 800 15884 1550
rect 15948 800 15976 4558
rect 16040 3602 16068 4626
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 16132 3534 16160 5510
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 16028 3392 16080 3398
rect 16028 3334 16080 3340
rect 16040 1358 16068 3334
rect 16118 3224 16174 3233
rect 16118 3159 16120 3168
rect 16172 3159 16174 3168
rect 16120 3130 16172 3136
rect 16224 2582 16252 50322
rect 16396 41472 16448 41478
rect 16396 41414 16448 41420
rect 16408 40526 16436 41414
rect 16396 40520 16448 40526
rect 16396 40462 16448 40468
rect 16304 39636 16356 39642
rect 16304 39578 16356 39584
rect 16316 36378 16344 39578
rect 16304 36372 16356 36378
rect 16304 36314 16356 36320
rect 16500 35986 16528 55558
rect 17038 55519 17094 55528
rect 17682 55584 17738 55593
rect 17682 55519 17738 55528
rect 17788 55350 17816 55694
rect 17776 55344 17828 55350
rect 17774 55312 17776 55321
rect 17828 55312 17830 55321
rect 17774 55247 17830 55256
rect 16580 42560 16632 42566
rect 16580 42502 16632 42508
rect 16592 41614 16620 42502
rect 16672 42220 16724 42226
rect 16672 42162 16724 42168
rect 16948 42220 17000 42226
rect 16948 42162 17000 42168
rect 16580 41608 16632 41614
rect 16580 41550 16632 41556
rect 16592 41274 16620 41550
rect 16580 41268 16632 41274
rect 16580 41210 16632 41216
rect 16684 41206 16712 42162
rect 16672 41200 16724 41206
rect 16672 41142 16724 41148
rect 16960 40390 16988 42162
rect 17316 42016 17368 42022
rect 17316 41958 17368 41964
rect 17328 41614 17356 41958
rect 17132 41608 17184 41614
rect 17132 41550 17184 41556
rect 17316 41608 17368 41614
rect 17316 41550 17368 41556
rect 17144 41274 17172 41550
rect 17960 41540 18012 41546
rect 17960 41482 18012 41488
rect 17776 41472 17828 41478
rect 17776 41414 17828 41420
rect 17132 41268 17184 41274
rect 17132 41210 17184 41216
rect 17040 41132 17092 41138
rect 17040 41074 17092 41080
rect 16948 40384 17000 40390
rect 16948 40326 17000 40332
rect 17052 40186 17080 41074
rect 17684 40928 17736 40934
rect 17684 40870 17736 40876
rect 17500 40384 17552 40390
rect 17500 40326 17552 40332
rect 17040 40180 17092 40186
rect 17040 40122 17092 40128
rect 16856 39296 16908 39302
rect 16856 39238 16908 39244
rect 16868 38962 16896 39238
rect 16856 38956 16908 38962
rect 16856 38898 16908 38904
rect 16764 38344 16816 38350
rect 16764 38286 16816 38292
rect 16776 38049 16804 38286
rect 16762 38040 16818 38049
rect 16762 37975 16818 37984
rect 16764 37460 16816 37466
rect 16764 37402 16816 37408
rect 16776 36854 16804 37402
rect 16764 36848 16816 36854
rect 16764 36790 16816 36796
rect 16408 35958 16528 35986
rect 16304 34672 16356 34678
rect 16304 34614 16356 34620
rect 16316 34474 16344 34614
rect 16304 34468 16356 34474
rect 16304 34410 16356 34416
rect 16304 33584 16356 33590
rect 16304 33526 16356 33532
rect 16316 32910 16344 33526
rect 16304 32904 16356 32910
rect 16304 32846 16356 32852
rect 16408 22094 16436 35958
rect 16488 35692 16540 35698
rect 16488 35634 16540 35640
rect 16500 33522 16528 35634
rect 16764 34604 16816 34610
rect 16764 34546 16816 34552
rect 16488 33516 16540 33522
rect 16488 33458 16540 33464
rect 16500 32978 16528 33458
rect 16488 32972 16540 32978
rect 16488 32914 16540 32920
rect 16580 31272 16632 31278
rect 16580 31214 16632 31220
rect 16672 31272 16724 31278
rect 16672 31214 16724 31220
rect 16592 30258 16620 31214
rect 16580 30252 16632 30258
rect 16580 30194 16632 30200
rect 16684 30054 16712 31214
rect 16776 30938 16804 34546
rect 16868 31822 16896 38898
rect 17052 38350 17080 40122
rect 17512 38554 17540 40326
rect 17500 38548 17552 38554
rect 17500 38490 17552 38496
rect 17040 38344 17092 38350
rect 17040 38286 17092 38292
rect 17132 38344 17184 38350
rect 17132 38286 17184 38292
rect 17144 37874 17172 38286
rect 17316 38208 17368 38214
rect 17316 38150 17368 38156
rect 17328 37874 17356 38150
rect 17132 37868 17184 37874
rect 17132 37810 17184 37816
rect 17316 37868 17368 37874
rect 17316 37810 17368 37816
rect 17408 37868 17460 37874
rect 17408 37810 17460 37816
rect 17420 37466 17448 37810
rect 17408 37460 17460 37466
rect 17408 37402 17460 37408
rect 17040 37256 17092 37262
rect 17040 37198 17092 37204
rect 17592 37256 17644 37262
rect 17592 37198 17644 37204
rect 17052 36786 17080 37198
rect 17316 37188 17368 37194
rect 17316 37130 17368 37136
rect 17040 36780 17092 36786
rect 17040 36722 17092 36728
rect 17052 35698 17080 36722
rect 17328 36106 17356 37130
rect 17604 36582 17632 37198
rect 17592 36576 17644 36582
rect 17592 36518 17644 36524
rect 17316 36100 17368 36106
rect 17316 36042 17368 36048
rect 17040 35692 17092 35698
rect 17040 35634 17092 35640
rect 17132 35012 17184 35018
rect 17132 34954 17184 34960
rect 17144 34746 17172 34954
rect 17132 34740 17184 34746
rect 17132 34682 17184 34688
rect 17328 34678 17356 36042
rect 17604 34746 17632 36518
rect 17696 35086 17724 40870
rect 17788 40050 17816 41414
rect 17972 41138 18000 41482
rect 17960 41132 18012 41138
rect 17960 41074 18012 41080
rect 17776 40044 17828 40050
rect 17776 39986 17828 39992
rect 17868 37732 17920 37738
rect 17868 37674 17920 37680
rect 17880 37398 17908 37674
rect 17960 37664 18012 37670
rect 17960 37606 18012 37612
rect 17868 37392 17920 37398
rect 17868 37334 17920 37340
rect 17776 37256 17828 37262
rect 17776 37198 17828 37204
rect 17788 36922 17816 37198
rect 17866 37088 17922 37097
rect 17866 37023 17922 37032
rect 17776 36916 17828 36922
rect 17776 36858 17828 36864
rect 17880 36786 17908 37023
rect 17868 36780 17920 36786
rect 17868 36722 17920 36728
rect 17776 35488 17828 35494
rect 17776 35430 17828 35436
rect 17684 35080 17736 35086
rect 17684 35022 17736 35028
rect 17592 34740 17644 34746
rect 17592 34682 17644 34688
rect 17316 34672 17368 34678
rect 17316 34614 17368 34620
rect 17328 34134 17356 34614
rect 17684 34604 17736 34610
rect 17788 34592 17816 35430
rect 17736 34564 17816 34592
rect 17868 34604 17920 34610
rect 17684 34546 17736 34552
rect 17868 34546 17920 34552
rect 17500 34468 17552 34474
rect 17500 34410 17552 34416
rect 17316 34128 17368 34134
rect 17316 34070 17368 34076
rect 17512 33998 17540 34410
rect 17880 34066 17908 34546
rect 17868 34060 17920 34066
rect 17868 34002 17920 34008
rect 17040 33992 17092 33998
rect 17500 33992 17552 33998
rect 17040 33934 17092 33940
rect 17328 33952 17500 33980
rect 16948 33856 17000 33862
rect 16948 33798 17000 33804
rect 16960 33318 16988 33798
rect 17052 33454 17080 33934
rect 17040 33448 17092 33454
rect 17040 33390 17092 33396
rect 16948 33312 17000 33318
rect 16948 33254 17000 33260
rect 17224 33040 17276 33046
rect 17224 32982 17276 32988
rect 16948 32904 17000 32910
rect 16948 32846 17000 32852
rect 16856 31816 16908 31822
rect 16856 31758 16908 31764
rect 16868 31521 16896 31758
rect 16854 31512 16910 31521
rect 16854 31447 16856 31456
rect 16908 31447 16910 31456
rect 16856 31418 16908 31424
rect 16868 31387 16896 31418
rect 16960 31346 16988 32846
rect 17236 31958 17264 32982
rect 17224 31952 17276 31958
rect 17224 31894 17276 31900
rect 16948 31340 17000 31346
rect 16948 31282 17000 31288
rect 16764 30932 16816 30938
rect 16764 30874 16816 30880
rect 16776 30682 16804 30874
rect 16776 30654 16896 30682
rect 16764 30184 16816 30190
rect 16764 30126 16816 30132
rect 16672 30048 16724 30054
rect 16672 29990 16724 29996
rect 16776 29510 16804 30126
rect 16764 29504 16816 29510
rect 16764 29446 16816 29452
rect 16672 27464 16724 27470
rect 16672 27406 16724 27412
rect 16580 27396 16632 27402
rect 16580 27338 16632 27344
rect 16592 25906 16620 27338
rect 16684 26246 16712 27406
rect 16776 26382 16804 29446
rect 16868 28694 16896 30654
rect 17132 29776 17184 29782
rect 17132 29718 17184 29724
rect 17040 29504 17092 29510
rect 17040 29446 17092 29452
rect 16856 28688 16908 28694
rect 16856 28630 16908 28636
rect 16948 28416 17000 28422
rect 16948 28358 17000 28364
rect 16960 28082 16988 28358
rect 16948 28076 17000 28082
rect 16948 28018 17000 28024
rect 17052 26432 17080 29446
rect 16960 26404 17080 26432
rect 16764 26376 16816 26382
rect 16762 26344 16764 26353
rect 16816 26344 16818 26353
rect 16762 26279 16818 26288
rect 16672 26240 16724 26246
rect 16672 26182 16724 26188
rect 16580 25900 16632 25906
rect 16580 25842 16632 25848
rect 16684 25362 16712 26182
rect 16672 25356 16724 25362
rect 16672 25298 16724 25304
rect 16672 25220 16724 25226
rect 16672 25162 16724 25168
rect 16580 24404 16632 24410
rect 16580 24346 16632 24352
rect 16592 22234 16620 24346
rect 16684 24206 16712 25162
rect 16764 24812 16816 24818
rect 16764 24754 16816 24760
rect 16672 24200 16724 24206
rect 16670 24168 16672 24177
rect 16724 24168 16726 24177
rect 16776 24138 16804 24754
rect 16670 24103 16726 24112
rect 16764 24132 16816 24138
rect 16684 23254 16712 24103
rect 16764 24074 16816 24080
rect 16672 23248 16724 23254
rect 16672 23190 16724 23196
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16684 22574 16712 22918
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16580 22228 16632 22234
rect 16580 22170 16632 22176
rect 16408 22066 16528 22094
rect 16304 14816 16356 14822
rect 16304 14758 16356 14764
rect 16316 14278 16344 14758
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 16316 13938 16344 14214
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 16120 2100 16172 2106
rect 16120 2042 16172 2048
rect 16028 1352 16080 1358
rect 16028 1294 16080 1300
rect 16132 800 16160 2042
rect 16316 1170 16344 3878
rect 16408 3058 16436 8774
rect 16500 8430 16528 22066
rect 16592 17134 16620 22170
rect 16684 21486 16712 22510
rect 16672 21480 16724 21486
rect 16672 21422 16724 21428
rect 16684 19378 16712 21422
rect 16776 20262 16804 24074
rect 16960 21894 16988 26404
rect 17038 26344 17094 26353
rect 17038 26279 17094 26288
rect 16948 21888 17000 21894
rect 16948 21830 17000 21836
rect 16960 21706 16988 21830
rect 16868 21678 16988 21706
rect 16868 21146 16896 21678
rect 16948 21548 17000 21554
rect 16948 21490 17000 21496
rect 16960 21146 16988 21490
rect 16856 21140 16908 21146
rect 16856 21082 16908 21088
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 16868 20874 16896 21082
rect 16856 20868 16908 20874
rect 16856 20810 16908 20816
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16856 20256 16908 20262
rect 16856 20198 16908 20204
rect 16776 19514 16804 20198
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16764 19372 16816 19378
rect 16764 19314 16816 19320
rect 16776 18970 16804 19314
rect 16764 18964 16816 18970
rect 16764 18906 16816 18912
rect 16868 18850 16896 20198
rect 16776 18822 16896 18850
rect 16580 17128 16632 17134
rect 16580 17070 16632 17076
rect 16592 10470 16620 17070
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16592 9081 16620 10066
rect 16578 9072 16634 9081
rect 16578 9007 16634 9016
rect 16684 8786 16712 12242
rect 16776 10062 16804 18822
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16868 18426 16896 18702
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 16868 16590 16896 17274
rect 16856 16584 16908 16590
rect 16856 16526 16908 16532
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16868 15366 16896 16050
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16868 14074 16896 15302
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16960 12102 16988 18158
rect 17052 14226 17080 26279
rect 17144 24682 17172 29718
rect 17328 27878 17356 33952
rect 17500 33934 17552 33940
rect 17776 33992 17828 33998
rect 17776 33934 17828 33940
rect 17788 33658 17816 33934
rect 17868 33924 17920 33930
rect 17868 33866 17920 33872
rect 17776 33652 17828 33658
rect 17776 33594 17828 33600
rect 17684 32904 17736 32910
rect 17684 32846 17736 32852
rect 17776 32904 17828 32910
rect 17776 32846 17828 32852
rect 17592 32768 17644 32774
rect 17592 32710 17644 32716
rect 17408 30252 17460 30258
rect 17408 30194 17460 30200
rect 17420 29510 17448 30194
rect 17500 30048 17552 30054
rect 17500 29990 17552 29996
rect 17512 29646 17540 29990
rect 17500 29640 17552 29646
rect 17500 29582 17552 29588
rect 17408 29504 17460 29510
rect 17408 29446 17460 29452
rect 17316 27872 17368 27878
rect 17316 27814 17368 27820
rect 17500 26988 17552 26994
rect 17500 26930 17552 26936
rect 17222 26480 17278 26489
rect 17222 26415 17224 26424
rect 17276 26415 17278 26424
rect 17224 26386 17276 26392
rect 17236 25906 17264 26386
rect 17512 26042 17540 26930
rect 17500 26036 17552 26042
rect 17500 25978 17552 25984
rect 17224 25900 17276 25906
rect 17224 25842 17276 25848
rect 17316 25220 17368 25226
rect 17316 25162 17368 25168
rect 17132 24676 17184 24682
rect 17132 24618 17184 24624
rect 17224 24132 17276 24138
rect 17224 24074 17276 24080
rect 17236 22030 17264 24074
rect 17224 22024 17276 22030
rect 17224 21966 17276 21972
rect 17132 18692 17184 18698
rect 17132 18634 17184 18640
rect 17144 16590 17172 18634
rect 17132 16584 17184 16590
rect 17132 16526 17184 16532
rect 17132 16448 17184 16454
rect 17132 16390 17184 16396
rect 17144 14346 17172 16390
rect 17236 15162 17264 21966
rect 17328 18766 17356 25162
rect 17408 25152 17460 25158
rect 17408 25094 17460 25100
rect 17420 24818 17448 25094
rect 17408 24812 17460 24818
rect 17408 24754 17460 24760
rect 17420 23594 17448 24754
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17408 23588 17460 23594
rect 17408 23530 17460 23536
rect 17408 22432 17460 22438
rect 17408 22374 17460 22380
rect 17420 22166 17448 22374
rect 17408 22160 17460 22166
rect 17408 22102 17460 22108
rect 17512 21962 17540 24142
rect 17500 21956 17552 21962
rect 17500 21898 17552 21904
rect 17512 20806 17540 21898
rect 17500 20800 17552 20806
rect 17500 20742 17552 20748
rect 17512 20398 17540 20742
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17604 20262 17632 32710
rect 17696 32570 17724 32846
rect 17684 32564 17736 32570
rect 17684 32506 17736 32512
rect 17696 32366 17724 32506
rect 17788 32434 17816 32846
rect 17776 32428 17828 32434
rect 17776 32370 17828 32376
rect 17684 32360 17736 32366
rect 17684 32302 17736 32308
rect 17880 32230 17908 33866
rect 17972 33114 18000 37606
rect 18052 34536 18104 34542
rect 18052 34478 18104 34484
rect 17960 33108 18012 33114
rect 17960 33050 18012 33056
rect 17960 32564 18012 32570
rect 17960 32506 18012 32512
rect 17972 32473 18000 32506
rect 17958 32464 18014 32473
rect 17958 32399 17960 32408
rect 18012 32399 18014 32408
rect 17960 32370 18012 32376
rect 17960 32292 18012 32298
rect 18064 32280 18092 34478
rect 18012 32252 18092 32280
rect 17960 32234 18012 32240
rect 17868 32224 17920 32230
rect 17868 32166 17920 32172
rect 17880 31686 17908 32166
rect 17972 31890 18000 32234
rect 17960 31884 18012 31890
rect 17960 31826 18012 31832
rect 17868 31680 17920 31686
rect 17868 31622 17920 31628
rect 17880 31278 17908 31622
rect 17868 31272 17920 31278
rect 17868 31214 17920 31220
rect 17880 30734 17908 31214
rect 17868 30728 17920 30734
rect 17868 30670 17920 30676
rect 18052 30660 18104 30666
rect 18052 30602 18104 30608
rect 18064 30326 18092 30602
rect 18052 30320 18104 30326
rect 18052 30262 18104 30268
rect 17960 30116 18012 30122
rect 17960 30058 18012 30064
rect 17868 29640 17920 29646
rect 17868 29582 17920 29588
rect 17880 29238 17908 29582
rect 17972 29578 18000 30058
rect 17960 29572 18012 29578
rect 17960 29514 18012 29520
rect 17972 29238 18000 29514
rect 17868 29232 17920 29238
rect 17868 29174 17920 29180
rect 17960 29232 18012 29238
rect 17960 29174 18012 29180
rect 17880 28994 17908 29174
rect 17788 28966 17908 28994
rect 17684 27872 17736 27878
rect 17684 27814 17736 27820
rect 17696 27334 17724 27814
rect 17684 27328 17736 27334
rect 17684 27270 17736 27276
rect 17696 25906 17724 27270
rect 17684 25900 17736 25906
rect 17684 25842 17736 25848
rect 17788 25294 17816 28966
rect 17960 28416 18012 28422
rect 17960 28358 18012 28364
rect 17972 28218 18000 28358
rect 17960 28212 18012 28218
rect 17960 28154 18012 28160
rect 17972 27606 18000 28154
rect 17960 27600 18012 27606
rect 17960 27542 18012 27548
rect 17868 26444 17920 26450
rect 17868 26386 17920 26392
rect 17880 26042 17908 26386
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 17868 26036 17920 26042
rect 17868 25978 17920 25984
rect 17776 25288 17828 25294
rect 17776 25230 17828 25236
rect 17972 25158 18000 26318
rect 17960 25152 18012 25158
rect 17960 25094 18012 25100
rect 17684 24676 17736 24682
rect 17684 24618 17736 24624
rect 17696 24410 17724 24618
rect 17684 24404 17736 24410
rect 17684 24346 17736 24352
rect 18052 22976 18104 22982
rect 18052 22918 18104 22924
rect 17776 22432 17828 22438
rect 17696 22392 17776 22420
rect 17696 20618 17724 22392
rect 17776 22374 17828 22380
rect 17868 22160 17920 22166
rect 17788 22108 17868 22114
rect 17788 22102 17920 22108
rect 17788 22098 17908 22102
rect 17776 22092 17908 22098
rect 17828 22086 17908 22092
rect 17776 22034 17828 22040
rect 18064 22030 18092 22918
rect 17868 22024 17920 22030
rect 17868 21966 17920 21972
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 17880 21690 17908 21966
rect 17868 21684 17920 21690
rect 17868 21626 17920 21632
rect 17880 20942 17908 21626
rect 17868 20936 17920 20942
rect 17868 20878 17920 20884
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17696 20590 17816 20618
rect 17682 20496 17738 20505
rect 17682 20431 17684 20440
rect 17736 20431 17738 20440
rect 17684 20402 17736 20408
rect 17592 20256 17644 20262
rect 17592 20198 17644 20204
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 17316 16516 17368 16522
rect 17316 16458 17368 16464
rect 17328 16250 17356 16458
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17224 15156 17276 15162
rect 17224 15098 17276 15104
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 17328 14822 17356 14962
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17132 14340 17184 14346
rect 17132 14282 17184 14288
rect 17052 14198 17264 14226
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 17236 11286 17264 14198
rect 17604 13802 17632 19450
rect 17788 17354 17816 20590
rect 17972 19854 18000 20742
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 18052 19508 18104 19514
rect 18052 19450 18104 19456
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 17696 17326 17816 17354
rect 17592 13796 17644 13802
rect 17592 13738 17644 13744
rect 17696 12646 17724 17326
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17788 16250 17816 16526
rect 17776 16244 17828 16250
rect 17776 16186 17828 16192
rect 17972 16182 18000 18226
rect 18064 18222 18092 19450
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 18156 17218 18184 56782
rect 18524 55894 18552 57258
rect 18708 57050 18736 57394
rect 18972 57248 19024 57254
rect 18972 57190 19024 57196
rect 18696 57044 18748 57050
rect 18696 56986 18748 56992
rect 18788 56976 18840 56982
rect 18788 56918 18840 56924
rect 18800 56506 18828 56918
rect 18788 56500 18840 56506
rect 18788 56442 18840 56448
rect 18984 56370 19012 57190
rect 19536 57050 19564 57394
rect 19984 57384 20036 57390
rect 19984 57326 20036 57332
rect 19996 57050 20024 57326
rect 20168 57248 20220 57254
rect 20168 57190 20220 57196
rect 19524 57044 19576 57050
rect 19524 56986 19576 56992
rect 19984 57044 20036 57050
rect 19984 56986 20036 56992
rect 19340 56976 19392 56982
rect 19340 56918 19392 56924
rect 19064 56772 19116 56778
rect 19064 56714 19116 56720
rect 18880 56364 18932 56370
rect 18880 56306 18932 56312
rect 18972 56364 19024 56370
rect 18972 56306 19024 56312
rect 18512 55888 18564 55894
rect 18512 55830 18564 55836
rect 18788 55752 18840 55758
rect 18788 55694 18840 55700
rect 18800 55350 18828 55694
rect 18788 55344 18840 55350
rect 18786 55312 18788 55321
rect 18840 55312 18842 55321
rect 18786 55247 18842 55256
rect 18604 42016 18656 42022
rect 18604 41958 18656 41964
rect 18616 41750 18644 41958
rect 18604 41744 18656 41750
rect 18604 41686 18656 41692
rect 18616 41138 18644 41686
rect 18696 41676 18748 41682
rect 18696 41618 18748 41624
rect 18708 41414 18736 41618
rect 18708 41386 18828 41414
rect 18604 41132 18656 41138
rect 18604 41074 18656 41080
rect 18696 41064 18748 41070
rect 18696 41006 18748 41012
rect 18604 40996 18656 41002
rect 18604 40938 18656 40944
rect 18420 40928 18472 40934
rect 18420 40870 18472 40876
rect 18328 40520 18380 40526
rect 18328 40462 18380 40468
rect 18340 39982 18368 40462
rect 18432 40118 18460 40870
rect 18616 40730 18644 40938
rect 18604 40724 18656 40730
rect 18604 40666 18656 40672
rect 18616 40390 18644 40666
rect 18604 40384 18656 40390
rect 18604 40326 18656 40332
rect 18420 40112 18472 40118
rect 18420 40054 18472 40060
rect 18328 39976 18380 39982
rect 18328 39918 18380 39924
rect 18340 39098 18368 39918
rect 18328 39092 18380 39098
rect 18328 39034 18380 39040
rect 18340 37874 18368 39034
rect 18328 37868 18380 37874
rect 18328 37810 18380 37816
rect 18512 37868 18564 37874
rect 18512 37810 18564 37816
rect 18524 37466 18552 37810
rect 18512 37460 18564 37466
rect 18512 37402 18564 37408
rect 18708 36718 18736 41006
rect 18696 36712 18748 36718
rect 18696 36654 18748 36660
rect 18512 35692 18564 35698
rect 18512 35634 18564 35640
rect 18524 34950 18552 35634
rect 18604 35148 18656 35154
rect 18604 35090 18656 35096
rect 18512 34944 18564 34950
rect 18512 34886 18564 34892
rect 18524 34066 18552 34886
rect 18616 34474 18644 35090
rect 18696 34604 18748 34610
rect 18696 34546 18748 34552
rect 18604 34468 18656 34474
rect 18604 34410 18656 34416
rect 18616 34202 18644 34410
rect 18604 34196 18656 34202
rect 18604 34138 18656 34144
rect 18512 34060 18564 34066
rect 18512 34002 18564 34008
rect 18328 33380 18380 33386
rect 18328 33322 18380 33328
rect 18340 32434 18368 33322
rect 18708 32842 18736 34546
rect 18420 32836 18472 32842
rect 18420 32778 18472 32784
rect 18696 32836 18748 32842
rect 18696 32778 18748 32784
rect 18432 32570 18460 32778
rect 18420 32564 18472 32570
rect 18420 32506 18472 32512
rect 18328 32428 18380 32434
rect 18328 32370 18380 32376
rect 18708 31346 18736 32778
rect 18696 31340 18748 31346
rect 18696 31282 18748 31288
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 18524 29850 18552 30194
rect 18604 30184 18656 30190
rect 18604 30126 18656 30132
rect 18512 29844 18564 29850
rect 18512 29786 18564 29792
rect 18616 29578 18644 30126
rect 18604 29572 18656 29578
rect 18604 29514 18656 29520
rect 18236 28008 18288 28014
rect 18236 27950 18288 27956
rect 18248 24138 18276 27950
rect 18328 26376 18380 26382
rect 18328 26318 18380 26324
rect 18340 25974 18368 26318
rect 18328 25968 18380 25974
rect 18328 25910 18380 25916
rect 18340 24886 18368 25910
rect 18328 24880 18380 24886
rect 18328 24822 18380 24828
rect 18340 24274 18368 24822
rect 18512 24812 18564 24818
rect 18512 24754 18564 24760
rect 18328 24268 18380 24274
rect 18328 24210 18380 24216
rect 18236 24132 18288 24138
rect 18236 24074 18288 24080
rect 18524 23866 18552 24754
rect 18616 24698 18644 29514
rect 18696 27056 18748 27062
rect 18696 26998 18748 27004
rect 18708 26382 18736 26998
rect 18696 26376 18748 26382
rect 18696 26318 18748 26324
rect 18708 24818 18736 26318
rect 18696 24812 18748 24818
rect 18696 24754 18748 24760
rect 18616 24670 18736 24698
rect 18512 23860 18564 23866
rect 18512 23802 18564 23808
rect 18524 23769 18552 23802
rect 18510 23760 18566 23769
rect 18510 23695 18566 23704
rect 18604 23724 18656 23730
rect 18604 23666 18656 23672
rect 18616 23050 18644 23666
rect 18604 23044 18656 23050
rect 18604 22986 18656 22992
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18524 22166 18552 22578
rect 18512 22160 18564 22166
rect 18512 22102 18564 22108
rect 18616 21622 18644 22986
rect 18604 21616 18656 21622
rect 18604 21558 18656 21564
rect 18708 18850 18736 24670
rect 18616 18822 18736 18850
rect 18236 18760 18288 18766
rect 18236 18702 18288 18708
rect 18248 18426 18276 18702
rect 18236 18420 18288 18426
rect 18236 18362 18288 18368
rect 18064 17190 18184 17218
rect 17960 16176 18012 16182
rect 17960 16118 18012 16124
rect 17776 13796 17828 13802
rect 17776 13738 17828 13744
rect 17788 13530 17816 13738
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 17788 13190 17816 13466
rect 17868 13252 17920 13258
rect 17868 13194 17920 13200
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 17684 12640 17736 12646
rect 17684 12582 17736 12588
rect 17788 12434 17816 13126
rect 17880 12986 17908 13194
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17788 12406 17908 12434
rect 17224 11280 17276 11286
rect 17224 11222 17276 11228
rect 17776 11076 17828 11082
rect 17776 11018 17828 11024
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 17684 8900 17736 8906
rect 17684 8842 17736 8848
rect 16592 8758 16712 8786
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16592 6662 16620 8758
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17144 8498 17172 8570
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 16856 8356 16908 8362
rect 16856 8298 16908 8304
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 16592 6458 16620 6598
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 16592 6254 16620 6394
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16592 5370 16620 5646
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 16488 4752 16540 4758
rect 16488 4694 16540 4700
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16396 2916 16448 2922
rect 16396 2858 16448 2864
rect 16224 1142 16344 1170
rect 16224 800 16252 1142
rect 16408 800 16436 2858
rect 16500 800 16528 4694
rect 16684 4146 16712 7686
rect 16868 7478 16896 8298
rect 17144 8090 17172 8434
rect 17500 8424 17552 8430
rect 17500 8366 17552 8372
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17144 7954 17172 8026
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 16856 7472 16908 7478
rect 16856 7414 16908 7420
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 16856 6724 16908 6730
rect 16856 6666 16908 6672
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 16776 5234 16804 5646
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16764 4616 16816 4622
rect 16764 4558 16816 4564
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16672 2848 16724 2854
rect 16672 2790 16724 2796
rect 16684 800 16712 2790
rect 16776 800 16804 4558
rect 16868 2446 16896 6666
rect 16960 6322 16988 7346
rect 17052 7274 17080 7346
rect 17040 7268 17092 7274
rect 17040 7210 17092 7216
rect 17052 6798 17080 7210
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 16960 5710 16988 6258
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 17052 5302 17080 6734
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 17328 5681 17356 5714
rect 17314 5672 17370 5681
rect 17314 5607 17370 5616
rect 17040 5296 17092 5302
rect 17040 5238 17092 5244
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17040 3120 17092 3126
rect 17040 3062 17092 3068
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 16960 800 16988 2994
rect 17052 800 17080 3062
rect 17236 800 17264 4082
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17328 800 17356 3878
rect 17420 3534 17448 6598
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17406 3224 17462 3233
rect 17406 3159 17408 3168
rect 17460 3159 17462 3168
rect 17408 3130 17460 3136
rect 17512 2774 17540 8366
rect 17696 8090 17724 8842
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17788 5846 17816 11018
rect 17880 7886 17908 12406
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17880 7546 17908 7822
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17776 5840 17828 5846
rect 17776 5782 17828 5788
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17592 5568 17644 5574
rect 17592 5510 17644 5516
rect 17604 5234 17632 5510
rect 17880 5234 17908 5646
rect 17592 5228 17644 5234
rect 17868 5228 17920 5234
rect 17644 5188 17724 5216
rect 17592 5170 17644 5176
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17420 2746 17540 2774
rect 17420 2310 17448 2746
rect 17500 2576 17552 2582
rect 17498 2544 17500 2553
rect 17552 2544 17554 2553
rect 17498 2479 17554 2488
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 17512 800 17540 2382
rect 17604 800 17632 4966
rect 17696 3738 17724 5188
rect 17868 5170 17920 5176
rect 17868 4072 17920 4078
rect 17868 4014 17920 4020
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 17682 2680 17738 2689
rect 17682 2615 17738 2624
rect 17696 2582 17724 2615
rect 17684 2576 17736 2582
rect 17684 2518 17736 2524
rect 17788 800 17816 3130
rect 17880 800 17908 4014
rect 17972 2378 18000 8774
rect 18064 3126 18092 17190
rect 18144 17060 18196 17066
rect 18144 17002 18196 17008
rect 18156 16590 18184 17002
rect 18616 16658 18644 18822
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18604 16652 18656 16658
rect 18604 16594 18656 16600
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18236 16040 18288 16046
rect 18236 15982 18288 15988
rect 18248 14550 18276 15982
rect 18432 15026 18460 16390
rect 18708 15570 18736 18702
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18708 15094 18736 15506
rect 18696 15088 18748 15094
rect 18696 15030 18748 15036
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 18236 14544 18288 14550
rect 18236 14486 18288 14492
rect 18340 14414 18368 14962
rect 18328 14408 18380 14414
rect 18328 14350 18380 14356
rect 18340 12850 18368 14350
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 18156 11898 18184 12786
rect 18420 12708 18472 12714
rect 18420 12650 18472 12656
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 18156 11354 18184 11698
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18248 11014 18276 11834
rect 18432 11762 18460 12650
rect 18524 11762 18552 13126
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18512 11756 18564 11762
rect 18512 11698 18564 11704
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 18524 11082 18552 11290
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 18432 8786 18460 10406
rect 18604 9172 18656 9178
rect 18604 9114 18656 9120
rect 18156 8758 18460 8786
rect 18156 8566 18184 8758
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 18144 8356 18196 8362
rect 18144 8298 18196 8304
rect 18156 7886 18184 8298
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18248 7818 18276 8570
rect 18432 8498 18460 8758
rect 18616 8498 18644 9114
rect 18800 9058 18828 41386
rect 18892 31754 18920 56306
rect 18972 38752 19024 38758
rect 18972 38694 19024 38700
rect 18984 37330 19012 38694
rect 18972 37324 19024 37330
rect 18972 37266 19024 37272
rect 18984 36922 19012 37266
rect 18972 36916 19024 36922
rect 18972 36858 19024 36864
rect 18892 31726 19012 31754
rect 18878 26480 18934 26489
rect 18878 26415 18880 26424
rect 18932 26415 18934 26424
rect 18880 26386 18932 26392
rect 18880 25900 18932 25906
rect 18880 25842 18932 25848
rect 18892 25770 18920 25842
rect 18880 25764 18932 25770
rect 18880 25706 18932 25712
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 18892 21486 18920 21966
rect 18880 21480 18932 21486
rect 18880 21422 18932 21428
rect 18880 21344 18932 21350
rect 18880 21286 18932 21292
rect 18892 21010 18920 21286
rect 18880 21004 18932 21010
rect 18880 20946 18932 20952
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18892 12170 18920 12582
rect 18880 12164 18932 12170
rect 18880 12106 18932 12112
rect 18984 9178 19012 31726
rect 19076 12434 19104 56714
rect 19352 55894 19380 56918
rect 20180 56846 20208 57190
rect 20168 56840 20220 56846
rect 20166 56808 20168 56817
rect 20220 56808 20222 56817
rect 20166 56743 20222 56752
rect 20720 56704 20772 56710
rect 20720 56646 20772 56652
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 20732 56438 20760 56646
rect 22204 56506 22232 57394
rect 23388 56704 23440 56710
rect 23388 56646 23440 56652
rect 22192 56500 22244 56506
rect 22192 56442 22244 56448
rect 19432 56432 19484 56438
rect 19432 56374 19484 56380
rect 20720 56432 20772 56438
rect 20720 56374 20772 56380
rect 19340 55888 19392 55894
rect 19340 55830 19392 55836
rect 19444 45554 19472 56374
rect 19984 56364 20036 56370
rect 19984 56306 20036 56312
rect 20904 56364 20956 56370
rect 20904 56306 20956 56312
rect 21732 56364 21784 56370
rect 21732 56306 21784 56312
rect 22560 56364 22612 56370
rect 22560 56306 22612 56312
rect 23020 56364 23072 56370
rect 23020 56306 23072 56312
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 19996 55350 20024 56306
rect 20168 56296 20220 56302
rect 20168 56238 20220 56244
rect 20076 56160 20128 56166
rect 20076 56102 20128 56108
rect 20088 55962 20116 56102
rect 20076 55956 20128 55962
rect 20076 55898 20128 55904
rect 20076 55820 20128 55826
rect 20076 55762 20128 55768
rect 19800 55344 19852 55350
rect 19798 55312 19800 55321
rect 19984 55344 20036 55350
rect 19852 55312 19854 55321
rect 19984 55286 20036 55292
rect 19798 55247 19854 55256
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 20088 45554 20116 55762
rect 19352 45526 19472 45554
rect 19996 45526 20116 45554
rect 19248 38276 19300 38282
rect 19248 38218 19300 38224
rect 19260 38010 19288 38218
rect 19248 38004 19300 38010
rect 19248 37946 19300 37952
rect 19248 36712 19300 36718
rect 19248 36654 19300 36660
rect 19156 35284 19208 35290
rect 19156 35226 19208 35232
rect 19168 33590 19196 35226
rect 19260 34474 19288 36654
rect 19248 34468 19300 34474
rect 19248 34410 19300 34416
rect 19156 33584 19208 33590
rect 19156 33526 19208 33532
rect 19352 31754 19380 45526
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19996 41721 20024 45526
rect 19982 41712 20038 41721
rect 19982 41647 20038 41656
rect 19984 41608 20036 41614
rect 19984 41550 20036 41556
rect 19432 41472 19484 41478
rect 19432 41414 19484 41420
rect 19444 40390 19472 41414
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19524 40928 19576 40934
rect 19524 40870 19576 40876
rect 19536 40526 19564 40870
rect 19524 40520 19576 40526
rect 19524 40462 19576 40468
rect 19432 40384 19484 40390
rect 19432 40326 19484 40332
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19996 40186 20024 41550
rect 20076 41132 20128 41138
rect 20076 41074 20128 41080
rect 19984 40180 20036 40186
rect 19984 40122 20036 40128
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19432 38344 19484 38350
rect 19432 38286 19484 38292
rect 19444 37670 19472 38286
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19616 38004 19668 38010
rect 19616 37946 19668 37952
rect 19432 37664 19484 37670
rect 19432 37606 19484 37612
rect 19444 36854 19472 37606
rect 19628 37194 19656 37946
rect 19996 37942 20024 40122
rect 19984 37936 20036 37942
rect 19984 37878 20036 37884
rect 20088 37874 20116 41074
rect 20076 37868 20128 37874
rect 20076 37810 20128 37816
rect 19984 37664 20036 37670
rect 19984 37606 20036 37612
rect 19616 37188 19668 37194
rect 19616 37130 19668 37136
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19432 36848 19484 36854
rect 19432 36790 19484 36796
rect 19996 36786 20024 37606
rect 19800 36780 19852 36786
rect 19800 36722 19852 36728
rect 19984 36780 20036 36786
rect 19984 36722 20036 36728
rect 19812 36582 19840 36722
rect 19984 36644 20036 36650
rect 19984 36586 20036 36592
rect 19432 36576 19484 36582
rect 19432 36518 19484 36524
rect 19800 36576 19852 36582
rect 19800 36518 19852 36524
rect 19444 35290 19472 36518
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19432 35284 19484 35290
rect 19432 35226 19484 35232
rect 19444 34610 19472 35226
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19432 34604 19484 34610
rect 19432 34546 19484 34552
rect 19800 34400 19852 34406
rect 19996 34388 20024 36586
rect 20088 34746 20116 37810
rect 20076 34740 20128 34746
rect 20076 34682 20128 34688
rect 19852 34360 20024 34388
rect 19800 34342 19852 34348
rect 19812 33998 19840 34342
rect 19800 33992 19852 33998
rect 19800 33934 19852 33940
rect 19984 33856 20036 33862
rect 19984 33798 20036 33804
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19996 32842 20024 33798
rect 19984 32836 20036 32842
rect 19984 32778 20036 32784
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19352 31726 19472 31754
rect 19340 30592 19392 30598
rect 19340 30534 19392 30540
rect 19352 30410 19380 30534
rect 19260 30382 19380 30410
rect 19260 30326 19288 30382
rect 19248 30320 19300 30326
rect 19248 30262 19300 30268
rect 19340 30252 19392 30258
rect 19340 30194 19392 30200
rect 19352 29850 19380 30194
rect 19340 29844 19392 29850
rect 19340 29786 19392 29792
rect 19340 29572 19392 29578
rect 19340 29514 19392 29520
rect 19352 29034 19380 29514
rect 19340 29028 19392 29034
rect 19340 28970 19392 28976
rect 19340 28008 19392 28014
rect 19340 27950 19392 27956
rect 19248 26988 19300 26994
rect 19248 26930 19300 26936
rect 19260 26586 19288 26930
rect 19248 26580 19300 26586
rect 19248 26522 19300 26528
rect 19156 25900 19208 25906
rect 19156 25842 19208 25848
rect 19168 24138 19196 25842
rect 19352 25378 19380 27950
rect 19260 25362 19380 25378
rect 19248 25356 19380 25362
rect 19300 25350 19380 25356
rect 19248 25298 19300 25304
rect 19156 24132 19208 24138
rect 19156 24074 19208 24080
rect 19168 23594 19196 24074
rect 19156 23588 19208 23594
rect 19156 23530 19208 23536
rect 19260 22094 19288 25298
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19352 22778 19380 23054
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19168 22066 19288 22094
rect 19168 16810 19196 22066
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 19248 21412 19300 21418
rect 19248 21354 19300 21360
rect 19260 19961 19288 21354
rect 19246 19952 19302 19961
rect 19246 19887 19302 19896
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19260 18426 19288 19110
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19260 18154 19288 18226
rect 19248 18148 19300 18154
rect 19248 18090 19300 18096
rect 19352 16998 19380 21830
rect 19444 17524 19472 31726
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19984 31340 20036 31346
rect 19984 31282 20036 31288
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19996 30326 20024 31282
rect 20076 30864 20128 30870
rect 20076 30806 20128 30812
rect 19708 30320 19760 30326
rect 19708 30262 19760 30268
rect 19984 30320 20036 30326
rect 19984 30262 20036 30268
rect 19616 30184 19668 30190
rect 19616 30126 19668 30132
rect 19628 29714 19656 30126
rect 19720 30122 19748 30262
rect 19708 30116 19760 30122
rect 19708 30058 19760 30064
rect 19616 29708 19668 29714
rect 19616 29650 19668 29656
rect 20088 29646 20116 30806
rect 20180 30054 20208 56238
rect 20916 55622 20944 56306
rect 21744 55622 21772 56306
rect 22572 55826 22600 56306
rect 22560 55820 22612 55826
rect 22560 55762 22612 55768
rect 23032 55622 23060 56306
rect 23400 56166 23428 56646
rect 24412 56506 24440 57394
rect 24676 57316 24728 57322
rect 24676 57258 24728 57264
rect 24688 56506 24716 57258
rect 24400 56500 24452 56506
rect 24400 56442 24452 56448
rect 24676 56500 24728 56506
rect 24676 56442 24728 56448
rect 23756 56364 23808 56370
rect 23756 56306 23808 56312
rect 24400 56364 24452 56370
rect 24400 56306 24452 56312
rect 25136 56364 25188 56370
rect 25136 56306 25188 56312
rect 23388 56160 23440 56166
rect 23388 56102 23440 56108
rect 23768 55622 23796 56306
rect 24412 55622 24440 56306
rect 25148 55622 25176 56306
rect 25332 56166 25360 57394
rect 26344 56506 26372 57462
rect 26976 57452 27028 57458
rect 26976 57394 27028 57400
rect 28448 57452 28500 57458
rect 28448 57394 28500 57400
rect 30104 57452 30156 57458
rect 30104 57394 30156 57400
rect 26988 56506 27016 57394
rect 28460 56506 28488 57394
rect 30116 56506 30144 57394
rect 26332 56500 26384 56506
rect 26332 56442 26384 56448
rect 26976 56500 27028 56506
rect 26976 56442 27028 56448
rect 28448 56500 28500 56506
rect 28448 56442 28500 56448
rect 30104 56500 30156 56506
rect 30104 56442 30156 56448
rect 26056 56364 26108 56370
rect 26056 56306 26108 56312
rect 26792 56364 26844 56370
rect 26792 56306 26844 56312
rect 27988 56364 28040 56370
rect 27988 56306 28040 56312
rect 29184 56364 29236 56370
rect 29184 56306 29236 56312
rect 29920 56364 29972 56370
rect 29920 56306 29972 56312
rect 25320 56160 25372 56166
rect 25320 56102 25372 56108
rect 26068 55622 26096 56306
rect 26804 55622 26832 56306
rect 28000 56166 28028 56306
rect 27988 56160 28040 56166
rect 27988 56102 28040 56108
rect 20260 55616 20312 55622
rect 20258 55584 20260 55593
rect 20904 55616 20956 55622
rect 20312 55584 20314 55593
rect 21732 55616 21784 55622
rect 20904 55558 20956 55564
rect 21730 55584 21732 55593
rect 23020 55616 23072 55622
rect 21784 55584 21786 55593
rect 20258 55519 20314 55528
rect 20916 50386 20944 55558
rect 21730 55519 21786 55528
rect 23018 55584 23020 55593
rect 23756 55616 23808 55622
rect 23072 55584 23074 55593
rect 23018 55519 23074 55528
rect 23754 55584 23756 55593
rect 24400 55616 24452 55622
rect 23808 55584 23810 55593
rect 24400 55558 24452 55564
rect 25136 55616 25188 55622
rect 25136 55558 25188 55564
rect 26056 55616 26108 55622
rect 26056 55558 26108 55564
rect 26792 55616 26844 55622
rect 26792 55558 26844 55564
rect 23754 55519 23810 55528
rect 20904 50380 20956 50386
rect 20904 50322 20956 50328
rect 24412 44878 24440 55558
rect 24400 44872 24452 44878
rect 24400 44814 24452 44820
rect 24308 41744 24360 41750
rect 24308 41686 24360 41692
rect 20260 41540 20312 41546
rect 20260 41482 20312 41488
rect 20272 41138 20300 41482
rect 24124 41268 24176 41274
rect 24124 41210 24176 41216
rect 20628 41200 20680 41206
rect 20628 41142 20680 41148
rect 20260 41132 20312 41138
rect 20260 41074 20312 41080
rect 20640 40390 20668 41142
rect 23756 40996 23808 41002
rect 23756 40938 23808 40944
rect 22100 40928 22152 40934
rect 22100 40870 22152 40876
rect 23020 40928 23072 40934
rect 23020 40870 23072 40876
rect 22112 40526 22140 40870
rect 22100 40520 22152 40526
rect 22100 40462 22152 40468
rect 22284 40520 22336 40526
rect 22284 40462 22336 40468
rect 22468 40520 22520 40526
rect 22468 40462 22520 40468
rect 20352 40384 20404 40390
rect 20352 40326 20404 40332
rect 20628 40384 20680 40390
rect 20628 40326 20680 40332
rect 22100 40384 22152 40390
rect 22100 40326 22152 40332
rect 20260 38344 20312 38350
rect 20260 38286 20312 38292
rect 20272 37738 20300 38286
rect 20260 37732 20312 37738
rect 20260 37674 20312 37680
rect 20272 37262 20300 37674
rect 20260 37256 20312 37262
rect 20260 37198 20312 37204
rect 20272 36650 20300 37198
rect 20260 36644 20312 36650
rect 20260 36586 20312 36592
rect 20364 36582 20392 40326
rect 20640 38282 20668 40326
rect 21456 40112 21508 40118
rect 21456 40054 21508 40060
rect 20996 40044 21048 40050
rect 20996 39986 21048 39992
rect 21008 39302 21036 39986
rect 20996 39296 21048 39302
rect 20996 39238 21048 39244
rect 20628 38276 20680 38282
rect 20628 38218 20680 38224
rect 20444 37868 20496 37874
rect 20444 37810 20496 37816
rect 20456 37466 20484 37810
rect 20444 37460 20496 37466
rect 20444 37402 20496 37408
rect 20444 37188 20496 37194
rect 20444 37130 20496 37136
rect 20536 37188 20588 37194
rect 20536 37130 20588 37136
rect 20352 36576 20404 36582
rect 20352 36518 20404 36524
rect 20352 35012 20404 35018
rect 20352 34954 20404 34960
rect 20260 34944 20312 34950
rect 20260 34886 20312 34892
rect 20272 34610 20300 34886
rect 20364 34746 20392 34954
rect 20352 34740 20404 34746
rect 20352 34682 20404 34688
rect 20260 34604 20312 34610
rect 20260 34546 20312 34552
rect 20272 33930 20300 34546
rect 20456 34066 20484 37130
rect 20548 36922 20576 37130
rect 20628 37120 20680 37126
rect 20628 37062 20680 37068
rect 20536 36916 20588 36922
rect 20536 36858 20588 36864
rect 20536 35080 20588 35086
rect 20536 35022 20588 35028
rect 20548 34678 20576 35022
rect 20536 34672 20588 34678
rect 20536 34614 20588 34620
rect 20640 34610 20668 37062
rect 21008 36242 21036 39238
rect 21468 39030 21496 40054
rect 22112 39370 22140 40326
rect 22296 40050 22324 40462
rect 22480 40050 22508 40462
rect 22744 40452 22796 40458
rect 22744 40394 22796 40400
rect 22756 40050 22784 40394
rect 23032 40050 23060 40870
rect 23388 40520 23440 40526
rect 23388 40462 23440 40468
rect 23112 40452 23164 40458
rect 23112 40394 23164 40400
rect 22284 40044 22336 40050
rect 22284 39986 22336 39992
rect 22468 40044 22520 40050
rect 22468 39986 22520 39992
rect 22652 40044 22704 40050
rect 22652 39986 22704 39992
rect 22744 40044 22796 40050
rect 22744 39986 22796 39992
rect 23020 40044 23072 40050
rect 23020 39986 23072 39992
rect 22480 39522 22508 39986
rect 22480 39494 22600 39522
rect 22572 39438 22600 39494
rect 22560 39432 22612 39438
rect 22560 39374 22612 39380
rect 22008 39364 22060 39370
rect 22008 39306 22060 39312
rect 22100 39364 22152 39370
rect 22100 39306 22152 39312
rect 22468 39364 22520 39370
rect 22468 39306 22520 39312
rect 21456 39024 21508 39030
rect 21456 38966 21508 38972
rect 21088 38208 21140 38214
rect 21088 38150 21140 38156
rect 20996 36236 21048 36242
rect 20996 36178 21048 36184
rect 20628 34604 20680 34610
rect 20628 34546 20680 34552
rect 20444 34060 20496 34066
rect 20444 34002 20496 34008
rect 20260 33924 20312 33930
rect 20260 33866 20312 33872
rect 20352 33108 20404 33114
rect 20352 33050 20404 33056
rect 20260 30592 20312 30598
rect 20260 30534 20312 30540
rect 20272 30190 20300 30534
rect 20260 30184 20312 30190
rect 20260 30126 20312 30132
rect 20168 30048 20220 30054
rect 20168 29990 20220 29996
rect 20166 29880 20222 29889
rect 20166 29815 20222 29824
rect 20076 29640 20128 29646
rect 19996 29600 20076 29628
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19892 29300 19944 29306
rect 19892 29242 19944 29248
rect 19904 29209 19932 29242
rect 19890 29200 19946 29209
rect 19996 29170 20024 29600
rect 20076 29582 20128 29588
rect 20074 29472 20130 29481
rect 20074 29407 20130 29416
rect 20088 29238 20116 29407
rect 20180 29288 20208 29815
rect 20272 29578 20300 30126
rect 20260 29572 20312 29578
rect 20260 29514 20312 29520
rect 20260 29300 20312 29306
rect 20180 29260 20260 29288
rect 20260 29242 20312 29248
rect 20076 29232 20128 29238
rect 20076 29174 20128 29180
rect 19890 29135 19946 29144
rect 19984 29164 20036 29170
rect 19984 29106 20036 29112
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 20088 28082 20116 29174
rect 20166 29064 20222 29073
rect 20166 28999 20222 29008
rect 20260 29028 20312 29034
rect 20076 28076 20128 28082
rect 20076 28018 20128 28024
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 20076 26784 20128 26790
rect 20076 26726 20128 26732
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19984 25900 20036 25906
rect 20088 25888 20116 26726
rect 20036 25860 20116 25888
rect 19984 25842 20036 25848
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19984 20936 20036 20942
rect 19984 20878 20036 20884
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19800 20528 19852 20534
rect 19996 20482 20024 20878
rect 19800 20470 19852 20476
rect 19524 20460 19576 20466
rect 19524 20402 19576 20408
rect 19536 20058 19564 20402
rect 19524 20052 19576 20058
rect 19524 19994 19576 20000
rect 19812 19802 19840 20470
rect 19904 20466 20024 20482
rect 19892 20460 20024 20466
rect 19944 20454 20024 20460
rect 19892 20402 19944 20408
rect 19904 19922 19932 20402
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19892 19916 19944 19922
rect 19892 19858 19944 19864
rect 19812 19786 19932 19802
rect 19812 19780 19944 19786
rect 19812 19774 19892 19780
rect 19892 19722 19944 19728
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 17678 20024 20198
rect 20088 19854 20116 25860
rect 20180 24342 20208 28999
rect 20260 28970 20312 28976
rect 20272 28014 20300 28970
rect 20260 28008 20312 28014
rect 20260 27950 20312 27956
rect 20168 24336 20220 24342
rect 20168 24278 20220 24284
rect 20364 22234 20392 33050
rect 20536 32496 20588 32502
rect 20536 32438 20588 32444
rect 20444 31816 20496 31822
rect 20444 31758 20496 31764
rect 20456 30326 20484 31758
rect 20444 30320 20496 30326
rect 20444 30262 20496 30268
rect 20444 30048 20496 30054
rect 20444 29990 20496 29996
rect 20456 23322 20484 29990
rect 20548 29209 20576 32438
rect 20996 31340 21048 31346
rect 20996 31282 21048 31288
rect 20720 31136 20772 31142
rect 20720 31078 20772 31084
rect 20628 30116 20680 30122
rect 20628 30058 20680 30064
rect 20640 29578 20668 30058
rect 20732 29714 20760 31078
rect 21008 30258 21036 31282
rect 20996 30252 21048 30258
rect 20996 30194 21048 30200
rect 20812 30048 20864 30054
rect 20812 29990 20864 29996
rect 20720 29708 20772 29714
rect 20720 29650 20772 29656
rect 20628 29572 20680 29578
rect 20628 29514 20680 29520
rect 20534 29200 20590 29209
rect 20534 29135 20590 29144
rect 20536 29028 20588 29034
rect 20536 28970 20588 28976
rect 20626 29008 20682 29017
rect 20444 23316 20496 23322
rect 20444 23258 20496 23264
rect 20444 22772 20496 22778
rect 20444 22714 20496 22720
rect 20352 22228 20404 22234
rect 20352 22170 20404 22176
rect 20260 21956 20312 21962
rect 20260 21898 20312 21904
rect 20272 21418 20300 21898
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20260 21412 20312 21418
rect 20260 21354 20312 21360
rect 20260 20868 20312 20874
rect 20260 20810 20312 20816
rect 20168 20800 20220 20806
rect 20168 20742 20220 20748
rect 20180 20602 20208 20742
rect 20168 20596 20220 20602
rect 20168 20538 20220 20544
rect 20168 20460 20220 20466
rect 20168 20402 20220 20408
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 19444 17496 20024 17524
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19168 16782 19380 16810
rect 19352 15706 19380 16782
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19444 16232 19472 16390
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19444 16204 19564 16232
rect 19432 16108 19484 16114
rect 19432 16050 19484 16056
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19352 14278 19380 15438
rect 19444 15162 19472 16050
rect 19536 15570 19564 16204
rect 19892 15972 19944 15978
rect 19892 15914 19944 15920
rect 19904 15706 19932 15914
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19524 15564 19576 15570
rect 19524 15506 19576 15512
rect 19536 15366 19564 15506
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19890 15056 19946 15065
rect 19890 14991 19946 15000
rect 19904 14958 19932 14991
rect 19892 14952 19944 14958
rect 19892 14894 19944 14900
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19444 14414 19472 14758
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19352 14006 19380 14214
rect 19444 14006 19472 14350
rect 19904 14346 19932 14894
rect 19892 14340 19944 14346
rect 19892 14282 19944 14288
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19156 12844 19208 12850
rect 19208 12804 19288 12832
rect 19156 12786 19208 12792
rect 19076 12406 19196 12434
rect 19064 11756 19116 11762
rect 19064 11698 19116 11704
rect 19076 10470 19104 11698
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 18972 9172 19024 9178
rect 18972 9114 19024 9120
rect 18800 9030 18920 9058
rect 18788 8900 18840 8906
rect 18788 8842 18840 8848
rect 18800 8634 18828 8842
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18236 7812 18288 7818
rect 18236 7754 18288 7760
rect 18696 7812 18748 7818
rect 18696 7754 18748 7760
rect 18144 7200 18196 7206
rect 18144 7142 18196 7148
rect 18156 6254 18184 7142
rect 18708 6866 18736 7754
rect 18788 7268 18840 7274
rect 18788 7210 18840 7216
rect 18696 6860 18748 6866
rect 18696 6802 18748 6808
rect 18512 6724 18564 6730
rect 18512 6666 18564 6672
rect 18696 6724 18748 6730
rect 18696 6666 18748 6672
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 18156 5710 18184 6054
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 18524 5642 18552 6666
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 18616 5914 18644 6258
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18512 5636 18564 5642
rect 18512 5578 18564 5584
rect 18524 5234 18552 5578
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 18144 4548 18196 4554
rect 18144 4490 18196 4496
rect 18052 3120 18104 3126
rect 18052 3062 18104 3068
rect 17960 2372 18012 2378
rect 17960 2314 18012 2320
rect 17972 1714 18000 2314
rect 17972 1686 18092 1714
rect 18064 800 18092 1686
rect 18156 800 18184 4490
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18340 800 18368 3470
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 18432 800 18460 2790
rect 18524 1170 18552 2994
rect 18616 2666 18644 4558
rect 18708 3058 18736 6666
rect 18800 6390 18828 7210
rect 18788 6384 18840 6390
rect 18788 6326 18840 6332
rect 18788 6248 18840 6254
rect 18788 6190 18840 6196
rect 18800 5234 18828 6190
rect 18788 5228 18840 5234
rect 18788 5170 18840 5176
rect 18892 5114 18920 9030
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 19076 7206 19104 7822
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 18800 5086 18920 5114
rect 18800 3942 18828 5086
rect 18880 5024 18932 5030
rect 18880 4966 18932 4972
rect 18892 4622 18920 4966
rect 18972 4752 19024 4758
rect 18972 4694 19024 4700
rect 18880 4616 18932 4622
rect 18880 4558 18932 4564
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18880 3392 18932 3398
rect 18786 3360 18842 3369
rect 18880 3334 18932 3340
rect 18786 3295 18842 3304
rect 18800 3126 18828 3295
rect 18788 3120 18840 3126
rect 18788 3062 18840 3068
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 18786 2680 18842 2689
rect 18616 2638 18736 2666
rect 18524 1142 18644 1170
rect 18616 800 18644 1142
rect 18708 800 18736 2638
rect 18786 2615 18842 2624
rect 18800 2582 18828 2615
rect 18788 2576 18840 2582
rect 18788 2518 18840 2524
rect 18892 2106 18920 3334
rect 18880 2100 18932 2106
rect 18880 2042 18932 2048
rect 18880 1760 18932 1766
rect 18880 1702 18932 1708
rect 18892 800 18920 1702
rect 18984 800 19012 4694
rect 19076 3126 19104 6598
rect 19168 3670 19196 12406
rect 19260 11014 19288 12804
rect 19444 12714 19472 13262
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19340 12708 19392 12714
rect 19340 12650 19392 12656
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 19352 12442 19380 12650
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19444 12306 19472 12650
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19340 11076 19392 11082
rect 19340 11018 19392 11024
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 19352 10470 19380 11018
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19616 10464 19668 10470
rect 19616 10406 19668 10412
rect 19628 10198 19656 10406
rect 19616 10192 19668 10198
rect 19616 10134 19668 10140
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19260 8974 19288 9454
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19260 5778 19288 8910
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19432 8492 19484 8498
rect 19352 8452 19432 8480
rect 19352 7410 19380 8452
rect 19432 8434 19484 8440
rect 19430 8392 19486 8401
rect 19430 8327 19486 8336
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 19352 5302 19380 6054
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 19156 3664 19208 3670
rect 19156 3606 19208 3612
rect 19248 3664 19300 3670
rect 19248 3606 19300 3612
rect 19064 3120 19116 3126
rect 19116 3080 19196 3108
rect 19064 3062 19116 3068
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 19076 2446 19104 2926
rect 19064 2440 19116 2446
rect 19064 2382 19116 2388
rect 19076 1766 19104 2382
rect 19064 1760 19116 1766
rect 19064 1702 19116 1708
rect 19168 800 19196 3080
rect 19260 2990 19288 3606
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 19352 2774 19380 4966
rect 19444 4128 19472 8327
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19996 6746 20024 17496
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 20088 14278 20116 14350
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 20180 13274 20208 20402
rect 20272 17678 20300 20810
rect 20364 20466 20392 21490
rect 20456 20942 20484 22714
rect 20444 20936 20496 20942
rect 20444 20878 20496 20884
rect 20548 20466 20576 28970
rect 20626 28943 20682 28952
rect 20640 26874 20668 28943
rect 20720 28484 20772 28490
rect 20720 28426 20772 28432
rect 20732 27470 20760 28426
rect 20720 27464 20772 27470
rect 20720 27406 20772 27412
rect 20824 27130 20852 29990
rect 20904 29572 20956 29578
rect 20904 29514 20956 29520
rect 20916 28966 20944 29514
rect 20904 28960 20956 28966
rect 20904 28902 20956 28908
rect 20996 27396 21048 27402
rect 20996 27338 21048 27344
rect 20812 27124 20864 27130
rect 20812 27066 20864 27072
rect 20640 26846 20760 26874
rect 20628 26784 20680 26790
rect 20628 26726 20680 26732
rect 20640 25974 20668 26726
rect 20628 25968 20680 25974
rect 20628 25910 20680 25916
rect 20640 24585 20668 25910
rect 20626 24576 20682 24585
rect 20626 24511 20682 24520
rect 20732 24154 20760 26846
rect 20812 26580 20864 26586
rect 20812 26522 20864 26528
rect 20824 26382 20852 26522
rect 20904 26444 20956 26450
rect 20904 26386 20956 26392
rect 20812 26376 20864 26382
rect 20812 26318 20864 26324
rect 20916 26246 20944 26386
rect 20904 26240 20956 26246
rect 20904 26182 20956 26188
rect 21008 25974 21036 27338
rect 20996 25968 21048 25974
rect 20996 25910 21048 25916
rect 20996 25696 21048 25702
rect 20996 25638 21048 25644
rect 21008 24614 21036 25638
rect 20904 24608 20956 24614
rect 20904 24550 20956 24556
rect 20996 24608 21048 24614
rect 20996 24550 21048 24556
rect 20916 24206 20944 24550
rect 20640 24126 20760 24154
rect 20904 24200 20956 24206
rect 20904 24142 20956 24148
rect 20996 24132 21048 24138
rect 20640 20942 20668 24126
rect 20996 24074 21048 24080
rect 21008 23662 21036 24074
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 20996 23316 21048 23322
rect 20996 23258 21048 23264
rect 20628 20936 20680 20942
rect 20628 20878 20680 20884
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20260 17672 20312 17678
rect 20260 17614 20312 17620
rect 20444 17536 20496 17542
rect 20444 17478 20496 17484
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 20272 15570 20300 16594
rect 20352 15904 20404 15910
rect 20352 15846 20404 15852
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20272 14822 20300 15506
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 20364 14618 20392 15846
rect 20352 14612 20404 14618
rect 20352 14554 20404 14560
rect 20180 13246 20300 13274
rect 20272 12918 20300 13246
rect 20260 12912 20312 12918
rect 20260 12854 20312 12860
rect 20168 12164 20220 12170
rect 20168 12106 20220 12112
rect 20180 11830 20208 12106
rect 20272 11898 20300 12854
rect 20260 11892 20312 11898
rect 20260 11834 20312 11840
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 20076 11008 20128 11014
rect 20076 10950 20128 10956
rect 20088 8090 20116 10950
rect 20456 10130 20484 17478
rect 20548 15008 20576 19858
rect 20628 19236 20680 19242
rect 20628 19178 20680 19184
rect 20640 18970 20668 19178
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20640 18222 20668 18906
rect 20904 18828 20956 18834
rect 20904 18770 20956 18776
rect 20812 18692 20864 18698
rect 20812 18634 20864 18640
rect 20628 18216 20680 18222
rect 20628 18158 20680 18164
rect 20720 16720 20772 16726
rect 20720 16662 20772 16668
rect 20732 16096 20760 16662
rect 20824 16250 20852 18634
rect 20916 17542 20944 18770
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20812 16108 20864 16114
rect 20732 16068 20812 16096
rect 20812 16050 20864 16056
rect 20824 15502 20852 16050
rect 20812 15496 20864 15502
rect 20810 15464 20812 15473
rect 20864 15464 20866 15473
rect 20810 15399 20866 15408
rect 20824 15373 20852 15399
rect 20916 15162 20944 17478
rect 20904 15156 20956 15162
rect 20904 15098 20956 15104
rect 20628 15020 20680 15026
rect 20548 14980 20628 15008
rect 20628 14962 20680 14968
rect 20640 14482 20668 14962
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20548 14006 20576 14418
rect 20628 14272 20680 14278
rect 20628 14214 20680 14220
rect 20536 14000 20588 14006
rect 20536 13942 20588 13948
rect 20534 13560 20590 13569
rect 20534 13495 20536 13504
rect 20588 13495 20590 13504
rect 20536 13466 20588 13472
rect 20548 12782 20576 13466
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 20548 11762 20576 12718
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20444 10124 20496 10130
rect 20444 10066 20496 10072
rect 20640 9654 20668 14214
rect 20916 12850 20944 15098
rect 20904 12844 20956 12850
rect 20904 12786 20956 12792
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20824 12306 20852 12582
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 20720 9988 20772 9994
rect 20720 9930 20772 9936
rect 20628 9648 20680 9654
rect 20628 9590 20680 9596
rect 20168 9580 20220 9586
rect 20168 9522 20220 9528
rect 20180 8838 20208 9522
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 20180 8566 20208 8774
rect 20168 8560 20220 8566
rect 20168 8502 20220 8508
rect 20076 8084 20128 8090
rect 20076 8026 20128 8032
rect 20088 7274 20116 8026
rect 20076 7268 20128 7274
rect 20076 7210 20128 7216
rect 19996 6718 20116 6746
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19444 4100 19564 4128
rect 19432 4004 19484 4010
rect 19432 3946 19484 3952
rect 19444 3040 19472 3946
rect 19536 3380 19564 4100
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 19720 3398 19748 3878
rect 19505 3352 19564 3380
rect 19708 3392 19760 3398
rect 19505 3176 19533 3352
rect 19708 3334 19760 3340
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19505 3148 19656 3176
rect 19444 3012 19564 3040
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 19260 2746 19380 2774
rect 19260 800 19288 2746
rect 19444 2446 19472 2858
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19444 1222 19472 2382
rect 19536 2360 19564 3012
rect 19628 2990 19656 3148
rect 19890 3088 19946 3097
rect 19996 3058 20024 6598
rect 20088 5302 20116 6718
rect 20444 6656 20496 6662
rect 20444 6598 20496 6604
rect 20168 6112 20220 6118
rect 20168 6054 20220 6060
rect 20076 5296 20128 5302
rect 20076 5238 20128 5244
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 19890 3023 19946 3032
rect 19984 3052 20036 3058
rect 19616 2984 19668 2990
rect 19616 2926 19668 2932
rect 19904 2922 19932 3023
rect 19984 2994 20036 3000
rect 19892 2916 19944 2922
rect 19892 2858 19944 2864
rect 19800 2848 19852 2854
rect 19798 2816 19800 2825
rect 19852 2816 19854 2825
rect 19798 2751 19854 2760
rect 19505 2332 19564 2360
rect 19505 2088 19533 2332
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19616 2100 19668 2106
rect 19505 2060 19564 2088
rect 19536 1358 19564 2060
rect 19616 2042 19668 2048
rect 19524 1352 19576 1358
rect 19524 1294 19576 1300
rect 19432 1216 19484 1222
rect 19628 1170 19656 2042
rect 19996 1442 20024 2994
rect 19432 1158 19484 1164
rect 19536 1142 19656 1170
rect 19720 1414 20024 1442
rect 19432 944 19484 950
rect 19432 886 19484 892
rect 19444 800 19472 886
rect 19536 800 19564 1142
rect 19720 800 19748 1414
rect 19800 1352 19852 1358
rect 19800 1294 19852 1300
rect 19984 1352 20036 1358
rect 19984 1294 20036 1300
rect 19812 800 19840 1294
rect 19996 800 20024 1294
rect 20088 800 20116 4966
rect 20180 3534 20208 6054
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 20258 3768 20314 3777
rect 20258 3703 20260 3712
rect 20312 3703 20314 3712
rect 20260 3674 20312 3680
rect 20168 3528 20220 3534
rect 20220 3488 20300 3516
rect 20168 3470 20220 3476
rect 20168 3392 20220 3398
rect 20168 3334 20220 3340
rect 20180 1086 20208 3334
rect 20272 1562 20300 3488
rect 20364 2990 20392 3878
rect 20456 3097 20484 6598
rect 20442 3088 20498 3097
rect 20442 3023 20498 3032
rect 20352 2984 20404 2990
rect 20548 2938 20576 9114
rect 20640 8974 20668 9590
rect 20732 9178 20760 9930
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20732 8634 20760 9114
rect 20720 8628 20772 8634
rect 20720 8570 20772 8576
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20732 6390 20760 7890
rect 20824 7886 20852 11018
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 20732 6202 20760 6326
rect 20732 6174 20852 6202
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20640 3126 20668 6054
rect 20628 3120 20680 3126
rect 20628 3062 20680 3068
rect 20352 2926 20404 2932
rect 20456 2910 20576 2938
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 20456 2774 20484 2910
rect 20536 2848 20588 2854
rect 20536 2790 20588 2796
rect 20364 2746 20484 2774
rect 20364 2650 20392 2746
rect 20352 2644 20404 2650
rect 20352 2586 20404 2592
rect 20352 2372 20404 2378
rect 20352 2314 20404 2320
rect 20260 1556 20312 1562
rect 20260 1498 20312 1504
rect 20364 1442 20392 2314
rect 20272 1414 20392 1442
rect 20168 1080 20220 1086
rect 20168 1022 20220 1028
rect 20272 800 20300 1414
rect 20352 1080 20404 1086
rect 20352 1022 20404 1028
rect 20364 800 20392 1022
rect 20548 800 20576 2790
rect 20640 800 20668 2926
rect 20732 2378 20760 6054
rect 20824 4826 20852 6174
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20812 4820 20864 4826
rect 20812 4762 20864 4768
rect 20812 3460 20864 3466
rect 20812 3402 20864 3408
rect 20720 2372 20772 2378
rect 20720 2314 20772 2320
rect 20732 1766 20760 2314
rect 20720 1760 20772 1766
rect 20720 1702 20772 1708
rect 20824 800 20852 3402
rect 20916 800 20944 4966
rect 21008 3738 21036 23258
rect 21100 22438 21128 38150
rect 21468 33930 21496 38966
rect 22020 37262 22048 39306
rect 22008 37256 22060 37262
rect 22008 37198 22060 37204
rect 22020 35154 22048 37198
rect 22284 37120 22336 37126
rect 22284 37062 22336 37068
rect 22296 36786 22324 37062
rect 22284 36780 22336 36786
rect 22284 36722 22336 36728
rect 22296 36582 22324 36722
rect 22284 36576 22336 36582
rect 22284 36518 22336 36524
rect 22296 36174 22324 36518
rect 22284 36168 22336 36174
rect 22284 36110 22336 36116
rect 22100 36032 22152 36038
rect 22100 35974 22152 35980
rect 22008 35148 22060 35154
rect 22008 35090 22060 35096
rect 21824 34672 21876 34678
rect 21824 34614 21876 34620
rect 21732 34604 21784 34610
rect 21732 34546 21784 34552
rect 21548 34536 21600 34542
rect 21548 34478 21600 34484
rect 21456 33924 21508 33930
rect 21456 33866 21508 33872
rect 21364 32836 21416 32842
rect 21364 32778 21416 32784
rect 21272 27464 21324 27470
rect 21272 27406 21324 27412
rect 21088 22432 21140 22438
rect 21088 22374 21140 22380
rect 21088 21548 21140 21554
rect 21088 21490 21140 21496
rect 21100 21350 21128 21490
rect 21088 21344 21140 21350
rect 21088 21286 21140 21292
rect 21180 21344 21232 21350
rect 21180 21286 21232 21292
rect 21192 19854 21220 21286
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 21088 19712 21140 19718
rect 21088 19654 21140 19660
rect 21100 19514 21128 19654
rect 21088 19508 21140 19514
rect 21088 19450 21140 19456
rect 21284 17218 21312 27406
rect 21376 23322 21404 32778
rect 21468 31346 21496 33866
rect 21456 31340 21508 31346
rect 21456 31282 21508 31288
rect 21456 25492 21508 25498
rect 21456 25434 21508 25440
rect 21468 24886 21496 25434
rect 21456 24880 21508 24886
rect 21456 24822 21508 24828
rect 21560 24138 21588 34478
rect 21640 24200 21692 24206
rect 21640 24142 21692 24148
rect 21548 24132 21600 24138
rect 21548 24074 21600 24080
rect 21652 23594 21680 24142
rect 21640 23588 21692 23594
rect 21640 23530 21692 23536
rect 21364 23316 21416 23322
rect 21364 23258 21416 23264
rect 21652 21078 21680 23530
rect 21744 22438 21772 34546
rect 21836 34202 21864 34614
rect 21824 34196 21876 34202
rect 21824 34138 21876 34144
rect 22020 34066 22048 35090
rect 22112 34542 22140 35974
rect 22296 35850 22324 36110
rect 22296 35822 22416 35850
rect 22388 35494 22416 35822
rect 22376 35488 22428 35494
rect 22376 35430 22428 35436
rect 22192 34944 22244 34950
rect 22192 34886 22244 34892
rect 22204 34610 22232 34886
rect 22192 34604 22244 34610
rect 22192 34546 22244 34552
rect 22100 34536 22152 34542
rect 22100 34478 22152 34484
rect 22008 34060 22060 34066
rect 21928 34020 22008 34048
rect 21928 33522 21956 34020
rect 22008 34002 22060 34008
rect 21916 33516 21968 33522
rect 21916 33458 21968 33464
rect 22100 32768 22152 32774
rect 22100 32710 22152 32716
rect 22112 32434 22140 32710
rect 22100 32428 22152 32434
rect 22100 32370 22152 32376
rect 22388 31754 22416 35430
rect 22480 34474 22508 39306
rect 22572 34950 22600 39374
rect 22664 39098 22692 39986
rect 22756 39370 22784 39986
rect 23032 39642 23060 39986
rect 23020 39636 23072 39642
rect 23020 39578 23072 39584
rect 22744 39364 22796 39370
rect 22744 39306 22796 39312
rect 22652 39092 22704 39098
rect 22652 39034 22704 39040
rect 23124 39030 23152 40394
rect 23296 40384 23348 40390
rect 23216 40344 23296 40372
rect 23216 39438 23244 40344
rect 23296 40326 23348 40332
rect 23204 39432 23256 39438
rect 23204 39374 23256 39380
rect 23400 39302 23428 40462
rect 23572 39840 23624 39846
rect 23572 39782 23624 39788
rect 23480 39636 23532 39642
rect 23480 39578 23532 39584
rect 23388 39296 23440 39302
rect 23388 39238 23440 39244
rect 23112 39024 23164 39030
rect 23112 38966 23164 38972
rect 23020 37664 23072 37670
rect 23020 37606 23072 37612
rect 23032 37398 23060 37606
rect 23020 37392 23072 37398
rect 23020 37334 23072 37340
rect 23032 37126 23060 37334
rect 23400 37262 23428 39238
rect 23492 38554 23520 39578
rect 23584 38962 23612 39782
rect 23572 38956 23624 38962
rect 23572 38898 23624 38904
rect 23480 38548 23532 38554
rect 23480 38490 23532 38496
rect 23480 37936 23532 37942
rect 23480 37878 23532 37884
rect 23388 37256 23440 37262
rect 23388 37198 23440 37204
rect 22928 37120 22980 37126
rect 22928 37062 22980 37068
rect 23020 37120 23072 37126
rect 23020 37062 23072 37068
rect 22652 36576 22704 36582
rect 22652 36518 22704 36524
rect 22560 34944 22612 34950
rect 22560 34886 22612 34892
rect 22468 34468 22520 34474
rect 22468 34410 22520 34416
rect 22296 31726 22416 31754
rect 22100 30184 22152 30190
rect 22100 30126 22152 30132
rect 21914 29336 21970 29345
rect 21914 29271 21970 29280
rect 21928 29238 21956 29271
rect 21916 29232 21968 29238
rect 21916 29174 21968 29180
rect 21914 29064 21970 29073
rect 21836 29022 21914 29050
rect 21836 28966 21864 29022
rect 21914 28999 21970 29008
rect 21824 28960 21876 28966
rect 21824 28902 21876 28908
rect 21916 27328 21968 27334
rect 21916 27270 21968 27276
rect 21824 25764 21876 25770
rect 21824 25706 21876 25712
rect 21836 24818 21864 25706
rect 21824 24812 21876 24818
rect 21928 24800 21956 27270
rect 22112 27062 22140 30126
rect 22190 29472 22246 29481
rect 22190 29407 22246 29416
rect 22204 29238 22232 29407
rect 22192 29232 22244 29238
rect 22192 29174 22244 29180
rect 22296 27878 22324 31726
rect 22480 30802 22508 34410
rect 22572 31822 22600 34886
rect 22560 31816 22612 31822
rect 22560 31758 22612 31764
rect 22572 30870 22600 31758
rect 22560 30864 22612 30870
rect 22560 30806 22612 30812
rect 22468 30796 22520 30802
rect 22468 30738 22520 30744
rect 22376 30592 22428 30598
rect 22376 30534 22428 30540
rect 22388 30258 22416 30534
rect 22376 30252 22428 30258
rect 22376 30194 22428 30200
rect 22480 29782 22508 30738
rect 22560 30320 22612 30326
rect 22560 30262 22612 30268
rect 22468 29776 22520 29782
rect 22468 29718 22520 29724
rect 22376 29708 22428 29714
rect 22376 29650 22428 29656
rect 22388 29170 22416 29650
rect 22572 29646 22600 30262
rect 22560 29640 22612 29646
rect 22560 29582 22612 29588
rect 22468 29504 22520 29510
rect 22468 29446 22520 29452
rect 22376 29164 22428 29170
rect 22376 29106 22428 29112
rect 22284 27872 22336 27878
rect 22284 27814 22336 27820
rect 22100 27056 22152 27062
rect 22100 26998 22152 27004
rect 22112 26586 22140 26998
rect 22100 26580 22152 26586
rect 22100 26522 22152 26528
rect 22192 26512 22244 26518
rect 22192 26454 22244 26460
rect 22204 26314 22232 26454
rect 22192 26308 22244 26314
rect 22192 26250 22244 26256
rect 22100 26036 22152 26042
rect 22100 25978 22152 25984
rect 22112 25770 22140 25978
rect 22192 25900 22244 25906
rect 22192 25842 22244 25848
rect 22100 25764 22152 25770
rect 22100 25706 22152 25712
rect 22008 24812 22060 24818
rect 21928 24772 22008 24800
rect 21824 24754 21876 24760
rect 22008 24754 22060 24760
rect 21836 24426 21864 24754
rect 22112 24682 22140 25706
rect 22204 25158 22232 25842
rect 22192 25152 22244 25158
rect 22192 25094 22244 25100
rect 22100 24676 22152 24682
rect 22100 24618 22152 24624
rect 22190 24576 22246 24585
rect 22190 24511 22246 24520
rect 21836 24398 22140 24426
rect 21824 24064 21876 24070
rect 21824 24006 21876 24012
rect 21916 24064 21968 24070
rect 21916 24006 21968 24012
rect 21836 22642 21864 24006
rect 21824 22636 21876 22642
rect 21824 22578 21876 22584
rect 21732 22432 21784 22438
rect 21732 22374 21784 22380
rect 21928 22030 21956 24006
rect 22008 22636 22060 22642
rect 22008 22578 22060 22584
rect 21916 22024 21968 22030
rect 21916 21966 21968 21972
rect 22020 21146 22048 22578
rect 22112 21690 22140 24398
rect 22204 24274 22232 24511
rect 22192 24268 22244 24274
rect 22192 24210 22244 24216
rect 22296 22778 22324 27814
rect 22376 27600 22428 27606
rect 22376 27542 22428 27548
rect 22284 22772 22336 22778
rect 22284 22714 22336 22720
rect 22100 21684 22152 21690
rect 22100 21626 22152 21632
rect 22008 21140 22060 21146
rect 22008 21082 22060 21088
rect 21640 21072 21692 21078
rect 21640 21014 21692 21020
rect 21916 19508 21968 19514
rect 21916 19450 21968 19456
rect 21928 18834 21956 19450
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 21916 18828 21968 18834
rect 21916 18770 21968 18776
rect 22112 18290 22140 19314
rect 22388 19310 22416 27542
rect 22480 23730 22508 29446
rect 22572 29102 22600 29582
rect 22560 29096 22612 29102
rect 22560 29038 22612 29044
rect 22572 28150 22600 29038
rect 22560 28144 22612 28150
rect 22560 28086 22612 28092
rect 22560 27396 22612 27402
rect 22560 27338 22612 27344
rect 22572 26790 22600 27338
rect 22560 26784 22612 26790
rect 22560 26726 22612 26732
rect 22572 23730 22600 26726
rect 22664 24206 22692 36518
rect 22744 35080 22796 35086
rect 22744 35022 22796 35028
rect 22756 34610 22784 35022
rect 22744 34604 22796 34610
rect 22744 34546 22796 34552
rect 22836 34400 22888 34406
rect 22836 34342 22888 34348
rect 22848 33998 22876 34342
rect 22836 33992 22888 33998
rect 22836 33934 22888 33940
rect 22744 31136 22796 31142
rect 22744 31078 22796 31084
rect 22756 30734 22784 31078
rect 22744 30728 22796 30734
rect 22744 30670 22796 30676
rect 22940 28234 22968 37062
rect 23032 36786 23060 37062
rect 23020 36780 23072 36786
rect 23020 36722 23072 36728
rect 23032 36106 23060 36722
rect 23492 36174 23520 37878
rect 23584 36786 23612 38898
rect 23572 36780 23624 36786
rect 23572 36722 23624 36728
rect 23664 36304 23716 36310
rect 23664 36246 23716 36252
rect 23480 36168 23532 36174
rect 23480 36110 23532 36116
rect 23020 36100 23072 36106
rect 23020 36042 23072 36048
rect 23032 35494 23060 36042
rect 23492 35766 23520 36110
rect 23676 36038 23704 36246
rect 23664 36032 23716 36038
rect 23664 35974 23716 35980
rect 23480 35760 23532 35766
rect 23480 35702 23532 35708
rect 23020 35488 23072 35494
rect 23020 35430 23072 35436
rect 23032 31754 23060 35430
rect 23492 33998 23520 35702
rect 23676 35698 23704 35974
rect 23664 35692 23716 35698
rect 23664 35634 23716 35640
rect 23480 33992 23532 33998
rect 23480 33934 23532 33940
rect 23492 32910 23520 33934
rect 23664 33312 23716 33318
rect 23664 33254 23716 33260
rect 23480 32904 23532 32910
rect 23480 32846 23532 32852
rect 23492 32298 23520 32846
rect 23676 32842 23704 33254
rect 23664 32836 23716 32842
rect 23664 32778 23716 32784
rect 23480 32292 23532 32298
rect 23480 32234 23532 32240
rect 23768 32230 23796 40938
rect 23848 39432 23900 39438
rect 23848 39374 23900 39380
rect 23860 38758 23888 39374
rect 23848 38752 23900 38758
rect 23848 38694 23900 38700
rect 24136 37874 24164 41210
rect 24124 37868 24176 37874
rect 24124 37810 24176 37816
rect 24136 37670 24164 37810
rect 24124 37664 24176 37670
rect 24124 37606 24176 37612
rect 23848 36100 23900 36106
rect 23848 36042 23900 36048
rect 23860 35154 23888 36042
rect 23848 35148 23900 35154
rect 23848 35090 23900 35096
rect 23940 34944 23992 34950
rect 23940 34886 23992 34892
rect 23848 33380 23900 33386
rect 23848 33322 23900 33328
rect 23756 32224 23808 32230
rect 23756 32166 23808 32172
rect 23756 32020 23808 32026
rect 23756 31962 23808 31968
rect 23768 31754 23796 31962
rect 23032 31726 23152 31754
rect 23124 29034 23152 31726
rect 23676 31726 23796 31754
rect 23388 31340 23440 31346
rect 23388 31282 23440 31288
rect 23204 30184 23256 30190
rect 23204 30126 23256 30132
rect 23216 29578 23244 30126
rect 23400 30122 23428 31282
rect 23388 30116 23440 30122
rect 23388 30058 23440 30064
rect 23400 29646 23428 30058
rect 23388 29640 23440 29646
rect 23388 29582 23440 29588
rect 23480 29640 23532 29646
rect 23480 29582 23532 29588
rect 23204 29572 23256 29578
rect 23204 29514 23256 29520
rect 23216 29170 23244 29514
rect 23204 29164 23256 29170
rect 23204 29106 23256 29112
rect 23112 29028 23164 29034
rect 23112 28970 23164 28976
rect 22848 28206 22968 28234
rect 22744 27328 22796 27334
rect 22744 27270 22796 27276
rect 22756 26246 22784 27270
rect 22744 26240 22796 26246
rect 22744 26182 22796 26188
rect 22756 24342 22784 26182
rect 22848 24818 22876 28206
rect 22928 27056 22980 27062
rect 22928 26998 22980 27004
rect 22940 25362 22968 26998
rect 22928 25356 22980 25362
rect 22928 25298 22980 25304
rect 23020 25152 23072 25158
rect 23020 25094 23072 25100
rect 23032 24818 23060 25094
rect 22836 24812 22888 24818
rect 22836 24754 22888 24760
rect 23020 24812 23072 24818
rect 23020 24754 23072 24760
rect 22744 24336 22796 24342
rect 22744 24278 22796 24284
rect 22652 24200 22704 24206
rect 22652 24142 22704 24148
rect 22756 24052 22784 24278
rect 22664 24024 22784 24052
rect 22468 23724 22520 23730
rect 22468 23666 22520 23672
rect 22560 23724 22612 23730
rect 22560 23666 22612 23672
rect 22468 22432 22520 22438
rect 22468 22374 22520 22380
rect 22560 22432 22612 22438
rect 22560 22374 22612 22380
rect 22376 19304 22428 19310
rect 22376 19246 22428 19252
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 21916 18216 21968 18222
rect 21916 18158 21968 18164
rect 21928 18086 21956 18158
rect 21916 18080 21968 18086
rect 21916 18022 21968 18028
rect 21824 17604 21876 17610
rect 21824 17546 21876 17552
rect 21836 17338 21864 17546
rect 21824 17332 21876 17338
rect 21824 17274 21876 17280
rect 21914 17232 21970 17241
rect 21284 17190 21496 17218
rect 21272 16992 21324 16998
rect 21272 16934 21324 16940
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 21192 15162 21220 15302
rect 21180 15156 21232 15162
rect 21180 15098 21232 15104
rect 21192 15026 21220 15098
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 21100 12306 21128 14554
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 21192 11354 21220 11834
rect 21284 11558 21312 16934
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21272 11280 21324 11286
rect 21272 11222 21324 11228
rect 21284 10266 21312 11222
rect 21468 11082 21496 17190
rect 21914 17167 21970 17176
rect 21928 17134 21956 17167
rect 21916 17128 21968 17134
rect 21916 17070 21968 17076
rect 22112 16658 22140 18226
rect 22192 17536 22244 17542
rect 22244 17496 22324 17524
rect 22192 17478 22244 17484
rect 22296 17202 22324 17496
rect 22284 17196 22336 17202
rect 22284 17138 22336 17144
rect 22284 17060 22336 17066
rect 22284 17002 22336 17008
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 22112 15706 22140 16050
rect 22100 15700 22152 15706
rect 22100 15642 22152 15648
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21652 12434 21680 15438
rect 22112 15434 22140 15642
rect 22100 15428 22152 15434
rect 22100 15370 22152 15376
rect 22192 15428 22244 15434
rect 22192 15370 22244 15376
rect 22204 15314 22232 15370
rect 22112 15286 22232 15314
rect 22112 15026 22140 15286
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 21732 14408 21784 14414
rect 21732 14350 21784 14356
rect 21916 14408 21968 14414
rect 21916 14350 21968 14356
rect 21744 13870 21772 14350
rect 21928 14074 21956 14350
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 22112 13938 22140 14962
rect 22190 14920 22246 14929
rect 22190 14855 22192 14864
rect 22244 14855 22246 14864
rect 22192 14826 22244 14832
rect 22296 14618 22324 17002
rect 22480 16794 22508 22374
rect 22572 22030 22600 22374
rect 22664 22234 22692 24024
rect 23124 23866 23152 28970
rect 23492 28490 23520 29582
rect 23676 29510 23704 31726
rect 23860 31346 23888 33322
rect 23848 31340 23900 31346
rect 23848 31282 23900 31288
rect 23860 30138 23888 31282
rect 23952 31226 23980 34886
rect 24032 32428 24084 32434
rect 24032 32370 24084 32376
rect 24044 31346 24072 32370
rect 24136 32026 24164 37606
rect 24320 34950 24348 41686
rect 24768 39840 24820 39846
rect 24768 39782 24820 39788
rect 24780 39370 24808 39782
rect 24768 39364 24820 39370
rect 24768 39306 24820 39312
rect 24676 38344 24728 38350
rect 24780 38332 24808 39306
rect 24728 38304 24808 38332
rect 24676 38286 24728 38292
rect 24400 38276 24452 38282
rect 24400 38218 24452 38224
rect 24412 38010 24440 38218
rect 24400 38004 24452 38010
rect 24400 37946 24452 37952
rect 24676 37732 24728 37738
rect 24676 37674 24728 37680
rect 24584 37664 24636 37670
rect 24584 37606 24636 37612
rect 24596 37194 24624 37606
rect 24584 37188 24636 37194
rect 24584 37130 24636 37136
rect 24492 37120 24544 37126
rect 24492 37062 24544 37068
rect 24504 36718 24532 37062
rect 24492 36712 24544 36718
rect 24492 36654 24544 36660
rect 24504 36174 24532 36654
rect 24492 36168 24544 36174
rect 24492 36110 24544 36116
rect 24400 36032 24452 36038
rect 24400 35974 24452 35980
rect 24412 35698 24440 35974
rect 24688 35834 24716 37674
rect 24780 37262 24808 38304
rect 24952 37868 25004 37874
rect 24952 37810 25004 37816
rect 24768 37256 24820 37262
rect 24768 37198 24820 37204
rect 24780 36922 24808 37198
rect 24768 36916 24820 36922
rect 24768 36858 24820 36864
rect 24676 35828 24728 35834
rect 24676 35770 24728 35776
rect 24400 35692 24452 35698
rect 24400 35634 24452 35640
rect 24412 35086 24440 35634
rect 24688 35086 24716 35770
rect 24400 35080 24452 35086
rect 24400 35022 24452 35028
rect 24676 35080 24728 35086
rect 24676 35022 24728 35028
rect 24308 34944 24360 34950
rect 24308 34886 24360 34892
rect 24492 33856 24544 33862
rect 24492 33798 24544 33804
rect 24400 33516 24452 33522
rect 24400 33458 24452 33464
rect 24308 33380 24360 33386
rect 24308 33322 24360 33328
rect 24320 32978 24348 33322
rect 24412 33114 24440 33458
rect 24400 33108 24452 33114
rect 24400 33050 24452 33056
rect 24308 32972 24360 32978
rect 24308 32914 24360 32920
rect 24216 32836 24268 32842
rect 24216 32778 24268 32784
rect 24124 32020 24176 32026
rect 24124 31962 24176 31968
rect 24032 31340 24084 31346
rect 24032 31282 24084 31288
rect 23952 31198 24072 31226
rect 24044 31142 24072 31198
rect 24032 31136 24084 31142
rect 24032 31078 24084 31084
rect 23860 30110 23980 30138
rect 23848 30048 23900 30054
rect 23848 29990 23900 29996
rect 23664 29504 23716 29510
rect 23664 29446 23716 29452
rect 23676 29102 23704 29446
rect 23756 29300 23808 29306
rect 23756 29242 23808 29248
rect 23664 29096 23716 29102
rect 23664 29038 23716 29044
rect 23768 28626 23796 29242
rect 23756 28620 23808 28626
rect 23756 28562 23808 28568
rect 23480 28484 23532 28490
rect 23480 28426 23532 28432
rect 23480 26988 23532 26994
rect 23480 26930 23532 26936
rect 23204 25696 23256 25702
rect 23204 25638 23256 25644
rect 23216 25294 23244 25638
rect 23204 25288 23256 25294
rect 23204 25230 23256 25236
rect 23204 24812 23256 24818
rect 23204 24754 23256 24760
rect 23388 24812 23440 24818
rect 23388 24754 23440 24760
rect 23216 24138 23244 24754
rect 23204 24132 23256 24138
rect 23204 24074 23256 24080
rect 23112 23860 23164 23866
rect 23112 23802 23164 23808
rect 23216 23798 23244 24074
rect 23204 23792 23256 23798
rect 23204 23734 23256 23740
rect 23400 23730 23428 24754
rect 23492 24614 23520 26930
rect 23572 25492 23624 25498
rect 23572 25434 23624 25440
rect 23584 24886 23612 25434
rect 23572 24880 23624 24886
rect 23572 24822 23624 24828
rect 23480 24608 23532 24614
rect 23480 24550 23532 24556
rect 23572 24608 23624 24614
rect 23572 24550 23624 24556
rect 23388 23724 23440 23730
rect 23388 23666 23440 23672
rect 23400 23594 23428 23666
rect 23388 23588 23440 23594
rect 23388 23530 23440 23536
rect 22836 23520 22888 23526
rect 22836 23462 22888 23468
rect 22848 23118 22876 23462
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 22928 22976 22980 22982
rect 22928 22918 22980 22924
rect 22652 22228 22704 22234
rect 22652 22170 22704 22176
rect 22560 22024 22612 22030
rect 22560 21966 22612 21972
rect 22664 21554 22692 22170
rect 22744 21888 22796 21894
rect 22744 21830 22796 21836
rect 22652 21548 22704 21554
rect 22652 21490 22704 21496
rect 22664 20806 22692 21490
rect 22756 20874 22784 21830
rect 22836 21548 22888 21554
rect 22836 21490 22888 21496
rect 22744 20868 22796 20874
rect 22744 20810 22796 20816
rect 22652 20800 22704 20806
rect 22652 20742 22704 20748
rect 22848 20058 22876 21490
rect 22836 20052 22888 20058
rect 22836 19994 22888 20000
rect 22940 17218 22968 22918
rect 23584 22642 23612 24550
rect 23572 22636 23624 22642
rect 23572 22578 23624 22584
rect 23112 22568 23164 22574
rect 23112 22510 23164 22516
rect 23124 22008 23152 22510
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 23400 22234 23428 22374
rect 23388 22228 23440 22234
rect 23388 22170 23440 22176
rect 23400 22030 23428 22170
rect 23204 22024 23256 22030
rect 23112 22002 23164 22008
rect 23204 21966 23256 21972
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 23112 21944 23164 21950
rect 23124 21622 23152 21944
rect 23216 21690 23244 21966
rect 23204 21684 23256 21690
rect 23204 21626 23256 21632
rect 23112 21616 23164 21622
rect 23032 21576 23112 21604
rect 23032 19514 23060 21576
rect 23112 21558 23164 21564
rect 23664 21616 23716 21622
rect 23664 21558 23716 21564
rect 23204 21412 23256 21418
rect 23204 21354 23256 21360
rect 23216 20942 23244 21354
rect 23296 21344 23348 21350
rect 23296 21286 23348 21292
rect 23204 20936 23256 20942
rect 23204 20878 23256 20884
rect 23112 20460 23164 20466
rect 23216 20448 23244 20878
rect 23308 20534 23336 21286
rect 23388 20868 23440 20874
rect 23388 20810 23440 20816
rect 23296 20528 23348 20534
rect 23296 20470 23348 20476
rect 23164 20420 23244 20448
rect 23112 20402 23164 20408
rect 23020 19508 23072 19514
rect 23020 19450 23072 19456
rect 23020 18896 23072 18902
rect 23020 18838 23072 18844
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22848 17190 22968 17218
rect 22572 17066 22600 17138
rect 22560 17060 22612 17066
rect 22560 17002 22612 17008
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 22100 13932 22152 13938
rect 22100 13874 22152 13880
rect 21732 13864 21784 13870
rect 21732 13806 21784 13812
rect 22100 13252 22152 13258
rect 22100 13194 22152 13200
rect 22112 12850 22140 13194
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22008 12640 22060 12646
rect 22008 12582 22060 12588
rect 21652 12406 21772 12434
rect 21548 12096 21600 12102
rect 21548 12038 21600 12044
rect 21560 11830 21588 12038
rect 21548 11824 21600 11830
rect 21548 11766 21600 11772
rect 21640 11688 21692 11694
rect 21640 11630 21692 11636
rect 21652 11218 21680 11630
rect 21640 11212 21692 11218
rect 21640 11154 21692 11160
rect 21456 11076 21508 11082
rect 21456 11018 21508 11024
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21284 10130 21312 10202
rect 21272 10124 21324 10130
rect 21272 10066 21324 10072
rect 21744 8974 21772 12406
rect 22020 12238 22048 12582
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 21836 12050 21864 12174
rect 22112 12050 22140 12786
rect 22572 12442 22600 17002
rect 22744 16652 22796 16658
rect 22744 16594 22796 16600
rect 22756 15094 22784 16594
rect 22744 15088 22796 15094
rect 22744 15030 22796 15036
rect 22756 14550 22784 15030
rect 22744 14544 22796 14550
rect 22744 14486 22796 14492
rect 22756 14074 22784 14486
rect 22744 14068 22796 14074
rect 22744 14010 22796 14016
rect 22560 12436 22612 12442
rect 22560 12378 22612 12384
rect 22572 12238 22600 12378
rect 22560 12232 22612 12238
rect 22560 12174 22612 12180
rect 21836 12022 22140 12050
rect 22112 11762 22140 12022
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22480 11558 22508 11834
rect 22652 11756 22704 11762
rect 22652 11698 22704 11704
rect 22192 11552 22244 11558
rect 22192 11494 22244 11500
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22204 11082 22232 11494
rect 22192 11076 22244 11082
rect 22192 11018 22244 11024
rect 22664 10810 22692 11698
rect 22744 11688 22796 11694
rect 22744 11630 22796 11636
rect 22756 11354 22784 11630
rect 22744 11348 22796 11354
rect 22744 11290 22796 11296
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 22192 10668 22244 10674
rect 22192 10610 22244 10616
rect 22204 10266 22232 10610
rect 22848 10538 22876 17190
rect 23032 17134 23060 18838
rect 23400 18834 23428 20810
rect 23676 19786 23704 21558
rect 23860 21486 23888 29990
rect 23952 22094 23980 30110
rect 24044 24954 24072 31078
rect 24124 30660 24176 30666
rect 24124 30602 24176 30608
rect 24136 26790 24164 30602
rect 24228 30326 24256 32778
rect 24320 32570 24348 32914
rect 24308 32564 24360 32570
rect 24308 32506 24360 32512
rect 24308 32428 24360 32434
rect 24308 32370 24360 32376
rect 24320 30734 24348 32370
rect 24400 32224 24452 32230
rect 24400 32166 24452 32172
rect 24308 30728 24360 30734
rect 24308 30670 24360 30676
rect 24216 30320 24268 30326
rect 24216 30262 24268 30268
rect 24412 29866 24440 32166
rect 24504 30258 24532 33798
rect 24688 33590 24716 35022
rect 24768 34400 24820 34406
rect 24768 34342 24820 34348
rect 24676 33584 24728 33590
rect 24676 33526 24728 33532
rect 24688 31890 24716 33526
rect 24780 33454 24808 34342
rect 24964 33522 24992 37810
rect 25044 37188 25096 37194
rect 25044 37130 25096 37136
rect 25056 35290 25084 37130
rect 25044 35284 25096 35290
rect 25044 35226 25096 35232
rect 25044 33924 25096 33930
rect 25044 33866 25096 33872
rect 24952 33516 25004 33522
rect 24952 33458 25004 33464
rect 24768 33448 24820 33454
rect 24768 33390 24820 33396
rect 24780 32473 24808 33390
rect 24964 32978 24992 33458
rect 24952 32972 25004 32978
rect 24952 32914 25004 32920
rect 24766 32464 24822 32473
rect 24766 32399 24822 32408
rect 24676 31884 24728 31890
rect 24676 31826 24728 31832
rect 24584 30728 24636 30734
rect 24584 30670 24636 30676
rect 24492 30252 24544 30258
rect 24492 30194 24544 30200
rect 24228 29838 24440 29866
rect 24124 26784 24176 26790
rect 24124 26726 24176 26732
rect 24136 25498 24164 26726
rect 24124 25492 24176 25498
rect 24124 25434 24176 25440
rect 24032 24948 24084 24954
rect 24032 24890 24084 24896
rect 24228 23769 24256 29838
rect 24400 29572 24452 29578
rect 24400 29514 24452 29520
rect 24412 29306 24440 29514
rect 24492 29504 24544 29510
rect 24492 29446 24544 29452
rect 24504 29345 24532 29446
rect 24490 29336 24546 29345
rect 24400 29300 24452 29306
rect 24490 29271 24546 29280
rect 24400 29242 24452 29248
rect 24504 29238 24532 29271
rect 24492 29232 24544 29238
rect 24492 29174 24544 29180
rect 24596 29170 24624 30670
rect 24676 30660 24728 30666
rect 24676 30602 24728 30608
rect 24688 29889 24716 30602
rect 24674 29880 24730 29889
rect 24674 29815 24730 29824
rect 24308 29164 24360 29170
rect 24308 29106 24360 29112
rect 24584 29164 24636 29170
rect 24584 29106 24636 29112
rect 24320 26518 24348 29106
rect 24780 28694 24808 32399
rect 24860 31816 24912 31822
rect 24860 31758 24912 31764
rect 24872 30190 24900 31758
rect 24964 30258 24992 32914
rect 25056 32774 25084 33866
rect 25044 32768 25096 32774
rect 25044 32710 25096 32716
rect 24952 30252 25004 30258
rect 24952 30194 25004 30200
rect 24860 30184 24912 30190
rect 24860 30126 24912 30132
rect 24964 29714 24992 30194
rect 25056 29782 25084 32710
rect 25044 29776 25096 29782
rect 25044 29718 25096 29724
rect 24952 29708 25004 29714
rect 24952 29650 25004 29656
rect 25044 29640 25096 29646
rect 25044 29582 25096 29588
rect 25056 29306 25084 29582
rect 25044 29300 25096 29306
rect 25044 29242 25096 29248
rect 24768 28688 24820 28694
rect 24768 28630 24820 28636
rect 24860 28552 24912 28558
rect 24860 28494 24912 28500
rect 24872 27878 24900 28494
rect 24860 27872 24912 27878
rect 24860 27814 24912 27820
rect 24768 27328 24820 27334
rect 24768 27270 24820 27276
rect 24780 26994 24808 27270
rect 25044 27124 25096 27130
rect 25044 27066 25096 27072
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24584 26920 24636 26926
rect 24584 26862 24636 26868
rect 24308 26512 24360 26518
rect 24308 26454 24360 26460
rect 24596 26450 24624 26862
rect 25056 26586 25084 27066
rect 25044 26580 25096 26586
rect 25044 26522 25096 26528
rect 24584 26444 24636 26450
rect 24584 26386 24636 26392
rect 24492 26376 24544 26382
rect 24492 26318 24544 26324
rect 24504 25906 24532 26318
rect 24596 25974 24624 26386
rect 24676 26376 24728 26382
rect 24728 26324 24900 26330
rect 24676 26318 24900 26324
rect 24688 26302 24900 26318
rect 24584 25968 24636 25974
rect 24584 25910 24636 25916
rect 24492 25900 24544 25906
rect 24492 25842 24544 25848
rect 24504 25226 24532 25842
rect 24872 25498 24900 26302
rect 24860 25492 24912 25498
rect 24860 25434 24912 25440
rect 24492 25220 24544 25226
rect 24492 25162 24544 25168
rect 24504 24206 24532 25162
rect 24492 24200 24544 24206
rect 24492 24142 24544 24148
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 24584 24132 24636 24138
rect 24584 24074 24636 24080
rect 24596 23866 24624 24074
rect 24584 23860 24636 23866
rect 24584 23802 24636 23808
rect 24492 23792 24544 23798
rect 24214 23760 24270 23769
rect 24214 23695 24270 23704
rect 24490 23760 24492 23769
rect 24544 23760 24546 23769
rect 24490 23695 24546 23704
rect 24492 23044 24544 23050
rect 24492 22986 24544 22992
rect 23952 22066 24164 22094
rect 23940 21548 23992 21554
rect 23940 21490 23992 21496
rect 23848 21480 23900 21486
rect 23848 21422 23900 21428
rect 23952 20806 23980 21490
rect 23940 20800 23992 20806
rect 23940 20742 23992 20748
rect 23664 19780 23716 19786
rect 23664 19722 23716 19728
rect 23388 18828 23440 18834
rect 23388 18770 23440 18776
rect 23388 18284 23440 18290
rect 23388 18226 23440 18232
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 23020 17128 23072 17134
rect 23020 17070 23072 17076
rect 22928 16652 22980 16658
rect 22928 16594 22980 16600
rect 22836 10532 22888 10538
rect 22836 10474 22888 10480
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 22100 10056 22152 10062
rect 22100 9998 22152 10004
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21732 8968 21784 8974
rect 21732 8910 21784 8916
rect 21284 8634 21312 8910
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 21836 8498 21864 8978
rect 22112 8498 22140 9998
rect 22468 9920 22520 9926
rect 22468 9862 22520 9868
rect 22284 9648 22336 9654
rect 22284 9590 22336 9596
rect 22296 9178 22324 9590
rect 22480 9586 22508 9862
rect 22468 9580 22520 9586
rect 22468 9522 22520 9528
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 22284 9172 22336 9178
rect 22284 9114 22336 9120
rect 21364 8492 21416 8498
rect 21364 8434 21416 8440
rect 21824 8492 21876 8498
rect 21824 8434 21876 8440
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21284 6866 21312 7686
rect 21376 7449 21404 8434
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 21362 7440 21418 7449
rect 21362 7375 21364 7384
rect 21416 7375 21418 7384
rect 21364 7346 21416 7352
rect 22112 7342 22140 7822
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 21272 6860 21324 6866
rect 21272 6802 21324 6808
rect 22480 6798 22508 9522
rect 22756 9382 22784 9522
rect 22940 9450 22968 16594
rect 23124 16590 23152 17614
rect 23400 17270 23428 18226
rect 23676 18154 23704 19722
rect 23664 18148 23716 18154
rect 23664 18090 23716 18096
rect 23388 17264 23440 17270
rect 23388 17206 23440 17212
rect 23664 17128 23716 17134
rect 23664 17070 23716 17076
rect 23112 16584 23164 16590
rect 23112 16526 23164 16532
rect 23124 16250 23152 16526
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 23388 16244 23440 16250
rect 23388 16186 23440 16192
rect 23112 14816 23164 14822
rect 23112 14758 23164 14764
rect 23124 14074 23152 14758
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 23204 13728 23256 13734
rect 23204 13670 23256 13676
rect 23216 13530 23244 13670
rect 23204 13524 23256 13530
rect 23204 13466 23256 13472
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 23112 13184 23164 13190
rect 23112 13126 23164 13132
rect 23020 11008 23072 11014
rect 23020 10950 23072 10956
rect 23032 10742 23060 10950
rect 23020 10736 23072 10742
rect 23020 10678 23072 10684
rect 23032 9654 23060 10678
rect 23020 9648 23072 9654
rect 23020 9590 23072 9596
rect 22928 9444 22980 9450
rect 22928 9386 22980 9392
rect 22744 9376 22796 9382
rect 22744 9318 22796 9324
rect 22756 9042 22784 9318
rect 22744 9036 22796 9042
rect 22744 8978 22796 8984
rect 22652 8492 22704 8498
rect 22652 8434 22704 8440
rect 22560 7744 22612 7750
rect 22560 7686 22612 7692
rect 22572 7478 22600 7686
rect 22560 7472 22612 7478
rect 22560 7414 22612 7420
rect 22664 7410 22692 8434
rect 23124 7546 23152 13126
rect 23216 10810 23244 13262
rect 23400 13258 23428 16186
rect 23480 16176 23532 16182
rect 23480 16118 23532 16124
rect 23492 15026 23520 16118
rect 23676 16114 23704 17070
rect 23664 16108 23716 16114
rect 23664 16050 23716 16056
rect 23572 16040 23624 16046
rect 23572 15982 23624 15988
rect 23480 15020 23532 15026
rect 23480 14962 23532 14968
rect 23584 14958 23612 15982
rect 23676 15706 23704 16050
rect 23664 15700 23716 15706
rect 23664 15642 23716 15648
rect 23848 15428 23900 15434
rect 23848 15370 23900 15376
rect 23860 15026 23888 15370
rect 23848 15020 23900 15026
rect 23848 14962 23900 14968
rect 23572 14952 23624 14958
rect 23492 14900 23572 14906
rect 23492 14894 23624 14900
rect 23492 14878 23612 14894
rect 23492 14414 23520 14878
rect 23572 14816 23624 14822
rect 23572 14758 23624 14764
rect 23848 14816 23900 14822
rect 23848 14758 23900 14764
rect 23480 14408 23532 14414
rect 23480 14350 23532 14356
rect 23492 13938 23520 14350
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23584 13734 23612 14758
rect 23860 14618 23888 14758
rect 23848 14612 23900 14618
rect 23848 14554 23900 14560
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23572 13728 23624 13734
rect 23572 13670 23624 13676
rect 23676 13530 23704 14214
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23388 13252 23440 13258
rect 23388 13194 23440 13200
rect 23572 11892 23624 11898
rect 23572 11834 23624 11840
rect 23584 11218 23612 11834
rect 23664 11756 23716 11762
rect 23664 11698 23716 11704
rect 23676 11558 23704 11698
rect 23664 11552 23716 11558
rect 23664 11494 23716 11500
rect 23572 11212 23624 11218
rect 23572 11154 23624 11160
rect 23676 11150 23704 11494
rect 23480 11144 23532 11150
rect 23400 11104 23480 11132
rect 23204 10804 23256 10810
rect 23204 10746 23256 10752
rect 23400 10062 23428 11104
rect 23480 11086 23532 11092
rect 23664 11144 23716 11150
rect 23664 11086 23716 11092
rect 23388 10056 23440 10062
rect 23388 9998 23440 10004
rect 23664 9172 23716 9178
rect 23664 9114 23716 9120
rect 23676 8498 23704 9114
rect 23664 8492 23716 8498
rect 23664 8434 23716 8440
rect 23296 8424 23348 8430
rect 23296 8366 23348 8372
rect 23204 8288 23256 8294
rect 23204 8230 23256 8236
rect 23216 7886 23244 8230
rect 23204 7880 23256 7886
rect 23204 7822 23256 7828
rect 23308 7546 23336 8366
rect 23480 8356 23532 8362
rect 23480 8298 23532 8304
rect 23112 7540 23164 7546
rect 23112 7482 23164 7488
rect 23296 7540 23348 7546
rect 23296 7482 23348 7488
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 23388 7404 23440 7410
rect 23388 7346 23440 7352
rect 22744 7336 22796 7342
rect 22744 7278 22796 7284
rect 21732 6792 21784 6798
rect 21732 6734 21784 6740
rect 22468 6792 22520 6798
rect 22468 6734 22520 6740
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 21284 6118 21312 6394
rect 21744 6254 21772 6734
rect 22756 6254 22784 7278
rect 23204 6656 23256 6662
rect 23204 6598 23256 6604
rect 21732 6248 21784 6254
rect 21732 6190 21784 6196
rect 22744 6248 22796 6254
rect 22744 6190 22796 6196
rect 21272 6112 21324 6118
rect 21272 6054 21324 6060
rect 21364 5568 21416 5574
rect 21364 5510 21416 5516
rect 20996 3732 21048 3738
rect 20996 3674 21048 3680
rect 21088 3732 21140 3738
rect 21088 3674 21140 3680
rect 20994 3224 21050 3233
rect 21100 3194 21128 3674
rect 21180 3596 21232 3602
rect 21180 3538 21232 3544
rect 20994 3159 21050 3168
rect 21088 3188 21140 3194
rect 21008 3126 21036 3159
rect 21088 3130 21140 3136
rect 20996 3120 21048 3126
rect 20996 3062 21048 3068
rect 21088 1760 21140 1766
rect 21088 1702 21140 1708
rect 21100 800 21128 1702
rect 21192 800 21220 3538
rect 21376 3126 21404 5510
rect 21548 5296 21600 5302
rect 21548 5238 21600 5244
rect 21456 4004 21508 4010
rect 21456 3946 21508 3952
rect 21364 3120 21416 3126
rect 21364 3062 21416 3068
rect 21270 2680 21326 2689
rect 21270 2615 21326 2624
rect 21284 2582 21312 2615
rect 21272 2576 21324 2582
rect 21272 2518 21324 2524
rect 21376 800 21404 3062
rect 21468 800 21496 3946
rect 21560 3602 21588 5238
rect 21744 4758 21772 6190
rect 22756 5710 22784 6190
rect 22744 5704 22796 5710
rect 22744 5646 22796 5652
rect 21916 5568 21968 5574
rect 21916 5510 21968 5516
rect 22926 5536 22982 5545
rect 21824 5024 21876 5030
rect 21824 4966 21876 4972
rect 21732 4752 21784 4758
rect 21732 4694 21784 4700
rect 21732 4616 21784 4622
rect 21732 4558 21784 4564
rect 21548 3596 21600 3602
rect 21548 3538 21600 3544
rect 21640 3528 21692 3534
rect 21640 3470 21692 3476
rect 21652 800 21680 3470
rect 21744 800 21772 4558
rect 21836 3534 21864 4966
rect 21824 3528 21876 3534
rect 21824 3470 21876 3476
rect 21928 2378 21956 5510
rect 22926 5471 22982 5480
rect 22192 5160 22244 5166
rect 22192 5102 22244 5108
rect 22100 4208 22152 4214
rect 22100 4150 22152 4156
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 21916 2372 21968 2378
rect 21916 2314 21968 2320
rect 21928 800 21956 2314
rect 22020 800 22048 3878
rect 22112 2446 22140 4150
rect 22204 3126 22232 5102
rect 22652 5092 22704 5098
rect 22652 5034 22704 5040
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 22192 3120 22244 3126
rect 22192 3062 22244 3068
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 22204 800 22232 3062
rect 22296 800 22324 4966
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 22374 3224 22430 3233
rect 22374 3159 22430 3168
rect 22388 3126 22416 3159
rect 22376 3120 22428 3126
rect 22376 3062 22428 3068
rect 22480 2854 22508 3878
rect 22468 2848 22520 2854
rect 22468 2790 22520 2796
rect 22376 2508 22428 2514
rect 22376 2450 22428 2456
rect 22388 1970 22416 2450
rect 22468 2032 22520 2038
rect 22468 1974 22520 1980
rect 22376 1964 22428 1970
rect 22376 1906 22428 1912
rect 22480 800 22508 1974
rect 22572 800 22600 4558
rect 22664 2446 22692 5034
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22848 3058 22876 3334
rect 22836 3052 22888 3058
rect 22836 2994 22888 3000
rect 22848 2938 22876 2994
rect 22756 2910 22876 2938
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 22664 2038 22692 2382
rect 22652 2032 22704 2038
rect 22652 1974 22704 1980
rect 22756 800 22784 2910
rect 22836 2848 22888 2854
rect 22836 2790 22888 2796
rect 22848 800 22876 2790
rect 22940 2650 22968 5471
rect 23112 4616 23164 4622
rect 23112 4558 23164 4564
rect 23018 3224 23074 3233
rect 23018 3159 23020 3168
rect 23072 3159 23074 3168
rect 23020 3130 23072 3136
rect 22928 2644 22980 2650
rect 22928 2586 22980 2592
rect 23020 2440 23072 2446
rect 23020 2382 23072 2388
rect 23032 800 23060 2382
rect 23124 800 23152 4558
rect 23216 4146 23244 6598
rect 23400 6338 23428 7346
rect 23492 6798 23520 8298
rect 23662 7576 23718 7585
rect 23662 7511 23718 7520
rect 23676 7478 23704 7511
rect 23664 7472 23716 7478
rect 23664 7414 23716 7420
rect 23480 6792 23532 6798
rect 23664 6792 23716 6798
rect 23532 6752 23612 6780
rect 23480 6734 23532 6740
rect 23400 6322 23520 6338
rect 23400 6316 23532 6322
rect 23400 6310 23480 6316
rect 23400 5710 23428 6310
rect 23480 6258 23532 6264
rect 23388 5704 23440 5710
rect 23388 5646 23440 5652
rect 23584 5574 23612 6752
rect 23664 6734 23716 6740
rect 23676 5914 23704 6734
rect 23664 5908 23716 5914
rect 23664 5850 23716 5856
rect 23768 5846 23796 13806
rect 23860 13802 23888 14214
rect 23848 13796 23900 13802
rect 23848 13738 23900 13744
rect 23940 13728 23992 13734
rect 23940 13670 23992 13676
rect 23952 13258 23980 13670
rect 23940 13252 23992 13258
rect 23940 13194 23992 13200
rect 23952 12442 23980 13194
rect 24136 12850 24164 22066
rect 24400 22024 24452 22030
rect 24400 21966 24452 21972
rect 24412 21622 24440 21966
rect 24504 21622 24532 22986
rect 24964 22642 24992 24142
rect 24952 22636 25004 22642
rect 24952 22578 25004 22584
rect 24400 21616 24452 21622
rect 24400 21558 24452 21564
rect 24492 21616 24544 21622
rect 24492 21558 24544 21564
rect 24584 21004 24636 21010
rect 24584 20946 24636 20952
rect 24492 20800 24544 20806
rect 24492 20742 24544 20748
rect 24400 20256 24452 20262
rect 24400 20198 24452 20204
rect 24412 19854 24440 20198
rect 24400 19848 24452 19854
rect 24400 19790 24452 19796
rect 24412 19378 24440 19790
rect 24400 19372 24452 19378
rect 24400 19314 24452 19320
rect 24504 18290 24532 20742
rect 24492 18284 24544 18290
rect 24492 18226 24544 18232
rect 24400 18216 24452 18222
rect 24400 18158 24452 18164
rect 24412 17678 24440 18158
rect 24400 17672 24452 17678
rect 24400 17614 24452 17620
rect 24400 14952 24452 14958
rect 24400 14894 24452 14900
rect 24412 14550 24440 14894
rect 24596 14550 24624 20946
rect 24860 20392 24912 20398
rect 24860 20334 24912 20340
rect 24676 19780 24728 19786
rect 24676 19722 24728 19728
rect 24688 19446 24716 19722
rect 24676 19440 24728 19446
rect 24676 19382 24728 19388
rect 24688 18290 24716 19382
rect 24676 18284 24728 18290
rect 24676 18226 24728 18232
rect 24872 18086 24900 20334
rect 24952 19304 25004 19310
rect 24952 19246 25004 19252
rect 24964 18290 24992 19246
rect 24952 18284 25004 18290
rect 24952 18226 25004 18232
rect 24860 18080 24912 18086
rect 24860 18022 24912 18028
rect 24860 17876 24912 17882
rect 24860 17818 24912 17824
rect 24872 16794 24900 17818
rect 24964 17134 24992 18226
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 24952 17128 25004 17134
rect 24952 17070 25004 17076
rect 25056 16794 25084 18022
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 25044 16788 25096 16794
rect 25044 16730 25096 16736
rect 25044 16584 25096 16590
rect 25042 16552 25044 16561
rect 25096 16552 25098 16561
rect 25042 16487 25098 16496
rect 25044 15020 25096 15026
rect 25044 14962 25096 14968
rect 25056 14550 25084 14962
rect 24400 14544 24452 14550
rect 24400 14486 24452 14492
rect 24584 14544 24636 14550
rect 24584 14486 24636 14492
rect 25044 14544 25096 14550
rect 25044 14486 25096 14492
rect 24308 13796 24360 13802
rect 24308 13738 24360 13744
rect 24216 13320 24268 13326
rect 24216 13262 24268 13268
rect 24124 12844 24176 12850
rect 24124 12786 24176 12792
rect 24032 12776 24084 12782
rect 24032 12718 24084 12724
rect 23940 12436 23992 12442
rect 23940 12378 23992 12384
rect 24044 10062 24072 12718
rect 24032 10056 24084 10062
rect 24032 9998 24084 10004
rect 24044 8498 24072 9998
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 24044 7410 24072 8434
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 23940 7336 23992 7342
rect 23940 7278 23992 7284
rect 23952 6730 23980 7278
rect 24044 6798 24072 7346
rect 24032 6792 24084 6798
rect 24032 6734 24084 6740
rect 23940 6724 23992 6730
rect 23940 6666 23992 6672
rect 24228 6458 24256 13262
rect 24320 12782 24348 13738
rect 24308 12776 24360 12782
rect 24308 12718 24360 12724
rect 24412 11762 24440 14486
rect 24596 13870 24624 14486
rect 24584 13864 24636 13870
rect 24584 13806 24636 13812
rect 24584 13320 24636 13326
rect 24584 13262 24636 13268
rect 24596 12714 24624 13262
rect 24860 13184 24912 13190
rect 24860 13126 24912 13132
rect 24676 12844 24728 12850
rect 24676 12786 24728 12792
rect 24584 12708 24636 12714
rect 24584 12650 24636 12656
rect 24688 12434 24716 12786
rect 24504 12406 24716 12434
rect 24504 12102 24532 12406
rect 24492 12096 24544 12102
rect 24492 12038 24544 12044
rect 24400 11756 24452 11762
rect 24400 11698 24452 11704
rect 24504 11286 24532 12038
rect 24492 11280 24544 11286
rect 24492 11222 24544 11228
rect 24584 11212 24636 11218
rect 24584 11154 24636 11160
rect 24596 10674 24624 11154
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24308 10600 24360 10606
rect 24308 10542 24360 10548
rect 24320 10130 24348 10542
rect 24308 10124 24360 10130
rect 24308 10066 24360 10072
rect 24320 8566 24348 10066
rect 24872 9674 24900 13126
rect 24952 12912 25004 12918
rect 24952 12854 25004 12860
rect 24964 12442 24992 12854
rect 24952 12436 25004 12442
rect 24952 12378 25004 12384
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 25044 12232 25096 12238
rect 25044 12174 25096 12180
rect 24964 11558 24992 12174
rect 24952 11552 25004 11558
rect 24952 11494 25004 11500
rect 25056 11082 25084 12174
rect 25044 11076 25096 11082
rect 25044 11018 25096 11024
rect 25056 10674 25084 11018
rect 25044 10668 25096 10674
rect 25044 10610 25096 10616
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 24964 9722 24992 9998
rect 24596 9646 24900 9674
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 24308 8560 24360 8566
rect 24308 8502 24360 8508
rect 24320 7342 24348 8502
rect 24308 7336 24360 7342
rect 24308 7278 24360 7284
rect 24596 6798 24624 9646
rect 24952 7880 25004 7886
rect 24952 7822 25004 7828
rect 24676 7744 24728 7750
rect 24676 7686 24728 7692
rect 24688 6905 24716 7686
rect 24768 7404 24820 7410
rect 24768 7346 24820 7352
rect 24674 6896 24730 6905
rect 24674 6831 24730 6840
rect 24308 6792 24360 6798
rect 24308 6734 24360 6740
rect 24584 6792 24636 6798
rect 24584 6734 24636 6740
rect 24320 6662 24348 6734
rect 24308 6656 24360 6662
rect 24308 6598 24360 6604
rect 24216 6452 24268 6458
rect 24216 6394 24268 6400
rect 24596 6254 24624 6734
rect 24780 6662 24808 7346
rect 24860 6792 24912 6798
rect 24860 6734 24912 6740
rect 24676 6656 24728 6662
rect 24676 6598 24728 6604
rect 24768 6656 24820 6662
rect 24768 6598 24820 6604
rect 24584 6248 24636 6254
rect 24584 6190 24636 6196
rect 24596 5846 24624 6190
rect 23756 5840 23808 5846
rect 23756 5782 23808 5788
rect 24584 5840 24636 5846
rect 24584 5782 24636 5788
rect 24584 5636 24636 5642
rect 24584 5578 24636 5584
rect 23572 5568 23624 5574
rect 23572 5510 23624 5516
rect 24596 5302 24624 5578
rect 24584 5296 24636 5302
rect 24584 5238 24636 5244
rect 24596 4826 24624 5238
rect 24584 4820 24636 4826
rect 24584 4762 24636 4768
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 23940 4616 23992 4622
rect 23940 4558 23992 4564
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23492 2774 23520 4558
rect 23952 3942 23980 4558
rect 24688 4554 24716 6598
rect 24768 6384 24820 6390
rect 24768 6326 24820 6332
rect 24780 5710 24808 6326
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 24676 4548 24728 4554
rect 24676 4490 24728 4496
rect 24032 4072 24084 4078
rect 24032 4014 24084 4020
rect 23940 3936 23992 3942
rect 23940 3878 23992 3884
rect 23664 3528 23716 3534
rect 23664 3470 23716 3476
rect 23400 2746 23520 2774
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 23308 800 23336 2382
rect 23400 800 23428 2746
rect 23676 800 23704 3470
rect 24044 2774 24072 4014
rect 24780 4010 24808 5646
rect 24872 5370 24900 6734
rect 24964 6118 24992 7822
rect 24952 6112 25004 6118
rect 24952 6054 25004 6060
rect 24860 5364 24912 5370
rect 24860 5306 24912 5312
rect 24964 4622 24992 6054
rect 24952 4616 25004 4622
rect 24952 4558 25004 4564
rect 24768 4004 24820 4010
rect 24768 3946 24820 3952
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 23952 2746 24072 2774
rect 23952 800 23980 2746
rect 24228 800 24256 3470
rect 24492 2984 24544 2990
rect 24492 2926 24544 2932
rect 24504 800 24532 2926
rect 24780 800 24808 3470
rect 25044 2848 25096 2854
rect 25044 2790 25096 2796
rect 25056 800 25084 2790
rect 25148 2106 25176 55558
rect 26068 41682 26096 55558
rect 26804 55321 26832 55558
rect 26790 55312 26846 55321
rect 26790 55247 26846 55256
rect 28000 44849 28028 56102
rect 29196 55622 29224 56306
rect 29932 56273 29960 56306
rect 29918 56264 29974 56273
rect 29918 56199 29920 56208
rect 29972 56199 29974 56208
rect 29920 56170 29972 56176
rect 30392 56166 30420 57462
rect 48700 57458 48728 59200
rect 50264 57882 50292 59200
rect 50172 57854 50292 57882
rect 50172 57458 50200 57854
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 51828 57458 51856 59200
rect 53392 57458 53420 59200
rect 32220 57452 32272 57458
rect 32220 57394 32272 57400
rect 33232 57452 33284 57458
rect 33232 57394 33284 57400
rect 40776 57452 40828 57458
rect 40776 57394 40828 57400
rect 42524 57452 42576 57458
rect 42524 57394 42576 57400
rect 44088 57452 44140 57458
rect 44088 57394 44140 57400
rect 44180 57452 44232 57458
rect 44180 57394 44232 57400
rect 47584 57452 47636 57458
rect 47584 57394 47636 57400
rect 48688 57452 48740 57458
rect 48688 57394 48740 57400
rect 50160 57452 50212 57458
rect 50160 57394 50212 57400
rect 51816 57452 51868 57458
rect 51816 57394 51868 57400
rect 53380 57452 53432 57458
rect 53380 57394 53432 57400
rect 32232 56506 32260 57394
rect 33244 56506 33272 57394
rect 37188 57316 37240 57322
rect 37188 57258 37240 57264
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 37200 56506 37228 57258
rect 40788 56710 40816 57394
rect 42536 56778 42564 57394
rect 42524 56772 42576 56778
rect 42524 56714 42576 56720
rect 40776 56704 40828 56710
rect 40776 56646 40828 56652
rect 32220 56500 32272 56506
rect 32220 56442 32272 56448
rect 33232 56500 33284 56506
rect 33232 56442 33284 56448
rect 37188 56500 37240 56506
rect 37188 56442 37240 56448
rect 30932 56364 30984 56370
rect 30932 56306 30984 56312
rect 32128 56364 32180 56370
rect 32128 56306 32180 56312
rect 35716 56364 35768 56370
rect 35716 56306 35768 56312
rect 30380 56160 30432 56166
rect 30380 56102 30432 56108
rect 30944 55622 30972 56306
rect 29184 55616 29236 55622
rect 29184 55558 29236 55564
rect 30932 55616 30984 55622
rect 30932 55558 30984 55564
rect 29196 47569 29224 55558
rect 30944 50289 30972 55558
rect 32140 53145 32168 56306
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 32126 53136 32182 53145
rect 32126 53071 32182 53080
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 30930 50280 30986 50289
rect 30930 50215 30986 50224
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 29182 47560 29238 47569
rect 29182 47495 29238 47504
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 27986 44840 28042 44849
rect 27986 44775 28042 44784
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 26056 41676 26108 41682
rect 26056 41618 26108 41624
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 27344 40520 27396 40526
rect 27344 40462 27396 40468
rect 31208 40520 31260 40526
rect 31208 40462 31260 40468
rect 27068 40044 27120 40050
rect 27068 39986 27120 39992
rect 27080 39846 27108 39986
rect 27068 39840 27120 39846
rect 27068 39782 27120 39788
rect 26976 38956 27028 38962
rect 26976 38898 27028 38904
rect 26792 38752 26844 38758
rect 26792 38694 26844 38700
rect 25504 38548 25556 38554
rect 25504 38490 25556 38496
rect 25228 36644 25280 36650
rect 25228 36586 25280 36592
rect 25240 35698 25268 36586
rect 25516 35894 25544 38490
rect 25964 38208 26016 38214
rect 25964 38150 26016 38156
rect 25976 37942 26004 38150
rect 25964 37936 26016 37942
rect 25964 37878 26016 37884
rect 26240 36100 26292 36106
rect 26240 36042 26292 36048
rect 25516 35866 25636 35894
rect 25228 35692 25280 35698
rect 25280 35652 25360 35680
rect 25228 35634 25280 35640
rect 25228 33856 25280 33862
rect 25228 33798 25280 33804
rect 25240 33522 25268 33798
rect 25228 33516 25280 33522
rect 25228 33458 25280 33464
rect 25332 31482 25360 35652
rect 25320 31476 25372 31482
rect 25320 31418 25372 31424
rect 25504 31340 25556 31346
rect 25424 31300 25504 31328
rect 25320 30592 25372 30598
rect 25320 30534 25372 30540
rect 25332 30258 25360 30534
rect 25320 30252 25372 30258
rect 25320 30194 25372 30200
rect 25320 30116 25372 30122
rect 25320 30058 25372 30064
rect 25332 29714 25360 30058
rect 25320 29708 25372 29714
rect 25320 29650 25372 29656
rect 25228 29300 25280 29306
rect 25228 29242 25280 29248
rect 25240 26518 25268 29242
rect 25332 27538 25360 29650
rect 25424 29170 25452 31300
rect 25504 31282 25556 31288
rect 25504 30252 25556 30258
rect 25504 30194 25556 30200
rect 25516 29850 25544 30194
rect 25504 29844 25556 29850
rect 25504 29786 25556 29792
rect 25608 29306 25636 35866
rect 26252 35834 26280 36042
rect 26240 35828 26292 35834
rect 26240 35770 26292 35776
rect 25872 35488 25924 35494
rect 25872 35430 25924 35436
rect 25884 34746 25912 35430
rect 25964 35216 26016 35222
rect 25964 35158 26016 35164
rect 25872 34740 25924 34746
rect 25872 34682 25924 34688
rect 25884 34202 25912 34682
rect 25872 34196 25924 34202
rect 25872 34138 25924 34144
rect 25884 33522 25912 34138
rect 25872 33516 25924 33522
rect 25872 33458 25924 33464
rect 25884 29306 25912 33458
rect 25976 31482 26004 35158
rect 26240 33312 26292 33318
rect 26240 33254 26292 33260
rect 26252 33114 26280 33254
rect 26240 33108 26292 33114
rect 26240 33050 26292 33056
rect 26700 32224 26752 32230
rect 26700 32166 26752 32172
rect 26056 31680 26108 31686
rect 26056 31622 26108 31628
rect 25964 31476 26016 31482
rect 25964 31418 26016 31424
rect 26068 31346 26096 31622
rect 26056 31340 26108 31346
rect 26056 31282 26108 31288
rect 26240 30660 26292 30666
rect 26240 30602 26292 30608
rect 26252 30326 26280 30602
rect 26240 30320 26292 30326
rect 26240 30262 26292 30268
rect 25596 29300 25648 29306
rect 25596 29242 25648 29248
rect 25872 29300 25924 29306
rect 25872 29242 25924 29248
rect 26146 29200 26202 29209
rect 25412 29164 25464 29170
rect 26146 29135 26148 29144
rect 25412 29106 25464 29112
rect 26200 29135 26202 29144
rect 26148 29106 26200 29112
rect 25424 28490 25452 29106
rect 25412 28484 25464 28490
rect 25412 28426 25464 28432
rect 25504 27872 25556 27878
rect 25504 27814 25556 27820
rect 25320 27532 25372 27538
rect 25320 27474 25372 27480
rect 25412 27396 25464 27402
rect 25412 27338 25464 27344
rect 25424 27130 25452 27338
rect 25412 27124 25464 27130
rect 25412 27066 25464 27072
rect 25320 26988 25372 26994
rect 25320 26930 25372 26936
rect 25332 26790 25360 26930
rect 25320 26784 25372 26790
rect 25320 26726 25372 26732
rect 25228 26512 25280 26518
rect 25228 26454 25280 26460
rect 25240 26382 25268 26454
rect 25228 26376 25280 26382
rect 25228 26318 25280 26324
rect 25240 26042 25268 26318
rect 25228 26036 25280 26042
rect 25228 25978 25280 25984
rect 25228 25424 25280 25430
rect 25228 25366 25280 25372
rect 25240 13326 25268 25366
rect 25412 24200 25464 24206
rect 25412 24142 25464 24148
rect 25320 24064 25372 24070
rect 25320 24006 25372 24012
rect 25332 23730 25360 24006
rect 25424 23769 25452 24142
rect 25410 23760 25466 23769
rect 25320 23724 25372 23730
rect 25410 23695 25466 23704
rect 25320 23666 25372 23672
rect 25320 23044 25372 23050
rect 25320 22986 25372 22992
rect 25332 17066 25360 22986
rect 25516 18630 25544 27814
rect 25596 26852 25648 26858
rect 25596 26794 25648 26800
rect 25608 26450 25636 26794
rect 25688 26784 25740 26790
rect 25688 26726 25740 26732
rect 25596 26444 25648 26450
rect 25596 26386 25648 26392
rect 25700 26234 25728 26726
rect 25700 26206 25820 26234
rect 25792 25906 25820 26206
rect 25780 25900 25832 25906
rect 25780 25842 25832 25848
rect 25872 25900 25924 25906
rect 25872 25842 25924 25848
rect 25884 24274 25912 25842
rect 25964 25220 26016 25226
rect 25964 25162 26016 25168
rect 25872 24268 25924 24274
rect 25872 24210 25924 24216
rect 25872 24064 25924 24070
rect 25976 24052 26004 25162
rect 26056 24676 26108 24682
rect 26056 24618 26108 24624
rect 26068 24206 26096 24618
rect 26240 24608 26292 24614
rect 26240 24550 26292 24556
rect 26252 24342 26280 24550
rect 26240 24336 26292 24342
rect 26240 24278 26292 24284
rect 26056 24200 26108 24206
rect 26056 24142 26108 24148
rect 26240 24200 26292 24206
rect 26240 24142 26292 24148
rect 25976 24024 26096 24052
rect 25872 24006 25924 24012
rect 25596 23792 25648 23798
rect 25596 23734 25648 23740
rect 25608 23118 25636 23734
rect 25884 23118 25912 24006
rect 26068 23526 26096 24024
rect 26056 23520 26108 23526
rect 26056 23462 26108 23468
rect 25596 23112 25648 23118
rect 25596 23054 25648 23060
rect 25872 23112 25924 23118
rect 25872 23054 25924 23060
rect 25608 22574 25636 23054
rect 25964 22636 26016 22642
rect 26068 22624 26096 23462
rect 26252 22778 26280 24142
rect 26240 22772 26292 22778
rect 26240 22714 26292 22720
rect 26016 22596 26096 22624
rect 25964 22578 26016 22584
rect 25596 22568 25648 22574
rect 25596 22510 25648 22516
rect 25608 22094 25636 22510
rect 25608 22066 25728 22094
rect 25700 21350 25728 22066
rect 25976 21894 26004 22578
rect 25964 21888 26016 21894
rect 25964 21830 26016 21836
rect 25688 21344 25740 21350
rect 25688 21286 25740 21292
rect 25964 21344 26016 21350
rect 25964 21286 26016 21292
rect 25700 19854 25728 21286
rect 25780 20936 25832 20942
rect 25780 20878 25832 20884
rect 25792 20058 25820 20878
rect 25872 20256 25924 20262
rect 25872 20198 25924 20204
rect 25780 20052 25832 20058
rect 25780 19994 25832 20000
rect 25884 19854 25912 20198
rect 25688 19848 25740 19854
rect 25872 19848 25924 19854
rect 25740 19796 25820 19802
rect 25688 19790 25820 19796
rect 25872 19790 25924 19796
rect 25700 19774 25820 19790
rect 25688 19372 25740 19378
rect 25688 19314 25740 19320
rect 25504 18624 25556 18630
rect 25504 18566 25556 18572
rect 25700 17882 25728 19314
rect 25792 18290 25820 19774
rect 25872 19712 25924 19718
rect 25872 19654 25924 19660
rect 25884 19446 25912 19654
rect 25872 19440 25924 19446
rect 25872 19382 25924 19388
rect 25780 18284 25832 18290
rect 25780 18226 25832 18232
rect 25688 17876 25740 17882
rect 25688 17818 25740 17824
rect 25412 17672 25464 17678
rect 25412 17614 25464 17620
rect 25320 17060 25372 17066
rect 25320 17002 25372 17008
rect 25424 14414 25452 17614
rect 25688 17604 25740 17610
rect 25688 17546 25740 17552
rect 25504 17536 25556 17542
rect 25504 17478 25556 17484
rect 25516 17338 25544 17478
rect 25700 17338 25728 17546
rect 25504 17332 25556 17338
rect 25504 17274 25556 17280
rect 25688 17332 25740 17338
rect 25688 17274 25740 17280
rect 25504 16992 25556 16998
rect 25504 16934 25556 16940
rect 25516 16590 25544 16934
rect 25504 16584 25556 16590
rect 25504 16526 25556 16532
rect 25516 16250 25544 16526
rect 25504 16244 25556 16250
rect 25504 16186 25556 16192
rect 25412 14408 25464 14414
rect 25412 14350 25464 14356
rect 25424 14074 25452 14350
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 25228 13320 25280 13326
rect 25228 13262 25280 13268
rect 25240 12986 25268 13262
rect 25228 12980 25280 12986
rect 25228 12922 25280 12928
rect 25424 12238 25452 14010
rect 25976 13938 26004 21286
rect 26712 21010 26740 32166
rect 26804 28762 26832 38694
rect 26884 33380 26936 33386
rect 26884 33322 26936 33328
rect 26896 32910 26924 33322
rect 26988 33318 27016 38898
rect 27080 38894 27108 39782
rect 27356 39438 27384 40462
rect 27620 40452 27672 40458
rect 27620 40394 27672 40400
rect 27632 40186 27660 40394
rect 28724 40384 28776 40390
rect 28724 40326 28776 40332
rect 27620 40180 27672 40186
rect 27620 40122 27672 40128
rect 28736 40118 28764 40326
rect 28724 40112 28776 40118
rect 28724 40054 28776 40060
rect 29092 40112 29144 40118
rect 29092 40054 29144 40060
rect 27988 40044 28040 40050
rect 27988 39986 28040 39992
rect 28264 40044 28316 40050
rect 28264 39986 28316 39992
rect 27344 39432 27396 39438
rect 27396 39380 27476 39386
rect 27344 39374 27476 39380
rect 27356 39358 27476 39374
rect 27068 38888 27120 38894
rect 27068 38830 27120 38836
rect 27080 36378 27108 38830
rect 27448 37670 27476 39358
rect 27528 39364 27580 39370
rect 27528 39306 27580 39312
rect 27540 39098 27568 39306
rect 28000 39098 28028 39986
rect 28276 39438 28304 39986
rect 28264 39432 28316 39438
rect 28264 39374 28316 39380
rect 27528 39092 27580 39098
rect 27528 39034 27580 39040
rect 27988 39092 28040 39098
rect 27988 39034 28040 39040
rect 28276 38962 28304 39374
rect 28632 39296 28684 39302
rect 28632 39238 28684 39244
rect 28264 38956 28316 38962
rect 28264 38898 28316 38904
rect 28080 38888 28132 38894
rect 28080 38830 28132 38836
rect 28092 38554 28120 38830
rect 28080 38548 28132 38554
rect 28080 38490 28132 38496
rect 28644 38350 28672 39238
rect 28632 38344 28684 38350
rect 28632 38286 28684 38292
rect 27436 37664 27488 37670
rect 27436 37606 27488 37612
rect 27448 36786 27476 37606
rect 28172 37120 28224 37126
rect 28172 37062 28224 37068
rect 27436 36780 27488 36786
rect 27436 36722 27488 36728
rect 27528 36780 27580 36786
rect 27528 36722 27580 36728
rect 27988 36780 28040 36786
rect 27988 36722 28040 36728
rect 27068 36372 27120 36378
rect 27068 36314 27120 36320
rect 27080 36174 27108 36314
rect 27448 36242 27476 36722
rect 27540 36378 27568 36722
rect 27528 36372 27580 36378
rect 27528 36314 27580 36320
rect 27436 36236 27488 36242
rect 27436 36178 27488 36184
rect 27068 36168 27120 36174
rect 27068 36110 27120 36116
rect 28000 35766 28028 36722
rect 28184 36174 28212 37062
rect 28448 36576 28500 36582
rect 28448 36518 28500 36524
rect 28172 36168 28224 36174
rect 28172 36110 28224 36116
rect 27988 35760 28040 35766
rect 27988 35702 28040 35708
rect 28184 35562 28212 36110
rect 28460 36106 28488 36518
rect 28448 36100 28500 36106
rect 28448 36042 28500 36048
rect 28264 35828 28316 35834
rect 28264 35770 28316 35776
rect 28172 35556 28224 35562
rect 28172 35498 28224 35504
rect 27712 34400 27764 34406
rect 27712 34342 27764 34348
rect 27068 33992 27120 33998
rect 27068 33934 27120 33940
rect 26976 33312 27028 33318
rect 26976 33254 27028 33260
rect 27080 32910 27108 33934
rect 27252 33924 27304 33930
rect 27252 33866 27304 33872
rect 27264 33658 27292 33866
rect 27252 33652 27304 33658
rect 27252 33594 27304 33600
rect 27724 33522 27752 34342
rect 28184 33522 28212 35498
rect 28276 34542 28304 35770
rect 28356 34672 28408 34678
rect 28356 34614 28408 34620
rect 28264 34536 28316 34542
rect 28264 34478 28316 34484
rect 27712 33516 27764 33522
rect 27712 33458 27764 33464
rect 28172 33516 28224 33522
rect 28172 33458 28224 33464
rect 28184 33114 28212 33458
rect 28172 33108 28224 33114
rect 28172 33050 28224 33056
rect 26884 32904 26936 32910
rect 26884 32846 26936 32852
rect 27068 32904 27120 32910
rect 27068 32846 27120 32852
rect 27252 32904 27304 32910
rect 27252 32846 27304 32852
rect 27264 32026 27292 32846
rect 28172 32360 28224 32366
rect 28172 32302 28224 32308
rect 27252 32020 27304 32026
rect 27252 31962 27304 31968
rect 27264 30802 27292 31962
rect 27896 31952 27948 31958
rect 27896 31894 27948 31900
rect 27252 30796 27304 30802
rect 27252 30738 27304 30744
rect 27264 29646 27292 30738
rect 27804 30048 27856 30054
rect 27804 29990 27856 29996
rect 27816 29850 27844 29990
rect 27804 29844 27856 29850
rect 27804 29786 27856 29792
rect 27816 29646 27844 29786
rect 27252 29640 27304 29646
rect 27252 29582 27304 29588
rect 27804 29640 27856 29646
rect 27804 29582 27856 29588
rect 26792 28756 26844 28762
rect 26792 28698 26844 28704
rect 26804 27614 26832 28698
rect 27160 28484 27212 28490
rect 27160 28426 27212 28432
rect 26804 27586 26924 27614
rect 26792 26784 26844 26790
rect 26792 26726 26844 26732
rect 26700 21004 26752 21010
rect 26700 20946 26752 20952
rect 26240 20800 26292 20806
rect 26240 20742 26292 20748
rect 26252 20466 26280 20742
rect 26240 20460 26292 20466
rect 26240 20402 26292 20408
rect 26424 20460 26476 20466
rect 26424 20402 26476 20408
rect 26148 20256 26200 20262
rect 26148 20198 26200 20204
rect 26160 19378 26188 20198
rect 26436 19718 26464 20402
rect 26424 19712 26476 19718
rect 26424 19654 26476 19660
rect 26700 19508 26752 19514
rect 26700 19450 26752 19456
rect 26148 19372 26200 19378
rect 26148 19314 26200 19320
rect 26424 19372 26476 19378
rect 26424 19314 26476 19320
rect 26240 18216 26292 18222
rect 26240 18158 26292 18164
rect 26148 17536 26200 17542
rect 26148 17478 26200 17484
rect 26160 17202 26188 17478
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 26148 17060 26200 17066
rect 26148 17002 26200 17008
rect 26160 16590 26188 17002
rect 26148 16584 26200 16590
rect 26148 16526 26200 16532
rect 26252 16522 26280 18158
rect 26332 16584 26384 16590
rect 26332 16526 26384 16532
rect 26240 16516 26292 16522
rect 26240 16458 26292 16464
rect 26252 16182 26280 16458
rect 26344 16250 26372 16526
rect 26332 16244 26384 16250
rect 26332 16186 26384 16192
rect 26240 16176 26292 16182
rect 26240 16118 26292 16124
rect 25964 13932 26016 13938
rect 25964 13874 26016 13880
rect 25976 13530 26004 13874
rect 25964 13524 26016 13530
rect 25964 13466 26016 13472
rect 25412 12232 25464 12238
rect 25412 12174 25464 12180
rect 25596 12164 25648 12170
rect 25596 12106 25648 12112
rect 25608 11898 25636 12106
rect 25964 12096 26016 12102
rect 25964 12038 26016 12044
rect 25596 11892 25648 11898
rect 25596 11834 25648 11840
rect 25976 11150 26004 12038
rect 26148 11756 26200 11762
rect 26148 11698 26200 11704
rect 26160 11354 26188 11698
rect 26332 11688 26384 11694
rect 26332 11630 26384 11636
rect 26148 11348 26200 11354
rect 26148 11290 26200 11296
rect 26344 11218 26372 11630
rect 26332 11212 26384 11218
rect 26332 11154 26384 11160
rect 25964 11144 26016 11150
rect 25964 11086 26016 11092
rect 25780 11076 25832 11082
rect 25780 11018 25832 11024
rect 25792 10674 25820 11018
rect 25320 10668 25372 10674
rect 25320 10610 25372 10616
rect 25780 10668 25832 10674
rect 25780 10610 25832 10616
rect 25332 10266 25360 10610
rect 25320 10260 25372 10266
rect 25320 10202 25372 10208
rect 25792 9722 25820 10610
rect 25976 10062 26004 11086
rect 26332 10464 26384 10470
rect 26332 10406 26384 10412
rect 25964 10056 26016 10062
rect 25964 9998 26016 10004
rect 26240 10056 26292 10062
rect 26240 9998 26292 10004
rect 25780 9716 25832 9722
rect 25780 9658 25832 9664
rect 25780 9444 25832 9450
rect 25780 9386 25832 9392
rect 25320 7812 25372 7818
rect 25320 7754 25372 7760
rect 25332 7342 25360 7754
rect 25792 7585 25820 9386
rect 26252 9382 26280 9998
rect 26344 9926 26372 10406
rect 26436 10266 26464 19314
rect 26712 18970 26740 19450
rect 26700 18964 26752 18970
rect 26700 18906 26752 18912
rect 26804 18698 26832 26726
rect 26896 25974 26924 27586
rect 26976 26240 27028 26246
rect 26976 26182 27028 26188
rect 26884 25968 26936 25974
rect 26884 25910 26936 25916
rect 26988 25294 27016 26182
rect 26976 25288 27028 25294
rect 26976 25230 27028 25236
rect 26988 23118 27016 25230
rect 26976 23112 27028 23118
rect 26976 23054 27028 23060
rect 26976 22976 27028 22982
rect 26976 22918 27028 22924
rect 26988 22710 27016 22918
rect 26976 22704 27028 22710
rect 26976 22646 27028 22652
rect 26884 20460 26936 20466
rect 26884 20402 26936 20408
rect 26792 18692 26844 18698
rect 26792 18634 26844 18640
rect 26516 18624 26568 18630
rect 26516 18566 26568 18572
rect 26424 10260 26476 10266
rect 26424 10202 26476 10208
rect 26332 9920 26384 9926
rect 26332 9862 26384 9868
rect 26344 9654 26372 9862
rect 26332 9648 26384 9654
rect 26332 9590 26384 9596
rect 26240 9376 26292 9382
rect 26240 9318 26292 9324
rect 26252 9042 26280 9318
rect 26240 9036 26292 9042
rect 26240 8978 26292 8984
rect 25964 8016 26016 8022
rect 25964 7958 26016 7964
rect 25778 7576 25834 7585
rect 25778 7511 25834 7520
rect 25792 7410 25820 7511
rect 25976 7410 26004 7958
rect 25780 7404 25832 7410
rect 25780 7346 25832 7352
rect 25964 7404 26016 7410
rect 25964 7346 26016 7352
rect 25320 7336 25372 7342
rect 25320 7278 25372 7284
rect 25792 5710 25820 7346
rect 26240 7336 26292 7342
rect 26240 7278 26292 7284
rect 26252 6798 26280 7278
rect 26240 6792 26292 6798
rect 26240 6734 26292 6740
rect 26148 6384 26200 6390
rect 26148 6326 26200 6332
rect 26160 5914 26188 6326
rect 26148 5908 26200 5914
rect 26148 5850 26200 5856
rect 25320 5704 25372 5710
rect 25320 5646 25372 5652
rect 25780 5704 25832 5710
rect 25780 5646 25832 5652
rect 25332 5234 25360 5646
rect 26252 5302 26280 6734
rect 26240 5296 26292 5302
rect 26240 5238 26292 5244
rect 26528 5234 26556 18566
rect 26700 17332 26752 17338
rect 26700 17274 26752 17280
rect 26608 17264 26660 17270
rect 26606 17232 26608 17241
rect 26660 17232 26662 17241
rect 26606 17167 26662 17176
rect 26712 16658 26740 17274
rect 26792 17196 26844 17202
rect 26792 17138 26844 17144
rect 26804 16794 26832 17138
rect 26792 16788 26844 16794
rect 26792 16730 26844 16736
rect 26700 16652 26752 16658
rect 26700 16594 26752 16600
rect 26608 16584 26660 16590
rect 26608 16526 26660 16532
rect 26620 16250 26648 16526
rect 26608 16244 26660 16250
rect 26608 16186 26660 16192
rect 26620 16114 26648 16186
rect 26608 16108 26660 16114
rect 26608 16050 26660 16056
rect 26712 15706 26740 16594
rect 26700 15700 26752 15706
rect 26700 15642 26752 15648
rect 26896 7750 26924 20402
rect 26988 19922 27016 22646
rect 27068 21004 27120 21010
rect 27068 20946 27120 20952
rect 26976 19916 27028 19922
rect 26976 19858 27028 19864
rect 26974 19816 27030 19825
rect 26974 19751 27030 19760
rect 26988 19514 27016 19751
rect 26976 19508 27028 19514
rect 26976 19450 27028 19456
rect 26976 18284 27028 18290
rect 26976 18226 27028 18232
rect 26988 17134 27016 18226
rect 26976 17128 27028 17134
rect 26976 17070 27028 17076
rect 27080 15638 27108 20946
rect 27172 19496 27200 28426
rect 27264 27470 27292 29582
rect 27344 29164 27396 29170
rect 27344 29106 27396 29112
rect 27252 27464 27304 27470
rect 27252 27406 27304 27412
rect 27356 22094 27384 29106
rect 27436 26988 27488 26994
rect 27436 26930 27488 26936
rect 27448 26314 27476 26930
rect 27436 26308 27488 26314
rect 27436 26250 27488 26256
rect 27448 25226 27476 26250
rect 27436 25220 27488 25226
rect 27436 25162 27488 25168
rect 27528 24948 27580 24954
rect 27528 24890 27580 24896
rect 27264 22066 27384 22094
rect 27264 20806 27292 22066
rect 27252 20800 27304 20806
rect 27252 20742 27304 20748
rect 27264 20466 27292 20742
rect 27436 20528 27488 20534
rect 27436 20470 27488 20476
rect 27252 20460 27304 20466
rect 27252 20402 27304 20408
rect 27172 19468 27292 19496
rect 27160 19372 27212 19378
rect 27160 19314 27212 19320
rect 27172 18154 27200 19314
rect 27160 18148 27212 18154
rect 27160 18090 27212 18096
rect 27264 17338 27292 19468
rect 27344 19168 27396 19174
rect 27344 19110 27396 19116
rect 27356 18970 27384 19110
rect 27344 18964 27396 18970
rect 27344 18906 27396 18912
rect 27448 18630 27476 20470
rect 27540 19446 27568 24890
rect 27620 23792 27672 23798
rect 27620 23734 27672 23740
rect 27632 22778 27660 23734
rect 27620 22772 27672 22778
rect 27620 22714 27672 22720
rect 27908 22094 27936 31894
rect 28184 31822 28212 32302
rect 28276 32065 28304 34478
rect 28368 33862 28396 34614
rect 28356 33856 28408 33862
rect 28356 33798 28408 33804
rect 28262 32056 28318 32065
rect 28262 31991 28318 32000
rect 28368 31822 28396 33798
rect 28460 32502 28488 36042
rect 28448 32496 28500 32502
rect 28448 32438 28500 32444
rect 28540 32428 28592 32434
rect 28540 32370 28592 32376
rect 28552 32178 28580 32370
rect 28460 32150 28580 32178
rect 28460 32026 28488 32150
rect 28538 32056 28594 32065
rect 28448 32020 28500 32026
rect 28538 31991 28594 32000
rect 28448 31962 28500 31968
rect 28172 31816 28224 31822
rect 28172 31758 28224 31764
rect 28356 31816 28408 31822
rect 28356 31758 28408 31764
rect 28460 31754 28488 31962
rect 28448 31748 28500 31754
rect 28448 31690 28500 31696
rect 28552 31414 28580 31991
rect 28644 31822 28672 38286
rect 28736 32434 28764 40054
rect 28816 38752 28868 38758
rect 28816 38694 28868 38700
rect 28828 37874 28856 38694
rect 29104 38282 29132 40054
rect 30288 39432 30340 39438
rect 30288 39374 30340 39380
rect 31116 39432 31168 39438
rect 31116 39374 31168 39380
rect 30196 38344 30248 38350
rect 30196 38286 30248 38292
rect 29092 38276 29144 38282
rect 29092 38218 29144 38224
rect 29552 38208 29604 38214
rect 29552 38150 29604 38156
rect 28816 37868 28868 37874
rect 28816 37810 28868 37816
rect 28828 36854 28856 37810
rect 28908 37664 28960 37670
rect 28908 37606 28960 37612
rect 28816 36848 28868 36854
rect 28816 36790 28868 36796
rect 28828 36310 28856 36790
rect 28816 36304 28868 36310
rect 28816 36246 28868 36252
rect 28724 32428 28776 32434
rect 28724 32370 28776 32376
rect 28724 32292 28776 32298
rect 28724 32234 28776 32240
rect 28632 31816 28684 31822
rect 28632 31758 28684 31764
rect 28540 31408 28592 31414
rect 28540 31350 28592 31356
rect 28080 31340 28132 31346
rect 28080 31282 28132 31288
rect 28092 31142 28120 31282
rect 28540 31272 28592 31278
rect 28540 31214 28592 31220
rect 28080 31136 28132 31142
rect 28080 31078 28132 31084
rect 27988 26988 28040 26994
rect 27988 26930 28040 26936
rect 28000 26042 28028 26930
rect 27988 26036 28040 26042
rect 27988 25978 28040 25984
rect 27988 22636 28040 22642
rect 27988 22578 28040 22584
rect 27816 22066 27936 22094
rect 27620 21548 27672 21554
rect 27620 21490 27672 21496
rect 27632 21350 27660 21490
rect 27712 21480 27764 21486
rect 27712 21422 27764 21428
rect 27620 21344 27672 21350
rect 27620 21286 27672 21292
rect 27632 20330 27660 21286
rect 27620 20324 27672 20330
rect 27620 20266 27672 20272
rect 27724 20210 27752 21422
rect 27632 20182 27752 20210
rect 27632 19718 27660 20182
rect 27620 19712 27672 19718
rect 27620 19654 27672 19660
rect 27528 19440 27580 19446
rect 27528 19382 27580 19388
rect 27632 18902 27660 19654
rect 27620 18896 27672 18902
rect 27620 18838 27672 18844
rect 27436 18624 27488 18630
rect 27436 18566 27488 18572
rect 27436 17604 27488 17610
rect 27436 17546 27488 17552
rect 27252 17332 27304 17338
rect 27252 17274 27304 17280
rect 27448 16794 27476 17546
rect 27436 16788 27488 16794
rect 27436 16730 27488 16736
rect 27252 16652 27304 16658
rect 27252 16594 27304 16600
rect 27264 15910 27292 16594
rect 27448 16182 27476 16730
rect 27528 16584 27580 16590
rect 27528 16526 27580 16532
rect 27436 16176 27488 16182
rect 27436 16118 27488 16124
rect 27540 16046 27568 16526
rect 27528 16040 27580 16046
rect 27528 15982 27580 15988
rect 27252 15904 27304 15910
rect 27252 15846 27304 15852
rect 27068 15632 27120 15638
rect 27068 15574 27120 15580
rect 27068 15496 27120 15502
rect 27068 15438 27120 15444
rect 27080 14958 27108 15438
rect 27264 15065 27292 15846
rect 27540 15502 27568 15982
rect 27528 15496 27580 15502
rect 27528 15438 27580 15444
rect 27250 15056 27306 15065
rect 27250 14991 27306 15000
rect 27068 14952 27120 14958
rect 27068 14894 27120 14900
rect 27344 14816 27396 14822
rect 27344 14758 27396 14764
rect 27712 14816 27764 14822
rect 27712 14758 27764 14764
rect 26976 14340 27028 14346
rect 26976 14282 27028 14288
rect 27160 14340 27212 14346
rect 27160 14282 27212 14288
rect 26988 13462 27016 14282
rect 27172 14074 27200 14282
rect 27160 14068 27212 14074
rect 27160 14010 27212 14016
rect 27068 13932 27120 13938
rect 27068 13874 27120 13880
rect 26976 13456 27028 13462
rect 26976 13398 27028 13404
rect 27080 12646 27108 13874
rect 27356 13308 27384 14758
rect 27528 13932 27580 13938
rect 27528 13874 27580 13880
rect 27540 13462 27568 13874
rect 27528 13456 27580 13462
rect 27528 13398 27580 13404
rect 27436 13320 27488 13326
rect 27356 13280 27436 13308
rect 27436 13262 27488 13268
rect 27068 12640 27120 12646
rect 27068 12582 27120 12588
rect 27080 9382 27108 12582
rect 27724 12102 27752 14758
rect 27816 13734 27844 22066
rect 28000 21690 28028 22578
rect 28092 22166 28120 31078
rect 28172 25696 28224 25702
rect 28172 25638 28224 25644
rect 28184 24886 28212 25638
rect 28264 25220 28316 25226
rect 28264 25162 28316 25168
rect 28172 24880 28224 24886
rect 28172 24822 28224 24828
rect 28184 24410 28212 24822
rect 28276 24818 28304 25162
rect 28264 24812 28316 24818
rect 28264 24754 28316 24760
rect 28172 24404 28224 24410
rect 28172 24346 28224 24352
rect 28276 23730 28304 24754
rect 28356 24676 28408 24682
rect 28356 24618 28408 24624
rect 28368 24138 28396 24618
rect 28356 24132 28408 24138
rect 28356 24074 28408 24080
rect 28448 24132 28500 24138
rect 28448 24074 28500 24080
rect 28264 23724 28316 23730
rect 28264 23666 28316 23672
rect 28172 22976 28224 22982
rect 28172 22918 28224 22924
rect 28080 22160 28132 22166
rect 28080 22102 28132 22108
rect 27988 21684 28040 21690
rect 27988 21626 28040 21632
rect 27988 18692 28040 18698
rect 27988 18634 28040 18640
rect 27896 15904 27948 15910
rect 27896 15846 27948 15852
rect 27804 13728 27856 13734
rect 27804 13670 27856 13676
rect 27804 13320 27856 13326
rect 27804 13262 27856 13268
rect 27816 12986 27844 13262
rect 27804 12980 27856 12986
rect 27804 12922 27856 12928
rect 27528 12096 27580 12102
rect 27528 12038 27580 12044
rect 27712 12096 27764 12102
rect 27712 12038 27764 12044
rect 27540 11762 27568 12038
rect 27528 11756 27580 11762
rect 27528 11698 27580 11704
rect 27160 10804 27212 10810
rect 27160 10746 27212 10752
rect 27068 9376 27120 9382
rect 27068 9318 27120 9324
rect 27080 9178 27108 9318
rect 27068 9172 27120 9178
rect 27068 9114 27120 9120
rect 27172 8090 27200 10746
rect 27724 10198 27752 12038
rect 27712 10192 27764 10198
rect 27712 10134 27764 10140
rect 27436 10056 27488 10062
rect 27436 9998 27488 10004
rect 27804 10056 27856 10062
rect 27804 9998 27856 10004
rect 27160 8084 27212 8090
rect 27160 8026 27212 8032
rect 26884 7744 26936 7750
rect 26884 7686 26936 7692
rect 26896 7410 26924 7686
rect 26884 7404 26936 7410
rect 26884 7346 26936 7352
rect 27344 7200 27396 7206
rect 27344 7142 27396 7148
rect 27160 6792 27212 6798
rect 27160 6734 27212 6740
rect 26884 6248 26936 6254
rect 26884 6190 26936 6196
rect 26896 5914 26924 6190
rect 26884 5908 26936 5914
rect 26884 5850 26936 5856
rect 25320 5228 25372 5234
rect 25320 5170 25372 5176
rect 26332 5228 26384 5234
rect 26332 5170 26384 5176
rect 26516 5228 26568 5234
rect 26516 5170 26568 5176
rect 26344 5030 26372 5170
rect 26332 5024 26384 5030
rect 26332 4966 26384 4972
rect 25688 3936 25740 3942
rect 25688 3878 25740 3884
rect 26240 3936 26292 3942
rect 26240 3878 26292 3884
rect 25700 3738 25728 3878
rect 25688 3732 25740 3738
rect 25688 3674 25740 3680
rect 26252 3670 26280 3878
rect 26240 3664 26292 3670
rect 26240 3606 26292 3612
rect 25596 3528 25648 3534
rect 25596 3470 25648 3476
rect 25320 2848 25372 2854
rect 25320 2790 25372 2796
rect 25136 2100 25188 2106
rect 25136 2042 25188 2048
rect 25332 800 25360 2790
rect 25608 800 25636 3470
rect 26344 2961 26372 4966
rect 27172 4690 27200 6734
rect 27356 6730 27384 7142
rect 27344 6724 27396 6730
rect 27344 6666 27396 6672
rect 27448 5778 27476 9998
rect 27528 9988 27580 9994
rect 27528 9930 27580 9936
rect 27540 9874 27568 9930
rect 27540 9846 27660 9874
rect 27632 8498 27660 9846
rect 27816 9110 27844 9998
rect 27804 9104 27856 9110
rect 27804 9046 27856 9052
rect 27620 8492 27672 8498
rect 27620 8434 27672 8440
rect 27620 8356 27672 8362
rect 27620 8298 27672 8304
rect 27632 7274 27660 8298
rect 27816 7886 27844 9046
rect 27908 8362 27936 15846
rect 28000 10266 28028 18634
rect 28080 13932 28132 13938
rect 28080 13874 28132 13880
rect 28092 13326 28120 13874
rect 28184 13569 28212 22918
rect 28276 21962 28304 23666
rect 28264 21956 28316 21962
rect 28264 21898 28316 21904
rect 28276 20874 28304 21898
rect 28460 21554 28488 24074
rect 28552 22094 28580 31214
rect 28632 29640 28684 29646
rect 28736 29628 28764 32234
rect 28828 31754 28856 36246
rect 28920 35018 28948 37606
rect 29276 37120 29328 37126
rect 29276 37062 29328 37068
rect 29288 36786 29316 37062
rect 29276 36780 29328 36786
rect 29276 36722 29328 36728
rect 29460 36780 29512 36786
rect 29460 36722 29512 36728
rect 29000 36712 29052 36718
rect 29000 36654 29052 36660
rect 29012 36038 29040 36654
rect 29472 36378 29500 36722
rect 29460 36372 29512 36378
rect 29460 36314 29512 36320
rect 29564 36122 29592 38150
rect 29644 37120 29696 37126
rect 29644 37062 29696 37068
rect 29656 36786 29684 37062
rect 29644 36780 29696 36786
rect 29644 36722 29696 36728
rect 29472 36106 29592 36122
rect 29460 36100 29592 36106
rect 29512 36094 29592 36100
rect 29460 36042 29512 36048
rect 29000 36032 29052 36038
rect 29000 35974 29052 35980
rect 28908 35012 28960 35018
rect 28908 34954 28960 34960
rect 29012 34474 29040 35974
rect 29276 35080 29328 35086
rect 29276 35022 29328 35028
rect 29000 34468 29052 34474
rect 29000 34410 29052 34416
rect 28828 31726 28948 31754
rect 28920 31142 28948 31726
rect 28908 31136 28960 31142
rect 28908 31078 28960 31084
rect 28920 30598 28948 31078
rect 28908 30592 28960 30598
rect 28908 30534 28960 30540
rect 29288 30326 29316 35022
rect 29368 32360 29420 32366
rect 29368 32302 29420 32308
rect 29276 30320 29328 30326
rect 29276 30262 29328 30268
rect 28816 30048 28868 30054
rect 28816 29990 28868 29996
rect 28828 29646 28856 29990
rect 28684 29600 28764 29628
rect 28816 29640 28868 29646
rect 28632 29582 28684 29588
rect 28816 29582 28868 29588
rect 29380 29170 29408 32302
rect 29472 29238 29500 36042
rect 29552 34944 29604 34950
rect 29552 34886 29604 34892
rect 29564 34610 29592 34886
rect 29552 34604 29604 34610
rect 29552 34546 29604 34552
rect 29552 33516 29604 33522
rect 29552 33458 29604 33464
rect 29564 33318 29592 33458
rect 29552 33312 29604 33318
rect 29552 33254 29604 33260
rect 29564 32570 29592 33254
rect 29552 32564 29604 32570
rect 29552 32506 29604 32512
rect 29656 32298 29684 36722
rect 30208 35086 30236 38286
rect 30300 37874 30328 39374
rect 30564 39296 30616 39302
rect 30564 39238 30616 39244
rect 30380 38276 30432 38282
rect 30380 38218 30432 38224
rect 30288 37868 30340 37874
rect 30288 37810 30340 37816
rect 30300 36786 30328 37810
rect 30392 36922 30420 38218
rect 30472 38208 30524 38214
rect 30472 38150 30524 38156
rect 30484 37874 30512 38150
rect 30472 37868 30524 37874
rect 30472 37810 30524 37816
rect 30380 36916 30432 36922
rect 30380 36858 30432 36864
rect 30288 36780 30340 36786
rect 30288 36722 30340 36728
rect 30472 36100 30524 36106
rect 30472 36042 30524 36048
rect 30380 36032 30432 36038
rect 30380 35974 30432 35980
rect 30196 35080 30248 35086
rect 30196 35022 30248 35028
rect 29828 35012 29880 35018
rect 29828 34954 29880 34960
rect 29736 34604 29788 34610
rect 29736 34546 29788 34552
rect 29748 34066 29776 34546
rect 29840 34542 29868 34954
rect 29828 34536 29880 34542
rect 29828 34478 29880 34484
rect 30196 34400 30248 34406
rect 30248 34348 30328 34354
rect 30196 34342 30328 34348
rect 30208 34326 30328 34342
rect 29736 34060 29788 34066
rect 29736 34002 29788 34008
rect 29920 33992 29972 33998
rect 29920 33934 29972 33940
rect 29932 32910 29960 33934
rect 30300 33454 30328 34326
rect 30392 33998 30420 35974
rect 30484 35018 30512 36042
rect 30576 35714 30604 39238
rect 31128 39030 31156 39374
rect 31116 39024 31168 39030
rect 31116 38966 31168 38972
rect 30656 37868 30708 37874
rect 30656 37810 30708 37816
rect 30668 35834 30696 37810
rect 31128 37806 31156 38966
rect 31220 38418 31248 40462
rect 31484 40452 31536 40458
rect 31484 40394 31536 40400
rect 31496 39642 31524 40394
rect 32036 40384 32088 40390
rect 32036 40326 32088 40332
rect 31484 39636 31536 39642
rect 31484 39578 31536 39584
rect 31300 39432 31352 39438
rect 31300 39374 31352 39380
rect 31312 39302 31340 39374
rect 32048 39370 32076 40326
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 31760 39364 31812 39370
rect 31760 39306 31812 39312
rect 32036 39364 32088 39370
rect 32036 39306 32088 39312
rect 31300 39296 31352 39302
rect 31300 39238 31352 39244
rect 31208 38412 31260 38418
rect 31208 38354 31260 38360
rect 31668 38412 31720 38418
rect 31668 38354 31720 38360
rect 31680 37806 31708 38354
rect 31772 38282 31800 39306
rect 31944 38344 31996 38350
rect 31944 38286 31996 38292
rect 31760 38276 31812 38282
rect 31760 38218 31812 38224
rect 31116 37800 31168 37806
rect 31116 37742 31168 37748
rect 31668 37800 31720 37806
rect 31668 37742 31720 37748
rect 30932 37664 30984 37670
rect 30932 37606 30984 37612
rect 30944 37194 30972 37606
rect 30932 37188 30984 37194
rect 30932 37130 30984 37136
rect 30656 35828 30708 35834
rect 30656 35770 30708 35776
rect 30576 35686 30696 35714
rect 30472 35012 30524 35018
rect 30472 34954 30524 34960
rect 30484 34762 30512 34954
rect 30484 34746 30604 34762
rect 30484 34740 30616 34746
rect 30484 34734 30564 34740
rect 30564 34682 30616 34688
rect 30380 33992 30432 33998
rect 30380 33934 30432 33940
rect 30564 33856 30616 33862
rect 30564 33798 30616 33804
rect 30576 33522 30604 33798
rect 30668 33658 30696 35686
rect 30748 34060 30800 34066
rect 30748 34002 30800 34008
rect 30656 33652 30708 33658
rect 30656 33594 30708 33600
rect 30760 33522 30788 34002
rect 30564 33516 30616 33522
rect 30564 33458 30616 33464
rect 30748 33516 30800 33522
rect 30800 33476 30972 33504
rect 30748 33458 30800 33464
rect 30288 33448 30340 33454
rect 30288 33390 30340 33396
rect 30104 33312 30156 33318
rect 30104 33254 30156 33260
rect 29920 32904 29972 32910
rect 29920 32846 29972 32852
rect 29736 32768 29788 32774
rect 29736 32710 29788 32716
rect 29644 32292 29696 32298
rect 29644 32234 29696 32240
rect 29552 30252 29604 30258
rect 29552 30194 29604 30200
rect 29564 29850 29592 30194
rect 29552 29844 29604 29850
rect 29552 29786 29604 29792
rect 29564 29306 29592 29786
rect 29552 29300 29604 29306
rect 29552 29242 29604 29248
rect 29460 29232 29512 29238
rect 29460 29174 29512 29180
rect 29368 29164 29420 29170
rect 29368 29106 29420 29112
rect 29184 29028 29236 29034
rect 29184 28970 29236 28976
rect 28908 28552 28960 28558
rect 28908 28494 28960 28500
rect 28920 26194 28948 28494
rect 29000 28416 29052 28422
rect 29000 28358 29052 28364
rect 29012 28218 29040 28358
rect 29000 28212 29052 28218
rect 29000 28154 29052 28160
rect 29000 27328 29052 27334
rect 29000 27270 29052 27276
rect 29012 26314 29040 27270
rect 29000 26308 29052 26314
rect 29000 26250 29052 26256
rect 28920 26166 29132 26194
rect 29000 25900 29052 25906
rect 29000 25842 29052 25848
rect 28908 24744 28960 24750
rect 28908 24686 28960 24692
rect 28816 24608 28868 24614
rect 28816 24550 28868 24556
rect 28828 24206 28856 24550
rect 28816 24200 28868 24206
rect 28816 24142 28868 24148
rect 28816 24064 28868 24070
rect 28816 24006 28868 24012
rect 28828 22982 28856 24006
rect 28920 23798 28948 24686
rect 29012 24410 29040 25842
rect 29104 25242 29132 26166
rect 29196 25430 29224 28970
rect 29380 28558 29408 29106
rect 29368 28552 29420 28558
rect 29368 28494 29420 28500
rect 29380 28082 29408 28494
rect 29368 28076 29420 28082
rect 29368 28018 29420 28024
rect 29276 27872 29328 27878
rect 29276 27814 29328 27820
rect 29288 26353 29316 27814
rect 29368 27124 29420 27130
rect 29368 27066 29420 27072
rect 29380 26790 29408 27066
rect 29368 26784 29420 26790
rect 29368 26726 29420 26732
rect 29748 26450 29776 32710
rect 30116 31822 30144 33254
rect 30104 31816 30156 31822
rect 30104 31758 30156 31764
rect 30300 30802 30328 33390
rect 30380 32768 30432 32774
rect 30380 32710 30432 32716
rect 30392 31754 30420 32710
rect 30840 32428 30892 32434
rect 30840 32370 30892 32376
rect 30748 32020 30800 32026
rect 30748 31962 30800 31968
rect 30392 31726 30512 31754
rect 30288 30796 30340 30802
rect 30288 30738 30340 30744
rect 30484 30734 30512 31726
rect 30760 31278 30788 31962
rect 30748 31272 30800 31278
rect 30748 31214 30800 31220
rect 30564 31136 30616 31142
rect 30564 31078 30616 31084
rect 30104 30728 30156 30734
rect 30104 30670 30156 30676
rect 30196 30728 30248 30734
rect 30196 30670 30248 30676
rect 30472 30728 30524 30734
rect 30472 30670 30524 30676
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29840 26450 29868 29582
rect 30116 28966 30144 30670
rect 30208 30394 30236 30670
rect 30380 30592 30432 30598
rect 30380 30534 30432 30540
rect 30392 30394 30420 30534
rect 30196 30388 30248 30394
rect 30196 30330 30248 30336
rect 30380 30388 30432 30394
rect 30380 30330 30432 30336
rect 30104 28960 30156 28966
rect 30104 28902 30156 28908
rect 30116 28762 30144 28902
rect 30104 28756 30156 28762
rect 30104 28698 30156 28704
rect 30104 28076 30156 28082
rect 30104 28018 30156 28024
rect 30116 27538 30144 28018
rect 30104 27532 30156 27538
rect 30104 27474 30156 27480
rect 29920 27328 29972 27334
rect 29920 27270 29972 27276
rect 29932 26858 29960 27270
rect 29920 26852 29972 26858
rect 29920 26794 29972 26800
rect 30288 26784 30340 26790
rect 30288 26726 30340 26732
rect 29368 26444 29420 26450
rect 29368 26386 29420 26392
rect 29736 26444 29788 26450
rect 29736 26386 29788 26392
rect 29828 26444 29880 26450
rect 29828 26386 29880 26392
rect 29274 26344 29330 26353
rect 29274 26279 29330 26288
rect 29184 25424 29236 25430
rect 29184 25366 29236 25372
rect 29104 25214 29224 25242
rect 29092 25152 29144 25158
rect 29092 25094 29144 25100
rect 29104 24682 29132 25094
rect 29092 24676 29144 24682
rect 29092 24618 29144 24624
rect 29000 24404 29052 24410
rect 29000 24346 29052 24352
rect 29092 23860 29144 23866
rect 29092 23802 29144 23808
rect 28908 23792 28960 23798
rect 28908 23734 28960 23740
rect 28816 22976 28868 22982
rect 28816 22918 28868 22924
rect 29104 22438 29132 23802
rect 29092 22432 29144 22438
rect 29092 22374 29144 22380
rect 28552 22066 28672 22094
rect 28445 21548 28497 21554
rect 28445 21490 28497 21496
rect 28264 20868 28316 20874
rect 28264 20810 28316 20816
rect 28460 20398 28488 21490
rect 28644 20466 28672 22066
rect 29104 22030 29132 22374
rect 29092 22024 29144 22030
rect 29092 21966 29144 21972
rect 28724 21888 28776 21894
rect 28724 21830 28776 21836
rect 28736 21690 28764 21830
rect 28724 21684 28776 21690
rect 28724 21626 28776 21632
rect 29092 20596 29144 20602
rect 29092 20538 29144 20544
rect 28632 20460 28684 20466
rect 28632 20402 28684 20408
rect 28448 20392 28500 20398
rect 28448 20334 28500 20340
rect 29000 20392 29052 20398
rect 29000 20334 29052 20340
rect 29012 20262 29040 20334
rect 29000 20256 29052 20262
rect 29000 20198 29052 20204
rect 29012 19854 29040 20198
rect 29000 19848 29052 19854
rect 29000 19790 29052 19796
rect 28816 18624 28868 18630
rect 28816 18566 28868 18572
rect 28828 18222 28856 18566
rect 28816 18216 28868 18222
rect 28816 18158 28868 18164
rect 28724 17128 28776 17134
rect 28724 17070 28776 17076
rect 28356 16992 28408 16998
rect 28356 16934 28408 16940
rect 28368 16522 28396 16934
rect 28356 16516 28408 16522
rect 28356 16458 28408 16464
rect 28262 15056 28318 15065
rect 28262 14991 28318 15000
rect 28632 15020 28684 15026
rect 28276 14482 28304 14991
rect 28632 14962 28684 14968
rect 28264 14476 28316 14482
rect 28264 14418 28316 14424
rect 28644 14414 28672 14962
rect 28632 14408 28684 14414
rect 28632 14350 28684 14356
rect 28448 14272 28500 14278
rect 28448 14214 28500 14220
rect 28460 14006 28488 14214
rect 28644 14006 28672 14350
rect 28448 14000 28500 14006
rect 28448 13942 28500 13948
rect 28632 14000 28684 14006
rect 28632 13942 28684 13948
rect 28170 13560 28226 13569
rect 28170 13495 28226 13504
rect 28080 13320 28132 13326
rect 28080 13262 28132 13268
rect 28184 12374 28212 13495
rect 28172 12368 28224 12374
rect 28172 12310 28224 12316
rect 28356 12164 28408 12170
rect 28356 12106 28408 12112
rect 28368 11694 28396 12106
rect 28356 11688 28408 11694
rect 28356 11630 28408 11636
rect 28540 10464 28592 10470
rect 28540 10406 28592 10412
rect 27988 10260 28040 10266
rect 27988 10202 28040 10208
rect 28264 10124 28316 10130
rect 28264 10066 28316 10072
rect 28276 8838 28304 10066
rect 28448 10056 28500 10062
rect 28448 9998 28500 10004
rect 28264 8832 28316 8838
rect 28264 8774 28316 8780
rect 28276 8498 28304 8774
rect 28264 8492 28316 8498
rect 28264 8434 28316 8440
rect 27896 8356 27948 8362
rect 27896 8298 27948 8304
rect 27804 7880 27856 7886
rect 27804 7822 27856 7828
rect 28276 7818 28304 8434
rect 28264 7812 28316 7818
rect 28264 7754 28316 7760
rect 28170 7440 28226 7449
rect 27804 7404 27856 7410
rect 27804 7346 27856 7352
rect 27988 7404 28040 7410
rect 28170 7375 28172 7384
rect 27988 7346 28040 7352
rect 28224 7375 28226 7384
rect 28172 7346 28224 7352
rect 27620 7268 27672 7274
rect 27620 7210 27672 7216
rect 27816 6458 27844 7346
rect 27804 6452 27856 6458
rect 27804 6394 27856 6400
rect 28000 6322 28028 7346
rect 27988 6316 28040 6322
rect 27988 6258 28040 6264
rect 27436 5772 27488 5778
rect 27436 5714 27488 5720
rect 27804 5568 27856 5574
rect 27804 5510 27856 5516
rect 27816 5234 27844 5510
rect 28000 5234 28028 6258
rect 28460 5710 28488 9998
rect 28552 9586 28580 10406
rect 28632 10192 28684 10198
rect 28632 10134 28684 10140
rect 28540 9580 28592 9586
rect 28540 9522 28592 9528
rect 28644 8566 28672 10134
rect 28632 8560 28684 8566
rect 28632 8502 28684 8508
rect 28736 8090 28764 17070
rect 28828 10742 28856 18158
rect 29104 17678 29132 20538
rect 29196 18306 29224 25214
rect 29276 24336 29328 24342
rect 29276 24278 29328 24284
rect 29288 20346 29316 24278
rect 29380 20602 29408 26386
rect 29644 26240 29696 26246
rect 29644 26182 29696 26188
rect 30300 26194 30328 26726
rect 30392 26314 30420 30330
rect 30472 29164 30524 29170
rect 30472 29106 30524 29112
rect 30484 28558 30512 29106
rect 30472 28552 30524 28558
rect 30472 28494 30524 28500
rect 30472 26784 30524 26790
rect 30472 26726 30524 26732
rect 30380 26308 30432 26314
rect 30380 26250 30432 26256
rect 29460 24812 29512 24818
rect 29460 24754 29512 24760
rect 29472 23866 29500 24754
rect 29460 23860 29512 23866
rect 29460 23802 29512 23808
rect 29656 20942 29684 26182
rect 30300 26166 30420 26194
rect 30288 25152 30340 25158
rect 30288 25094 30340 25100
rect 30012 24268 30064 24274
rect 30012 24210 30064 24216
rect 30024 23662 30052 24210
rect 30300 24206 30328 25094
rect 30104 24200 30156 24206
rect 30104 24142 30156 24148
rect 30288 24200 30340 24206
rect 30288 24142 30340 24148
rect 30116 23730 30144 24142
rect 30104 23724 30156 23730
rect 30104 23666 30156 23672
rect 30012 23656 30064 23662
rect 30012 23598 30064 23604
rect 30012 23520 30064 23526
rect 30012 23462 30064 23468
rect 30024 22438 30052 23462
rect 30012 22432 30064 22438
rect 30012 22374 30064 22380
rect 29644 20936 29696 20942
rect 29644 20878 29696 20884
rect 29920 20936 29972 20942
rect 29920 20878 29972 20884
rect 29644 20800 29696 20806
rect 29644 20742 29696 20748
rect 29368 20596 29420 20602
rect 29368 20538 29420 20544
rect 29460 20460 29512 20466
rect 29460 20402 29512 20408
rect 29288 20318 29408 20346
rect 29380 20262 29408 20318
rect 29368 20256 29420 20262
rect 29368 20198 29420 20204
rect 29196 18290 29316 18306
rect 29196 18284 29328 18290
rect 29196 18278 29276 18284
rect 29276 18226 29328 18232
rect 29092 17672 29144 17678
rect 29092 17614 29144 17620
rect 29184 17332 29236 17338
rect 29184 17274 29236 17280
rect 28908 16516 28960 16522
rect 28908 16458 28960 16464
rect 28920 16250 28948 16458
rect 28908 16244 28960 16250
rect 28908 16186 28960 16192
rect 29092 15020 29144 15026
rect 29092 14962 29144 14968
rect 29104 14822 29132 14962
rect 29092 14816 29144 14822
rect 29092 14758 29144 14764
rect 29092 13932 29144 13938
rect 29092 13874 29144 13880
rect 29104 13802 29132 13874
rect 29092 13796 29144 13802
rect 29092 13738 29144 13744
rect 29104 12918 29132 13738
rect 29196 13190 29224 17274
rect 29288 15994 29316 18226
rect 29380 17882 29408 20198
rect 29368 17876 29420 17882
rect 29368 17818 29420 17824
rect 29368 16992 29420 16998
rect 29368 16934 29420 16940
rect 29380 16114 29408 16934
rect 29368 16108 29420 16114
rect 29368 16050 29420 16056
rect 29288 15966 29408 15994
rect 29276 13728 29328 13734
rect 29276 13670 29328 13676
rect 29184 13184 29236 13190
rect 29184 13126 29236 13132
rect 29092 12912 29144 12918
rect 29092 12854 29144 12860
rect 29092 11212 29144 11218
rect 29092 11154 29144 11160
rect 28816 10736 28868 10742
rect 28816 10678 28868 10684
rect 29104 10538 29132 11154
rect 29092 10532 29144 10538
rect 29092 10474 29144 10480
rect 29288 10198 29316 13670
rect 29380 13258 29408 15966
rect 29368 13252 29420 13258
rect 29368 13194 29420 13200
rect 29368 10532 29420 10538
rect 29368 10474 29420 10480
rect 29380 10266 29408 10474
rect 29368 10260 29420 10266
rect 29368 10202 29420 10208
rect 29276 10192 29328 10198
rect 29276 10134 29328 10140
rect 28816 10056 28868 10062
rect 28816 9998 28868 10004
rect 28828 8974 28856 9998
rect 28816 8968 28868 8974
rect 28816 8910 28868 8916
rect 28828 8430 28856 8910
rect 29276 8492 29328 8498
rect 29276 8434 29328 8440
rect 28816 8424 28868 8430
rect 28816 8366 28868 8372
rect 28724 8084 28776 8090
rect 28724 8026 28776 8032
rect 28632 7200 28684 7206
rect 28632 7142 28684 7148
rect 28644 6322 28672 7142
rect 29288 6662 29316 8434
rect 29276 6656 29328 6662
rect 29276 6598 29328 6604
rect 28632 6316 28684 6322
rect 28632 6258 28684 6264
rect 28448 5704 28500 5710
rect 28448 5646 28500 5652
rect 27804 5228 27856 5234
rect 27804 5170 27856 5176
rect 27988 5228 28040 5234
rect 27988 5170 28040 5176
rect 27252 5024 27304 5030
rect 27252 4966 27304 4972
rect 27160 4684 27212 4690
rect 27160 4626 27212 4632
rect 27264 4622 27292 4966
rect 28460 4826 28488 5646
rect 28644 5642 28672 6258
rect 29288 6254 29316 6598
rect 29472 6458 29500 20402
rect 29656 19854 29684 20742
rect 29932 20398 29960 20878
rect 29920 20392 29972 20398
rect 29920 20334 29972 20340
rect 29736 20052 29788 20058
rect 29736 19994 29788 20000
rect 29644 19848 29696 19854
rect 29644 19790 29696 19796
rect 29748 19446 29776 19994
rect 29736 19440 29788 19446
rect 29736 19382 29788 19388
rect 29828 19372 29880 19378
rect 29828 19314 29880 19320
rect 29644 18624 29696 18630
rect 29644 18566 29696 18572
rect 29656 18426 29684 18566
rect 29644 18420 29696 18426
rect 29644 18362 29696 18368
rect 29736 18080 29788 18086
rect 29736 18022 29788 18028
rect 29552 16584 29604 16590
rect 29552 16526 29604 16532
rect 29564 15502 29592 16526
rect 29552 15496 29604 15502
rect 29552 15438 29604 15444
rect 29564 13326 29592 15438
rect 29644 15428 29696 15434
rect 29644 15370 29696 15376
rect 29656 15162 29684 15370
rect 29644 15156 29696 15162
rect 29644 15098 29696 15104
rect 29644 14340 29696 14346
rect 29644 14282 29696 14288
rect 29656 14074 29684 14282
rect 29644 14068 29696 14074
rect 29644 14010 29696 14016
rect 29656 13462 29684 14010
rect 29644 13456 29696 13462
rect 29644 13398 29696 13404
rect 29552 13320 29604 13326
rect 29552 13262 29604 13268
rect 29552 13184 29604 13190
rect 29552 13126 29604 13132
rect 29564 12986 29592 13126
rect 29552 12980 29604 12986
rect 29552 12922 29604 12928
rect 29564 6882 29592 12922
rect 29748 12442 29776 18022
rect 29840 17202 29868 19314
rect 30024 18086 30052 22374
rect 30392 22094 30420 26166
rect 30484 24954 30512 26726
rect 30472 24948 30524 24954
rect 30472 24890 30524 24896
rect 30392 22066 30512 22094
rect 30484 22030 30512 22066
rect 30472 22024 30524 22030
rect 30472 21966 30524 21972
rect 30288 21480 30340 21486
rect 30288 21422 30340 21428
rect 30104 21344 30156 21350
rect 30104 21286 30156 21292
rect 30116 21146 30144 21286
rect 30104 21140 30156 21146
rect 30104 21082 30156 21088
rect 30104 20800 30156 20806
rect 30104 20742 30156 20748
rect 30116 18766 30144 20742
rect 30196 20256 30248 20262
rect 30196 20198 30248 20204
rect 30208 19990 30236 20198
rect 30196 19984 30248 19990
rect 30196 19926 30248 19932
rect 30104 18760 30156 18766
rect 30104 18702 30156 18708
rect 30012 18080 30064 18086
rect 30012 18022 30064 18028
rect 29828 17196 29880 17202
rect 29828 17138 29880 17144
rect 30012 17196 30064 17202
rect 30012 17138 30064 17144
rect 30024 16454 30052 17138
rect 30104 16516 30156 16522
rect 30104 16458 30156 16464
rect 30012 16448 30064 16454
rect 30012 16390 30064 16396
rect 30116 16130 30144 16458
rect 30024 16102 30144 16130
rect 30196 16108 30248 16114
rect 30024 16046 30052 16102
rect 30196 16050 30248 16056
rect 30012 16040 30064 16046
rect 30012 15982 30064 15988
rect 30104 16040 30156 16046
rect 30104 15982 30156 15988
rect 30024 15722 30052 15982
rect 29932 15706 30052 15722
rect 29920 15700 30052 15706
rect 29972 15694 30052 15700
rect 29920 15642 29972 15648
rect 30012 15360 30064 15366
rect 30012 15302 30064 15308
rect 29920 15156 29972 15162
rect 29920 15098 29972 15104
rect 29828 14272 29880 14278
rect 29828 14214 29880 14220
rect 29840 13938 29868 14214
rect 29828 13932 29880 13938
rect 29828 13874 29880 13880
rect 29932 13394 29960 15098
rect 30024 14074 30052 15302
rect 30116 14822 30144 15982
rect 30208 15366 30236 16050
rect 30196 15360 30248 15366
rect 30196 15302 30248 15308
rect 30104 14816 30156 14822
rect 30104 14758 30156 14764
rect 30012 14068 30064 14074
rect 30012 14010 30064 14016
rect 30116 13870 30144 14758
rect 30208 14006 30236 15302
rect 30196 14000 30248 14006
rect 30196 13942 30248 13948
rect 30104 13864 30156 13870
rect 30104 13806 30156 13812
rect 29920 13388 29972 13394
rect 29920 13330 29972 13336
rect 30104 13252 30156 13258
rect 30104 13194 30156 13200
rect 29736 12436 29788 12442
rect 29736 12378 29788 12384
rect 29644 9988 29696 9994
rect 29644 9930 29696 9936
rect 29656 9722 29684 9930
rect 29644 9716 29696 9722
rect 30116 9674 30144 13194
rect 30196 11348 30248 11354
rect 30196 11290 30248 11296
rect 30208 11150 30236 11290
rect 30196 11144 30248 11150
rect 30196 11086 30248 11092
rect 29644 9658 29696 9664
rect 29828 9648 29880 9654
rect 29828 9590 29880 9596
rect 29932 9646 30144 9674
rect 29840 7342 29868 9590
rect 29828 7336 29880 7342
rect 29828 7278 29880 7284
rect 29564 6854 29684 6882
rect 29460 6452 29512 6458
rect 29460 6394 29512 6400
rect 29276 6248 29328 6254
rect 29276 6190 29328 6196
rect 28632 5636 28684 5642
rect 28632 5578 28684 5584
rect 28448 4820 28500 4826
rect 28448 4762 28500 4768
rect 27252 4616 27304 4622
rect 27252 4558 27304 4564
rect 26700 3528 26752 3534
rect 26700 3470 26752 3476
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 28632 3528 28684 3534
rect 28632 3470 28684 3476
rect 26330 2952 26386 2961
rect 26330 2887 26386 2896
rect 26148 2848 26200 2854
rect 26148 2790 26200 2796
rect 25872 2440 25924 2446
rect 25872 2382 25924 2388
rect 25884 800 25912 2382
rect 26160 800 26188 2790
rect 26424 2576 26476 2582
rect 26424 2518 26476 2524
rect 26436 800 26464 2518
rect 26712 800 26740 3470
rect 26976 2848 27028 2854
rect 26976 2790 27028 2796
rect 26988 800 27016 2790
rect 27252 2440 27304 2446
rect 27252 2382 27304 2388
rect 27264 800 27292 2382
rect 27540 800 27568 3470
rect 27804 2848 27856 2854
rect 27804 2790 27856 2796
rect 28080 2848 28132 2854
rect 28080 2790 28132 2796
rect 27816 800 27844 2790
rect 28092 800 28120 2790
rect 28356 2576 28408 2582
rect 28356 2518 28408 2524
rect 28368 800 28396 2518
rect 28644 800 28672 3470
rect 29184 2848 29236 2854
rect 29184 2790 29236 2796
rect 28908 2440 28960 2446
rect 28908 2382 28960 2388
rect 28920 800 28948 2382
rect 29196 800 29224 2790
rect 29472 2774 29500 6394
rect 29550 5672 29606 5681
rect 29550 5607 29606 5616
rect 29564 5574 29592 5607
rect 29552 5568 29604 5574
rect 29552 5510 29604 5516
rect 29380 2746 29500 2774
rect 29380 2417 29408 2746
rect 29460 2440 29512 2446
rect 29366 2408 29422 2417
rect 29460 2382 29512 2388
rect 29366 2343 29422 2352
rect 29472 800 29500 2382
rect 29564 1970 29592 5510
rect 29656 5166 29684 6854
rect 29840 6798 29868 7278
rect 29828 6792 29880 6798
rect 29828 6734 29880 6740
rect 29932 5681 29960 9646
rect 30300 8634 30328 21422
rect 30472 19848 30524 19854
rect 30472 19790 30524 19796
rect 30380 19440 30432 19446
rect 30380 19382 30432 19388
rect 30392 18834 30420 19382
rect 30484 19378 30512 19790
rect 30472 19372 30524 19378
rect 30472 19314 30524 19320
rect 30472 19168 30524 19174
rect 30472 19110 30524 19116
rect 30484 18970 30512 19110
rect 30472 18964 30524 18970
rect 30472 18906 30524 18912
rect 30380 18828 30432 18834
rect 30380 18770 30432 18776
rect 30576 18766 30604 31078
rect 30760 29238 30788 31214
rect 30748 29232 30800 29238
rect 30748 29174 30800 29180
rect 30760 28626 30788 29174
rect 30748 28620 30800 28626
rect 30748 28562 30800 28568
rect 30852 28218 30880 32370
rect 30944 31822 30972 33476
rect 31128 33386 31156 37742
rect 31680 37398 31708 37742
rect 31668 37392 31720 37398
rect 31668 37334 31720 37340
rect 31680 37262 31708 37334
rect 31668 37256 31720 37262
rect 31668 37198 31720 37204
rect 31392 36712 31444 36718
rect 31392 36654 31444 36660
rect 31404 36174 31432 36654
rect 31392 36168 31444 36174
rect 31392 36110 31444 36116
rect 31208 35012 31260 35018
rect 31208 34954 31260 34960
rect 31220 33930 31248 34954
rect 31576 34944 31628 34950
rect 31576 34886 31628 34892
rect 31588 34746 31616 34886
rect 31576 34740 31628 34746
rect 31576 34682 31628 34688
rect 31208 33924 31260 33930
rect 31208 33866 31260 33872
rect 31392 33924 31444 33930
rect 31392 33866 31444 33872
rect 31116 33380 31168 33386
rect 31116 33322 31168 33328
rect 31024 32020 31076 32026
rect 31024 31962 31076 31968
rect 30932 31816 30984 31822
rect 30932 31758 30984 31764
rect 30932 31340 30984 31346
rect 30932 31282 30984 31288
rect 30944 30258 30972 31282
rect 31036 30326 31064 31962
rect 31024 30320 31076 30326
rect 31024 30262 31076 30268
rect 30932 30252 30984 30258
rect 30932 30194 30984 30200
rect 31128 29850 31156 33322
rect 31220 32570 31248 33866
rect 31208 32564 31260 32570
rect 31208 32506 31260 32512
rect 31404 32026 31432 33866
rect 31392 32020 31444 32026
rect 31392 31962 31444 31968
rect 31588 31414 31616 34682
rect 31680 33522 31708 37198
rect 31956 37126 31984 38286
rect 31944 37120 31996 37126
rect 31944 37062 31996 37068
rect 31760 35692 31812 35698
rect 31760 35634 31812 35640
rect 31772 35086 31800 35634
rect 31760 35080 31812 35086
rect 31760 35022 31812 35028
rect 31668 33516 31720 33522
rect 31668 33458 31720 33464
rect 31772 32910 31800 35022
rect 31760 32904 31812 32910
rect 31760 32846 31812 32852
rect 31576 31408 31628 31414
rect 31576 31350 31628 31356
rect 31956 31346 31984 37062
rect 31208 31340 31260 31346
rect 31208 31282 31260 31288
rect 31944 31340 31996 31346
rect 31944 31282 31996 31288
rect 31220 30666 31248 31282
rect 31208 30660 31260 30666
rect 31208 30602 31260 30608
rect 31220 30326 31248 30602
rect 31208 30320 31260 30326
rect 31208 30262 31260 30268
rect 32048 30258 32076 39306
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 32312 38208 32364 38214
rect 32312 38150 32364 38156
rect 32324 37262 32352 38150
rect 32588 37868 32640 37874
rect 32588 37810 32640 37816
rect 32312 37256 32364 37262
rect 32312 37198 32364 37204
rect 32324 36310 32352 37198
rect 32600 36922 32628 37810
rect 33784 37664 33836 37670
rect 33784 37606 33836 37612
rect 35532 37664 35584 37670
rect 35532 37606 35584 37612
rect 33508 37256 33560 37262
rect 33508 37198 33560 37204
rect 32588 36916 32640 36922
rect 32588 36858 32640 36864
rect 33416 36916 33468 36922
rect 33416 36858 33468 36864
rect 33140 36780 33192 36786
rect 33140 36722 33192 36728
rect 32312 36304 32364 36310
rect 32312 36246 32364 36252
rect 33152 35834 33180 36722
rect 33428 36038 33456 36858
rect 33520 36786 33548 37198
rect 33508 36780 33560 36786
rect 33508 36722 33560 36728
rect 33520 36174 33548 36722
rect 33508 36168 33560 36174
rect 33508 36110 33560 36116
rect 33416 36032 33468 36038
rect 33416 35974 33468 35980
rect 33140 35828 33192 35834
rect 33140 35770 33192 35776
rect 33324 35216 33376 35222
rect 33324 35158 33376 35164
rect 33336 34406 33364 35158
rect 33324 34400 33376 34406
rect 33324 34342 33376 34348
rect 32312 33584 32364 33590
rect 32312 33526 32364 33532
rect 32324 32978 32352 33526
rect 32956 33516 33008 33522
rect 32956 33458 33008 33464
rect 32312 32972 32364 32978
rect 32312 32914 32364 32920
rect 32128 32904 32180 32910
rect 32128 32846 32180 32852
rect 32140 31482 32168 32846
rect 32324 32502 32352 32914
rect 32404 32768 32456 32774
rect 32404 32710 32456 32716
rect 32312 32496 32364 32502
rect 32312 32438 32364 32444
rect 32128 31476 32180 31482
rect 32128 31418 32180 31424
rect 32220 31136 32272 31142
rect 32220 31078 32272 31084
rect 32232 30734 32260 31078
rect 32324 30870 32352 32438
rect 32416 32434 32444 32710
rect 32968 32570 32996 33458
rect 32956 32564 33008 32570
rect 32956 32506 33008 32512
rect 32404 32428 32456 32434
rect 32404 32370 32456 32376
rect 32588 32428 32640 32434
rect 32588 32370 32640 32376
rect 32600 32026 32628 32370
rect 32588 32020 32640 32026
rect 32588 31962 32640 31968
rect 32404 31680 32456 31686
rect 32404 31622 32456 31628
rect 32416 31346 32444 31622
rect 32404 31340 32456 31346
rect 32404 31282 32456 31288
rect 32312 30864 32364 30870
rect 32312 30806 32364 30812
rect 32220 30728 32272 30734
rect 32220 30670 32272 30676
rect 32036 30252 32088 30258
rect 32036 30194 32088 30200
rect 31208 30116 31260 30122
rect 31208 30058 31260 30064
rect 31116 29844 31168 29850
rect 31116 29786 31168 29792
rect 30932 29640 30984 29646
rect 30932 29582 30984 29588
rect 30840 28212 30892 28218
rect 30840 28154 30892 28160
rect 30748 28144 30800 28150
rect 30748 28086 30800 28092
rect 30760 22094 30788 28086
rect 30852 27402 30880 28154
rect 30840 27396 30892 27402
rect 30840 27338 30892 27344
rect 30944 27062 30972 29582
rect 31220 29034 31248 30058
rect 31392 30048 31444 30054
rect 31392 29990 31444 29996
rect 31208 29028 31260 29034
rect 31208 28970 31260 28976
rect 30932 27056 30984 27062
rect 30932 26998 30984 27004
rect 30840 26308 30892 26314
rect 30840 26250 30892 26256
rect 30852 26042 30880 26250
rect 30840 26036 30892 26042
rect 30840 25978 30892 25984
rect 30944 25906 30972 26998
rect 30932 25900 30984 25906
rect 30932 25842 30984 25848
rect 30944 25294 30972 25842
rect 30932 25288 30984 25294
rect 30932 25230 30984 25236
rect 30944 24818 30972 25230
rect 31024 24880 31076 24886
rect 31024 24822 31076 24828
rect 30932 24812 30984 24818
rect 30932 24754 30984 24760
rect 30760 22066 30880 22094
rect 30852 21010 30880 22066
rect 30932 21548 30984 21554
rect 30932 21490 30984 21496
rect 30944 21146 30972 21490
rect 30932 21140 30984 21146
rect 30932 21082 30984 21088
rect 30840 21004 30892 21010
rect 30840 20946 30892 20952
rect 30654 20496 30710 20505
rect 30654 20431 30710 20440
rect 30668 19174 30696 20431
rect 30932 19712 30984 19718
rect 30932 19654 30984 19660
rect 30840 19304 30892 19310
rect 30840 19246 30892 19252
rect 30656 19168 30708 19174
rect 30656 19110 30708 19116
rect 30564 18760 30616 18766
rect 30564 18702 30616 18708
rect 30564 18624 30616 18630
rect 30564 18566 30616 18572
rect 30576 18358 30604 18566
rect 30564 18352 30616 18358
rect 30564 18294 30616 18300
rect 30380 17876 30432 17882
rect 30380 17818 30432 17824
rect 30392 11354 30420 17818
rect 30656 17264 30708 17270
rect 30656 17206 30708 17212
rect 30472 15360 30524 15366
rect 30472 15302 30524 15308
rect 30484 15026 30512 15302
rect 30472 15020 30524 15026
rect 30472 14962 30524 14968
rect 30380 11348 30432 11354
rect 30380 11290 30432 11296
rect 30472 11076 30524 11082
rect 30472 11018 30524 11024
rect 30564 11076 30616 11082
rect 30564 11018 30616 11024
rect 30484 9586 30512 11018
rect 30576 10674 30604 11018
rect 30564 10668 30616 10674
rect 30564 10610 30616 10616
rect 30668 10266 30696 17206
rect 30748 13864 30800 13870
rect 30748 13806 30800 13812
rect 30760 13258 30788 13806
rect 30852 13734 30880 19246
rect 30944 18902 30972 19654
rect 31036 19446 31064 24822
rect 31116 20868 31168 20874
rect 31116 20810 31168 20816
rect 31128 20602 31156 20810
rect 31404 20806 31432 29990
rect 32324 29306 32352 30806
rect 32312 29300 32364 29306
rect 32312 29242 32364 29248
rect 31484 28416 31536 28422
rect 31484 28358 31536 28364
rect 31496 28150 31524 28358
rect 31484 28144 31536 28150
rect 31484 28086 31536 28092
rect 32416 27946 32444 31282
rect 32600 29034 32628 31962
rect 33428 31958 33456 35974
rect 33520 34610 33548 36110
rect 33692 36100 33744 36106
rect 33692 36042 33744 36048
rect 33704 35698 33732 36042
rect 33796 35766 33824 37606
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34888 37392 34940 37398
rect 34888 37334 34940 37340
rect 34152 37188 34204 37194
rect 34152 37130 34204 37136
rect 33876 37120 33928 37126
rect 33876 37062 33928 37068
rect 33888 36854 33916 37062
rect 33876 36848 33928 36854
rect 33876 36790 33928 36796
rect 33784 35760 33836 35766
rect 33784 35702 33836 35708
rect 33692 35692 33744 35698
rect 33692 35634 33744 35640
rect 33704 35494 33732 35634
rect 33692 35488 33744 35494
rect 33692 35430 33744 35436
rect 33508 34604 33560 34610
rect 33508 34546 33560 34552
rect 33520 33998 33548 34546
rect 33704 34134 33732 35430
rect 33692 34128 33744 34134
rect 33692 34070 33744 34076
rect 33508 33992 33560 33998
rect 33508 33934 33560 33940
rect 33520 32366 33548 33934
rect 33508 32360 33560 32366
rect 33508 32302 33560 32308
rect 33416 31952 33468 31958
rect 33416 31894 33468 31900
rect 33232 31340 33284 31346
rect 33232 31282 33284 31288
rect 33140 30592 33192 30598
rect 33140 30534 33192 30540
rect 33152 30326 33180 30534
rect 33140 30320 33192 30326
rect 33140 30262 33192 30268
rect 33244 30054 33272 31282
rect 33508 31272 33560 31278
rect 33508 31214 33560 31220
rect 33324 30796 33376 30802
rect 33324 30738 33376 30744
rect 33232 30048 33284 30054
rect 33232 29990 33284 29996
rect 32588 29028 32640 29034
rect 32588 28970 32640 28976
rect 32404 27940 32456 27946
rect 32404 27882 32456 27888
rect 32600 26382 32628 28970
rect 33140 28008 33192 28014
rect 33140 27950 33192 27956
rect 32956 27872 33008 27878
rect 32956 27814 33008 27820
rect 32588 26376 32640 26382
rect 32588 26318 32640 26324
rect 31760 25220 31812 25226
rect 31760 25162 31812 25168
rect 31772 24410 31800 25162
rect 32968 24886 32996 27814
rect 33152 27010 33180 27950
rect 33060 26994 33180 27010
rect 33244 26994 33272 29990
rect 33336 29510 33364 30738
rect 33520 30734 33548 31214
rect 33796 30734 33824 35702
rect 33888 34728 33916 36790
rect 34164 36378 34192 37130
rect 34900 36786 34928 37334
rect 35544 37274 35572 37606
rect 35544 37262 35664 37274
rect 35544 37256 35676 37262
rect 35544 37246 35624 37256
rect 35624 37198 35676 37204
rect 35348 37120 35400 37126
rect 35348 37062 35400 37068
rect 34244 36780 34296 36786
rect 34244 36722 34296 36728
rect 34888 36780 34940 36786
rect 34888 36722 34940 36728
rect 34152 36372 34204 36378
rect 34152 36314 34204 36320
rect 34256 35562 34284 36722
rect 34704 36712 34756 36718
rect 34900 36666 34928 36722
rect 34704 36654 34756 36660
rect 34716 36378 34744 36654
rect 34808 36638 34928 36666
rect 34704 36372 34756 36378
rect 34704 36314 34756 36320
rect 34808 36242 34836 36638
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34796 36236 34848 36242
rect 34796 36178 34848 36184
rect 35360 36174 35388 37062
rect 35440 36916 35492 36922
rect 35440 36858 35492 36864
rect 35348 36168 35400 36174
rect 35348 36110 35400 36116
rect 35452 36106 35480 36858
rect 35440 36100 35492 36106
rect 35440 36042 35492 36048
rect 34704 36032 34756 36038
rect 34704 35974 34756 35980
rect 34244 35556 34296 35562
rect 34244 35498 34296 35504
rect 34244 34944 34296 34950
rect 34244 34886 34296 34892
rect 33968 34740 34020 34746
rect 33888 34700 33968 34728
rect 33968 34682 34020 34688
rect 33876 34400 33928 34406
rect 33876 34342 33928 34348
rect 33888 33998 33916 34342
rect 33980 34066 34008 34682
rect 34256 34610 34284 34886
rect 34244 34604 34296 34610
rect 34244 34546 34296 34552
rect 33968 34060 34020 34066
rect 33968 34002 34020 34008
rect 33876 33992 33928 33998
rect 33876 33934 33928 33940
rect 33416 30728 33468 30734
rect 33416 30670 33468 30676
rect 33508 30728 33560 30734
rect 33508 30670 33560 30676
rect 33784 30728 33836 30734
rect 33784 30670 33836 30676
rect 33428 30258 33456 30670
rect 33600 30660 33652 30666
rect 33600 30602 33652 30608
rect 33416 30252 33468 30258
rect 33416 30194 33468 30200
rect 33428 29646 33456 30194
rect 33416 29640 33468 29646
rect 33416 29582 33468 29588
rect 33324 29504 33376 29510
rect 33324 29446 33376 29452
rect 33336 28506 33364 29446
rect 33428 29170 33456 29582
rect 33612 29578 33640 30602
rect 33888 30598 33916 33934
rect 33980 32978 34008 34002
rect 34152 33856 34204 33862
rect 34152 33798 34204 33804
rect 34164 33590 34192 33798
rect 34152 33584 34204 33590
rect 34152 33526 34204 33532
rect 34152 33312 34204 33318
rect 34152 33254 34204 33260
rect 33968 32972 34020 32978
rect 33968 32914 34020 32920
rect 34164 32842 34192 33254
rect 34152 32836 34204 32842
rect 34152 32778 34204 32784
rect 34060 30864 34112 30870
rect 34060 30806 34112 30812
rect 33876 30592 33928 30598
rect 33876 30534 33928 30540
rect 33600 29572 33652 29578
rect 33600 29514 33652 29520
rect 33876 29572 33928 29578
rect 33876 29514 33928 29520
rect 33888 29238 33916 29514
rect 33876 29232 33928 29238
rect 33876 29174 33928 29180
rect 33416 29164 33468 29170
rect 33416 29106 33468 29112
rect 33428 28626 33456 29106
rect 33508 29028 33560 29034
rect 33508 28970 33560 28976
rect 33416 28620 33468 28626
rect 33416 28562 33468 28568
rect 33336 28478 33456 28506
rect 33324 27464 33376 27470
rect 33324 27406 33376 27412
rect 33336 27062 33364 27406
rect 33324 27056 33376 27062
rect 33324 26998 33376 27004
rect 33048 26988 33180 26994
rect 33100 26982 33180 26988
rect 33232 26988 33284 26994
rect 33048 26930 33100 26936
rect 33232 26930 33284 26936
rect 33140 26376 33192 26382
rect 33140 26318 33192 26324
rect 33048 26240 33100 26246
rect 33048 26182 33100 26188
rect 33060 25906 33088 26182
rect 33152 26042 33180 26318
rect 33232 26240 33284 26246
rect 33232 26182 33284 26188
rect 33140 26036 33192 26042
rect 33140 25978 33192 25984
rect 33244 25974 33272 26182
rect 33232 25968 33284 25974
rect 33232 25910 33284 25916
rect 33048 25900 33100 25906
rect 33048 25842 33100 25848
rect 33060 25362 33088 25842
rect 33336 25702 33364 26998
rect 33428 26382 33456 28478
rect 33416 26376 33468 26382
rect 33416 26318 33468 26324
rect 33324 25696 33376 25702
rect 33324 25638 33376 25644
rect 33048 25356 33100 25362
rect 33048 25298 33100 25304
rect 32956 24880 33008 24886
rect 32956 24822 33008 24828
rect 31760 24404 31812 24410
rect 31760 24346 31812 24352
rect 31576 24064 31628 24070
rect 31576 24006 31628 24012
rect 31588 23594 31616 24006
rect 31576 23588 31628 23594
rect 31576 23530 31628 23536
rect 31392 20800 31444 20806
rect 31392 20742 31444 20748
rect 31116 20596 31168 20602
rect 31116 20538 31168 20544
rect 31116 19984 31168 19990
rect 31116 19926 31168 19932
rect 31024 19440 31076 19446
rect 31024 19382 31076 19388
rect 31128 19174 31156 19926
rect 31484 19848 31536 19854
rect 31484 19790 31536 19796
rect 31208 19780 31260 19786
rect 31208 19722 31260 19728
rect 31116 19168 31168 19174
rect 31116 19110 31168 19116
rect 30932 18896 30984 18902
rect 30932 18838 30984 18844
rect 30932 18760 30984 18766
rect 30932 18702 30984 18708
rect 30944 17134 30972 18702
rect 30932 17128 30984 17134
rect 30932 17070 30984 17076
rect 31220 15706 31248 19722
rect 31496 19242 31524 19790
rect 31484 19236 31536 19242
rect 31484 19178 31536 19184
rect 31300 17672 31352 17678
rect 31300 17614 31352 17620
rect 31312 16794 31340 17614
rect 31392 17196 31444 17202
rect 31392 17138 31444 17144
rect 31300 16788 31352 16794
rect 31300 16730 31352 16736
rect 31312 16114 31340 16730
rect 31300 16108 31352 16114
rect 31300 16050 31352 16056
rect 31404 15910 31432 17138
rect 31588 17134 31616 23530
rect 32220 23316 32272 23322
rect 32220 23258 32272 23264
rect 31852 23044 31904 23050
rect 31852 22986 31904 22992
rect 31864 22642 31892 22986
rect 31852 22636 31904 22642
rect 31852 22578 31904 22584
rect 32128 22568 32180 22574
rect 32128 22510 32180 22516
rect 32140 22438 32168 22510
rect 32128 22432 32180 22438
rect 32128 22374 32180 22380
rect 32232 22030 32260 23258
rect 33048 23180 33100 23186
rect 33048 23122 33100 23128
rect 32772 22976 32824 22982
rect 32772 22918 32824 22924
rect 32588 22704 32640 22710
rect 32588 22646 32640 22652
rect 32496 22636 32548 22642
rect 32496 22578 32548 22584
rect 32220 22024 32272 22030
rect 32220 21966 32272 21972
rect 32404 22024 32456 22030
rect 32404 21966 32456 21972
rect 31668 20596 31720 20602
rect 31668 20538 31720 20544
rect 31680 19854 31708 20538
rect 31760 20460 31812 20466
rect 31760 20402 31812 20408
rect 32036 20460 32088 20466
rect 32036 20402 32088 20408
rect 31772 19922 31800 20402
rect 31760 19916 31812 19922
rect 31760 19858 31812 19864
rect 31668 19848 31720 19854
rect 31668 19790 31720 19796
rect 32048 19334 32076 20402
rect 32232 20346 32260 21966
rect 32416 20534 32444 21966
rect 32404 20528 32456 20534
rect 32404 20470 32456 20476
rect 32508 20466 32536 22578
rect 32600 20534 32628 22646
rect 32680 22500 32732 22506
rect 32680 22442 32732 22448
rect 32692 21690 32720 22442
rect 32784 21962 32812 22918
rect 33060 22658 33088 23122
rect 33416 23112 33468 23118
rect 33416 23054 33468 23060
rect 33232 23044 33284 23050
rect 33232 22986 33284 22992
rect 33324 23044 33376 23050
rect 33324 22986 33376 22992
rect 33060 22642 33180 22658
rect 32864 22636 32916 22642
rect 32864 22578 32916 22584
rect 33060 22636 33192 22642
rect 33060 22630 33140 22636
rect 32876 22506 32904 22578
rect 32864 22500 32916 22506
rect 32864 22442 32916 22448
rect 32956 22092 33008 22098
rect 32956 22034 33008 22040
rect 32772 21956 32824 21962
rect 32772 21898 32824 21904
rect 32680 21684 32732 21690
rect 32680 21626 32732 21632
rect 32784 21622 32812 21898
rect 32968 21690 32996 22034
rect 33060 22030 33088 22630
rect 33140 22578 33192 22584
rect 33048 22024 33100 22030
rect 33048 21966 33100 21972
rect 33048 21888 33100 21894
rect 33048 21830 33100 21836
rect 32956 21684 33008 21690
rect 32956 21626 33008 21632
rect 32772 21616 32824 21622
rect 32772 21558 32824 21564
rect 32772 21480 32824 21486
rect 32772 21422 32824 21428
rect 32588 20528 32640 20534
rect 32588 20470 32640 20476
rect 32496 20460 32548 20466
rect 32496 20402 32548 20408
rect 32140 20318 32260 20346
rect 32140 20058 32168 20318
rect 32220 20256 32272 20262
rect 32220 20198 32272 20204
rect 32128 20052 32180 20058
rect 32128 19994 32180 20000
rect 32140 19786 32168 19994
rect 32128 19780 32180 19786
rect 32128 19722 32180 19728
rect 31956 19306 32076 19334
rect 31956 18766 31984 19306
rect 32232 19242 32260 20198
rect 32600 19334 32628 20470
rect 32680 20460 32732 20466
rect 32680 20402 32732 20408
rect 32692 20058 32720 20402
rect 32680 20052 32732 20058
rect 32680 19994 32732 20000
rect 32784 19786 32812 21422
rect 33060 21078 33088 21830
rect 33244 21350 33272 22986
rect 33336 22778 33364 22986
rect 33324 22772 33376 22778
rect 33324 22714 33376 22720
rect 33324 22024 33376 22030
rect 33324 21966 33376 21972
rect 33232 21344 33284 21350
rect 33232 21286 33284 21292
rect 33048 21072 33100 21078
rect 33048 21014 33100 21020
rect 33336 20806 33364 21966
rect 32864 20800 32916 20806
rect 32864 20742 32916 20748
rect 33324 20800 33376 20806
rect 33324 20742 33376 20748
rect 32876 20466 32904 20742
rect 32864 20460 32916 20466
rect 32864 20402 32916 20408
rect 32876 20330 32904 20402
rect 32864 20324 32916 20330
rect 32864 20266 32916 20272
rect 32772 19780 32824 19786
rect 32772 19722 32824 19728
rect 32600 19306 32720 19334
rect 32220 19236 32272 19242
rect 32220 19178 32272 19184
rect 31944 18760 31996 18766
rect 31944 18702 31996 18708
rect 31668 18624 31720 18630
rect 31668 18566 31720 18572
rect 31680 18222 31708 18566
rect 31944 18352 31996 18358
rect 31944 18294 31996 18300
rect 31668 18216 31720 18222
rect 31668 18158 31720 18164
rect 31956 17814 31984 18294
rect 32232 18290 32260 19178
rect 32496 18896 32548 18902
rect 32496 18838 32548 18844
rect 32508 18426 32536 18838
rect 32692 18834 32720 19306
rect 32680 18828 32732 18834
rect 32680 18770 32732 18776
rect 32496 18420 32548 18426
rect 32496 18362 32548 18368
rect 32220 18284 32272 18290
rect 32220 18226 32272 18232
rect 32588 18080 32640 18086
rect 32588 18022 32640 18028
rect 31944 17808 31996 17814
rect 31944 17750 31996 17756
rect 31956 17678 31984 17750
rect 31944 17672 31996 17678
rect 31944 17614 31996 17620
rect 32404 17672 32456 17678
rect 32404 17614 32456 17620
rect 32416 17202 32444 17614
rect 32600 17202 32628 18022
rect 32692 17954 32720 18770
rect 32784 18358 32812 19722
rect 32772 18352 32824 18358
rect 32772 18294 32824 18300
rect 32692 17926 32812 17954
rect 32784 17814 32812 17926
rect 32772 17808 32824 17814
rect 32772 17750 32824 17756
rect 32784 17202 32812 17750
rect 32404 17196 32456 17202
rect 32404 17138 32456 17144
rect 32588 17196 32640 17202
rect 32772 17196 32824 17202
rect 32588 17138 32640 17144
rect 32692 17156 32772 17184
rect 31576 17128 31628 17134
rect 31576 17070 31628 17076
rect 31588 16998 31616 17070
rect 31576 16992 31628 16998
rect 31576 16934 31628 16940
rect 31392 15904 31444 15910
rect 31392 15846 31444 15852
rect 31208 15700 31260 15706
rect 31208 15642 31260 15648
rect 31220 15502 31248 15642
rect 31208 15496 31260 15502
rect 31208 15438 31260 15444
rect 31404 15434 31432 15846
rect 31392 15428 31444 15434
rect 31392 15370 31444 15376
rect 31404 14414 31432 15370
rect 31392 14408 31444 14414
rect 31392 14350 31444 14356
rect 30840 13728 30892 13734
rect 30840 13670 30892 13676
rect 30748 13252 30800 13258
rect 30748 13194 30800 13200
rect 31588 12986 31616 16934
rect 31760 15360 31812 15366
rect 31760 15302 31812 15308
rect 31772 15094 31800 15302
rect 31760 15088 31812 15094
rect 31760 15030 31812 15036
rect 32416 15026 32444 17138
rect 32692 16590 32720 17156
rect 32772 17138 32824 17144
rect 32680 16584 32732 16590
rect 32680 16526 32732 16532
rect 32496 16108 32548 16114
rect 32496 16050 32548 16056
rect 32508 15366 32536 16050
rect 32496 15360 32548 15366
rect 32496 15302 32548 15308
rect 32404 15020 32456 15026
rect 32404 14962 32456 14968
rect 32508 13530 32536 15302
rect 32496 13524 32548 13530
rect 32496 13466 32548 13472
rect 31944 13252 31996 13258
rect 31944 13194 31996 13200
rect 32128 13252 32180 13258
rect 32128 13194 32180 13200
rect 31576 12980 31628 12986
rect 31576 12922 31628 12928
rect 31300 12844 31352 12850
rect 31300 12786 31352 12792
rect 31312 12238 31340 12786
rect 31852 12776 31904 12782
rect 31852 12718 31904 12724
rect 31300 12232 31352 12238
rect 31300 12174 31352 12180
rect 31484 12232 31536 12238
rect 31484 12174 31536 12180
rect 30748 11756 30800 11762
rect 30748 11698 30800 11704
rect 30760 10742 30788 11698
rect 31312 11150 31340 12174
rect 31496 11898 31524 12174
rect 31864 12170 31892 12718
rect 31852 12164 31904 12170
rect 31852 12106 31904 12112
rect 31484 11892 31536 11898
rect 31484 11834 31536 11840
rect 31864 11218 31892 12106
rect 31956 11762 31984 13194
rect 32036 12232 32088 12238
rect 32036 12174 32088 12180
rect 32048 12102 32076 12174
rect 32036 12096 32088 12102
rect 32036 12038 32088 12044
rect 31944 11756 31996 11762
rect 31944 11698 31996 11704
rect 31852 11212 31904 11218
rect 31852 11154 31904 11160
rect 30840 11144 30892 11150
rect 30840 11086 30892 11092
rect 31300 11144 31352 11150
rect 31300 11086 31352 11092
rect 30852 10810 30880 11086
rect 30840 10804 30892 10810
rect 30840 10746 30892 10752
rect 30748 10736 30800 10742
rect 30748 10678 30800 10684
rect 30656 10260 30708 10266
rect 30656 10202 30708 10208
rect 30668 10062 30696 10202
rect 30656 10056 30708 10062
rect 30656 9998 30708 10004
rect 30760 9994 30788 10678
rect 30840 10668 30892 10674
rect 30840 10610 30892 10616
rect 30748 9988 30800 9994
rect 30748 9930 30800 9936
rect 30472 9580 30524 9586
rect 30472 9522 30524 9528
rect 30760 8974 30788 9930
rect 30852 9722 30880 10610
rect 30840 9716 30892 9722
rect 30840 9658 30892 9664
rect 31576 9716 31628 9722
rect 31576 9658 31628 9664
rect 31588 9042 31616 9658
rect 31864 9654 31892 11154
rect 32036 11144 32088 11150
rect 32036 11086 32088 11092
rect 31852 9648 31904 9654
rect 31852 9590 31904 9596
rect 32048 9586 32076 11086
rect 32036 9580 32088 9586
rect 32036 9522 32088 9528
rect 31576 9036 31628 9042
rect 31576 8978 31628 8984
rect 30748 8968 30800 8974
rect 30748 8910 30800 8916
rect 31668 8968 31720 8974
rect 31668 8910 31720 8916
rect 31392 8900 31444 8906
rect 31392 8842 31444 8848
rect 30288 8628 30340 8634
rect 30288 8570 30340 8576
rect 31404 8566 31432 8842
rect 31392 8560 31444 8566
rect 31392 8502 31444 8508
rect 30656 7744 30708 7750
rect 30656 7686 30708 7692
rect 30472 7404 30524 7410
rect 30472 7346 30524 7352
rect 30012 6792 30064 6798
rect 30012 6734 30064 6740
rect 30024 6390 30052 6734
rect 30116 6458 30328 6474
rect 30484 6458 30512 7346
rect 30104 6452 30328 6458
rect 30156 6446 30328 6452
rect 30104 6394 30156 6400
rect 30012 6384 30064 6390
rect 30012 6326 30064 6332
rect 30300 6322 30328 6446
rect 30472 6452 30524 6458
rect 30472 6394 30524 6400
rect 30668 6322 30696 7686
rect 31404 6662 31432 8502
rect 31680 7886 31708 8910
rect 32140 8634 32168 13194
rect 32404 13184 32456 13190
rect 32404 13126 32456 13132
rect 32416 12850 32444 13126
rect 32404 12844 32456 12850
rect 32404 12786 32456 12792
rect 32404 12096 32456 12102
rect 32404 12038 32456 12044
rect 32416 11762 32444 12038
rect 32404 11756 32456 11762
rect 32404 11698 32456 11704
rect 32312 11620 32364 11626
rect 32312 11562 32364 11568
rect 32324 11150 32352 11562
rect 32312 11144 32364 11150
rect 32312 11086 32364 11092
rect 32508 10266 32536 13466
rect 32496 10260 32548 10266
rect 32496 10202 32548 10208
rect 32312 9580 32364 9586
rect 32312 9522 32364 9528
rect 32324 9178 32352 9522
rect 32312 9172 32364 9178
rect 32312 9114 32364 9120
rect 32404 8968 32456 8974
rect 32404 8910 32456 8916
rect 32312 8900 32364 8906
rect 32312 8842 32364 8848
rect 32128 8628 32180 8634
rect 32128 8570 32180 8576
rect 32324 8566 32352 8842
rect 32312 8560 32364 8566
rect 32312 8502 32364 8508
rect 32128 8492 32180 8498
rect 32128 8434 32180 8440
rect 31668 7880 31720 7886
rect 31668 7822 31720 7828
rect 31484 7812 31536 7818
rect 31484 7754 31536 7760
rect 31208 6656 31260 6662
rect 31208 6598 31260 6604
rect 31392 6656 31444 6662
rect 31392 6598 31444 6604
rect 30196 6316 30248 6322
rect 30196 6258 30248 6264
rect 30288 6316 30340 6322
rect 30288 6258 30340 6264
rect 30564 6316 30616 6322
rect 30564 6258 30616 6264
rect 30656 6316 30708 6322
rect 30656 6258 30708 6264
rect 30104 6112 30156 6118
rect 30104 6054 30156 6060
rect 30116 5778 30144 6054
rect 30104 5772 30156 5778
rect 30104 5714 30156 5720
rect 30208 5710 30236 6258
rect 30288 5908 30340 5914
rect 30288 5850 30340 5856
rect 30196 5704 30248 5710
rect 29918 5672 29974 5681
rect 30196 5646 30248 5652
rect 29918 5607 29974 5616
rect 30208 5234 30236 5646
rect 30300 5234 30328 5850
rect 30576 5556 30604 6258
rect 30656 5704 30708 5710
rect 30654 5672 30656 5681
rect 30708 5672 30710 5681
rect 30654 5607 30710 5616
rect 30656 5568 30708 5574
rect 30576 5528 30656 5556
rect 30576 5370 30604 5528
rect 30656 5510 30708 5516
rect 30932 5568 30984 5574
rect 30932 5510 30984 5516
rect 30564 5364 30616 5370
rect 30564 5306 30616 5312
rect 30196 5228 30248 5234
rect 30196 5170 30248 5176
rect 30288 5228 30340 5234
rect 30288 5170 30340 5176
rect 29644 5160 29696 5166
rect 29642 5128 29644 5137
rect 29696 5128 29698 5137
rect 29642 5063 29698 5072
rect 30840 5024 30892 5030
rect 30840 4966 30892 4972
rect 30852 3466 30880 4966
rect 30944 4622 30972 5510
rect 31220 4690 31248 6598
rect 31496 6254 31524 7754
rect 31680 7546 31708 7822
rect 31668 7540 31720 7546
rect 31668 7482 31720 7488
rect 31484 6248 31536 6254
rect 31484 6190 31536 6196
rect 31496 5642 31524 6190
rect 32140 5710 32168 8434
rect 32416 5710 32444 8910
rect 32508 6798 32536 10202
rect 32876 9654 32904 20266
rect 33324 19372 33376 19378
rect 33324 19314 33376 19320
rect 33336 18970 33364 19314
rect 33324 18964 33376 18970
rect 33324 18906 33376 18912
rect 33428 18358 33456 23054
rect 33520 22778 33548 28970
rect 33784 28552 33836 28558
rect 33784 28494 33836 28500
rect 33796 28082 33824 28494
rect 33784 28076 33836 28082
rect 33784 28018 33836 28024
rect 33692 27328 33744 27334
rect 33692 27270 33744 27276
rect 33704 26382 33732 27270
rect 33796 27130 33824 28018
rect 33888 28014 33916 29174
rect 33876 28008 33928 28014
rect 33876 27950 33928 27956
rect 33784 27124 33836 27130
rect 33784 27066 33836 27072
rect 33968 26784 34020 26790
rect 33968 26726 34020 26732
rect 33692 26376 33744 26382
rect 33692 26318 33744 26324
rect 33600 24336 33652 24342
rect 33600 24278 33652 24284
rect 33508 22772 33560 22778
rect 33508 22714 33560 22720
rect 33612 22574 33640 24278
rect 33784 23520 33836 23526
rect 33784 23462 33836 23468
rect 33600 22568 33652 22574
rect 33600 22510 33652 22516
rect 33508 22432 33560 22438
rect 33508 22374 33560 22380
rect 33520 22234 33548 22374
rect 33508 22228 33560 22234
rect 33508 22170 33560 22176
rect 33796 21554 33824 23462
rect 33784 21548 33836 21554
rect 33784 21490 33836 21496
rect 33692 21480 33744 21486
rect 33692 21422 33744 21428
rect 33600 20256 33652 20262
rect 33600 20198 33652 20204
rect 33612 19378 33640 20198
rect 33600 19372 33652 19378
rect 33600 19314 33652 19320
rect 33416 18352 33468 18358
rect 33416 18294 33468 18300
rect 33416 17536 33468 17542
rect 33416 17478 33468 17484
rect 33428 16522 33456 17478
rect 33508 17332 33560 17338
rect 33508 17274 33560 17280
rect 33416 16516 33468 16522
rect 33416 16458 33468 16464
rect 33048 15496 33100 15502
rect 33048 15438 33100 15444
rect 32956 13252 33008 13258
rect 32956 13194 33008 13200
rect 32968 12986 32996 13194
rect 32956 12980 33008 12986
rect 32956 12922 33008 12928
rect 33060 11762 33088 15438
rect 32956 11756 33008 11762
rect 32956 11698 33008 11704
rect 33048 11756 33100 11762
rect 33048 11698 33100 11704
rect 32864 9648 32916 9654
rect 32864 9590 32916 9596
rect 32680 9376 32732 9382
rect 32680 9318 32732 9324
rect 32588 9036 32640 9042
rect 32588 8978 32640 8984
rect 32600 8498 32628 8978
rect 32588 8492 32640 8498
rect 32588 8434 32640 8440
rect 32692 6798 32720 9318
rect 32968 8974 32996 11698
rect 33060 11354 33088 11698
rect 33048 11348 33100 11354
rect 33048 11290 33100 11296
rect 33520 9178 33548 17274
rect 33600 17128 33652 17134
rect 33600 17070 33652 17076
rect 33612 16590 33640 17070
rect 33600 16584 33652 16590
rect 33600 16526 33652 16532
rect 33612 16250 33640 16526
rect 33600 16244 33652 16250
rect 33600 16186 33652 16192
rect 33600 15496 33652 15502
rect 33600 15438 33652 15444
rect 33612 15026 33640 15438
rect 33600 15020 33652 15026
rect 33600 14962 33652 14968
rect 33612 13870 33640 14962
rect 33600 13864 33652 13870
rect 33600 13806 33652 13812
rect 33508 9172 33560 9178
rect 33508 9114 33560 9120
rect 32956 8968 33008 8974
rect 32956 8910 33008 8916
rect 33704 8634 33732 21422
rect 33876 20800 33928 20806
rect 33876 20742 33928 20748
rect 33888 9110 33916 20742
rect 33980 16998 34008 26726
rect 34072 22794 34100 30806
rect 34164 26994 34192 32778
rect 34256 30122 34284 34546
rect 34612 33992 34664 33998
rect 34612 33934 34664 33940
rect 34428 33924 34480 33930
rect 34428 33866 34480 33872
rect 34440 33658 34468 33866
rect 34428 33652 34480 33658
rect 34428 33594 34480 33600
rect 34244 30116 34296 30122
rect 34244 30058 34296 30064
rect 34256 29102 34284 30058
rect 34440 29646 34468 33594
rect 34624 32774 34652 33934
rect 34612 32768 34664 32774
rect 34612 32710 34664 32716
rect 34428 29640 34480 29646
rect 34428 29582 34480 29588
rect 34336 29504 34388 29510
rect 34336 29446 34388 29452
rect 34244 29096 34296 29102
rect 34244 29038 34296 29044
rect 34244 28960 34296 28966
rect 34244 28902 34296 28908
rect 34152 26988 34204 26994
rect 34152 26930 34204 26936
rect 34256 26314 34284 28902
rect 34244 26308 34296 26314
rect 34244 26250 34296 26256
rect 34244 23316 34296 23322
rect 34244 23258 34296 23264
rect 34072 22766 34192 22794
rect 34060 22636 34112 22642
rect 34060 22578 34112 22584
rect 34072 17610 34100 22578
rect 34164 22094 34192 22766
rect 34256 22642 34284 23258
rect 34244 22636 34296 22642
rect 34244 22578 34296 22584
rect 34164 22066 34284 22094
rect 34256 22030 34284 22066
rect 34244 22024 34296 22030
rect 34244 21966 34296 21972
rect 34348 21622 34376 29446
rect 34624 29238 34652 32710
rect 34716 31754 34744 35974
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34796 34468 34848 34474
rect 34796 34410 34848 34416
rect 34808 34202 34836 34410
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34796 34196 34848 34202
rect 34796 34138 34848 34144
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34716 31726 34836 31754
rect 34612 29232 34664 29238
rect 34612 29174 34664 29180
rect 34520 29164 34572 29170
rect 34520 29106 34572 29112
rect 34428 28484 34480 28490
rect 34428 28426 34480 28432
rect 34440 28218 34468 28426
rect 34428 28212 34480 28218
rect 34428 28154 34480 28160
rect 34532 27690 34560 29106
rect 34704 28416 34756 28422
rect 34704 28358 34756 28364
rect 34532 27662 34652 27690
rect 34624 27402 34652 27662
rect 34612 27396 34664 27402
rect 34612 27338 34664 27344
rect 34520 27056 34572 27062
rect 34520 26998 34572 27004
rect 34532 26042 34560 26998
rect 34624 26994 34652 27338
rect 34612 26988 34664 26994
rect 34612 26930 34664 26936
rect 34520 26036 34572 26042
rect 34520 25978 34572 25984
rect 34520 22976 34572 22982
rect 34520 22918 34572 22924
rect 34428 22432 34480 22438
rect 34428 22374 34480 22380
rect 34440 21962 34468 22374
rect 34532 22098 34560 22918
rect 34612 22568 34664 22574
rect 34612 22510 34664 22516
rect 34520 22092 34572 22098
rect 34520 22034 34572 22040
rect 34428 21956 34480 21962
rect 34428 21898 34480 21904
rect 34336 21616 34388 21622
rect 34336 21558 34388 21564
rect 34520 19712 34572 19718
rect 34520 19654 34572 19660
rect 34428 19440 34480 19446
rect 34428 19382 34480 19388
rect 34440 18970 34468 19382
rect 34428 18964 34480 18970
rect 34428 18906 34480 18912
rect 34532 18902 34560 19654
rect 34520 18896 34572 18902
rect 34520 18838 34572 18844
rect 34428 18352 34480 18358
rect 34428 18294 34480 18300
rect 34060 17604 34112 17610
rect 34060 17546 34112 17552
rect 33968 16992 34020 16998
rect 33968 16934 34020 16940
rect 34072 16794 34100 17546
rect 34440 17270 34468 18294
rect 34624 17338 34652 22510
rect 34716 21690 34744 28358
rect 34808 28082 34836 31726
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35348 30728 35400 30734
rect 35348 30670 35400 30676
rect 35164 30660 35216 30666
rect 35164 30602 35216 30608
rect 35176 30190 35204 30602
rect 35164 30184 35216 30190
rect 35164 30126 35216 30132
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35360 29714 35388 30670
rect 35348 29708 35400 29714
rect 35348 29650 35400 29656
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35452 28558 35480 36042
rect 35532 30252 35584 30258
rect 35532 30194 35584 30200
rect 35544 29850 35572 30194
rect 35532 29844 35584 29850
rect 35532 29786 35584 29792
rect 35544 29306 35572 29786
rect 35532 29300 35584 29306
rect 35532 29242 35584 29248
rect 35532 28688 35584 28694
rect 35636 28676 35664 37198
rect 35584 28648 35664 28676
rect 35532 28630 35584 28636
rect 35440 28552 35492 28558
rect 35440 28494 35492 28500
rect 35544 28218 35572 28630
rect 35532 28212 35584 28218
rect 35532 28154 35584 28160
rect 34796 28076 34848 28082
rect 34796 28018 34848 28024
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34796 26784 34848 26790
rect 34796 26726 34848 26732
rect 34808 26382 34836 26726
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34796 26376 34848 26382
rect 34796 26318 34848 26324
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35348 23112 35400 23118
rect 35348 23054 35400 23060
rect 35624 23112 35676 23118
rect 35624 23054 35676 23060
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34704 21684 34756 21690
rect 34704 21626 34756 21632
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35360 20058 35388 23054
rect 35636 22574 35664 23054
rect 35624 22568 35676 22574
rect 35624 22510 35676 22516
rect 35348 20052 35400 20058
rect 35348 19994 35400 20000
rect 35360 19854 35388 19994
rect 35348 19848 35400 19854
rect 35348 19790 35400 19796
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34612 17332 34664 17338
rect 34612 17274 34664 17280
rect 34428 17264 34480 17270
rect 34428 17206 34480 17212
rect 35624 17196 35676 17202
rect 35624 17138 35676 17144
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35636 16794 35664 17138
rect 34060 16788 34112 16794
rect 34060 16730 34112 16736
rect 35624 16788 35676 16794
rect 35624 16730 35676 16736
rect 35348 16040 35400 16046
rect 35348 15982 35400 15988
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34704 15564 34756 15570
rect 34704 15506 34756 15512
rect 34716 14550 34744 15506
rect 35360 14958 35388 15982
rect 35440 15020 35492 15026
rect 35440 14962 35492 14968
rect 35348 14952 35400 14958
rect 35346 14920 35348 14929
rect 35400 14920 35402 14929
rect 35346 14855 35402 14864
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34704 14544 34756 14550
rect 34704 14486 34756 14492
rect 34796 14544 34848 14550
rect 34796 14486 34848 14492
rect 35348 14544 35400 14550
rect 35348 14486 35400 14492
rect 34716 14414 34744 14486
rect 34704 14408 34756 14414
rect 34704 14350 34756 14356
rect 34808 14074 34836 14486
rect 34796 14068 34848 14074
rect 34796 14010 34848 14016
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35360 13326 35388 14486
rect 35452 14346 35480 14962
rect 35532 14408 35584 14414
rect 35532 14350 35584 14356
rect 35440 14340 35492 14346
rect 35440 14282 35492 14288
rect 35348 13320 35400 13326
rect 35348 13262 35400 13268
rect 35256 13184 35308 13190
rect 35256 13126 35308 13132
rect 35268 12918 35296 13126
rect 35360 12986 35388 13262
rect 35348 12980 35400 12986
rect 35348 12922 35400 12928
rect 35256 12912 35308 12918
rect 35256 12854 35308 12860
rect 34612 12708 34664 12714
rect 34612 12650 34664 12656
rect 34520 11552 34572 11558
rect 34520 11494 34572 11500
rect 34532 11354 34560 11494
rect 34520 11348 34572 11354
rect 34520 11290 34572 11296
rect 34520 9444 34572 9450
rect 34520 9386 34572 9392
rect 33876 9104 33928 9110
rect 33876 9046 33928 9052
rect 34532 8634 34560 9386
rect 33692 8628 33744 8634
rect 33692 8570 33744 8576
rect 34520 8628 34572 8634
rect 34520 8570 34572 8576
rect 34624 7546 34652 12650
rect 34704 12640 34756 12646
rect 34704 12582 34756 12588
rect 34716 11898 34744 12582
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34796 12232 34848 12238
rect 34796 12174 34848 12180
rect 34704 11892 34756 11898
rect 34704 11834 34756 11840
rect 34808 10674 34836 12174
rect 35348 12164 35400 12170
rect 35348 12106 35400 12112
rect 35256 12096 35308 12102
rect 35256 12038 35308 12044
rect 35268 11830 35296 12038
rect 35256 11824 35308 11830
rect 35256 11766 35308 11772
rect 35360 11762 35388 12106
rect 35452 11778 35480 14282
rect 35544 13258 35572 14350
rect 35532 13252 35584 13258
rect 35532 13194 35584 13200
rect 35624 13252 35676 13258
rect 35624 13194 35676 13200
rect 35544 12170 35572 13194
rect 35636 12986 35664 13194
rect 35624 12980 35676 12986
rect 35624 12922 35676 12928
rect 35532 12164 35584 12170
rect 35532 12106 35584 12112
rect 35452 11762 35572 11778
rect 35348 11756 35400 11762
rect 35452 11756 35584 11762
rect 35452 11750 35532 11756
rect 35348 11698 35400 11704
rect 35532 11698 35584 11704
rect 35624 11756 35676 11762
rect 35624 11698 35676 11704
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35256 11144 35308 11150
rect 35256 11086 35308 11092
rect 35360 11098 35388 11698
rect 35440 11552 35492 11558
rect 35440 11494 35492 11500
rect 35452 11218 35480 11494
rect 35440 11212 35492 11218
rect 35440 11154 35492 11160
rect 34796 10668 34848 10674
rect 34796 10610 34848 10616
rect 34808 9654 34836 10610
rect 35268 10554 35296 11086
rect 35360 11070 35480 11098
rect 35348 11008 35400 11014
rect 35348 10950 35400 10956
rect 35360 10674 35388 10950
rect 35348 10668 35400 10674
rect 35348 10610 35400 10616
rect 35268 10526 35388 10554
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35360 10282 35388 10526
rect 35268 10254 35388 10282
rect 34796 9648 34848 9654
rect 34796 9590 34848 9596
rect 34704 9580 34756 9586
rect 34704 9522 34756 9528
rect 34716 7562 34744 9522
rect 34808 8974 34836 9590
rect 35268 9450 35296 10254
rect 35452 9466 35480 11070
rect 35256 9444 35308 9450
rect 35256 9386 35308 9392
rect 35360 9438 35480 9466
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34796 8968 34848 8974
rect 34796 8910 34848 8916
rect 34980 8900 35032 8906
rect 34980 8842 35032 8848
rect 34992 8634 35020 8842
rect 34980 8628 35032 8634
rect 34980 8570 35032 8576
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35360 7954 35388 9438
rect 35440 9376 35492 9382
rect 35440 9318 35492 9324
rect 35452 8498 35480 9318
rect 35440 8492 35492 8498
rect 35440 8434 35492 8440
rect 35348 7948 35400 7954
rect 35348 7890 35400 7896
rect 35360 7834 35388 7890
rect 35544 7886 35572 11698
rect 35636 9586 35664 11698
rect 35624 9580 35676 9586
rect 35624 9522 35676 9528
rect 35636 9178 35664 9522
rect 35624 9172 35676 9178
rect 35624 9114 35676 9120
rect 35268 7806 35388 7834
rect 35532 7880 35584 7886
rect 35532 7822 35584 7828
rect 35624 7880 35676 7886
rect 35624 7822 35676 7828
rect 34612 7540 34664 7546
rect 34716 7534 34836 7562
rect 34612 7482 34664 7488
rect 34704 7472 34756 7478
rect 34704 7414 34756 7420
rect 32496 6792 32548 6798
rect 32496 6734 32548 6740
rect 32680 6792 32732 6798
rect 32680 6734 32732 6740
rect 34336 6792 34388 6798
rect 34336 6734 34388 6740
rect 32508 6458 32536 6734
rect 32496 6452 32548 6458
rect 32496 6394 32548 6400
rect 32508 5914 32536 6394
rect 34348 6390 34376 6734
rect 34336 6384 34388 6390
rect 34336 6326 34388 6332
rect 32496 5908 32548 5914
rect 32496 5850 32548 5856
rect 34716 5846 34744 7414
rect 34808 7410 34836 7534
rect 35268 7410 35296 7806
rect 35544 7478 35572 7822
rect 35636 7546 35664 7822
rect 35624 7540 35676 7546
rect 35624 7482 35676 7488
rect 35532 7472 35584 7478
rect 35532 7414 35584 7420
rect 34796 7404 34848 7410
rect 34796 7346 34848 7352
rect 35256 7404 35308 7410
rect 35256 7346 35308 7352
rect 34808 6254 34836 7346
rect 35348 7268 35400 7274
rect 35348 7210 35400 7216
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35360 6322 35388 7210
rect 35532 6792 35584 6798
rect 35532 6734 35584 6740
rect 35440 6656 35492 6662
rect 35440 6598 35492 6604
rect 35348 6316 35400 6322
rect 35348 6258 35400 6264
rect 34796 6248 34848 6254
rect 34796 6190 34848 6196
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34704 5840 34756 5846
rect 34704 5782 34756 5788
rect 32128 5704 32180 5710
rect 32128 5646 32180 5652
rect 32404 5704 32456 5710
rect 32404 5646 32456 5652
rect 31484 5636 31536 5642
rect 31484 5578 31536 5584
rect 31208 4684 31260 4690
rect 31208 4626 31260 4632
rect 30932 4616 30984 4622
rect 30932 4558 30984 4564
rect 31220 3466 31248 4626
rect 32140 3738 32168 5646
rect 32416 4826 32444 5646
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 32404 4820 32456 4826
rect 32404 4762 32456 4768
rect 35452 4146 35480 6598
rect 35544 6458 35572 6734
rect 35532 6452 35584 6458
rect 35532 6394 35584 6400
rect 35440 4140 35492 4146
rect 35440 4082 35492 4088
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 32128 3732 32180 3738
rect 32128 3674 32180 3680
rect 34704 3528 34756 3534
rect 34704 3470 34756 3476
rect 35348 3528 35400 3534
rect 35348 3470 35400 3476
rect 30840 3460 30892 3466
rect 30840 3402 30892 3408
rect 31208 3460 31260 3466
rect 31208 3402 31260 3408
rect 32772 2984 32824 2990
rect 32772 2926 32824 2932
rect 29736 2848 29788 2854
rect 29736 2790 29788 2796
rect 30012 2848 30064 2854
rect 30012 2790 30064 2796
rect 30564 2848 30616 2854
rect 30564 2790 30616 2796
rect 31668 2848 31720 2854
rect 31668 2790 31720 2796
rect 32220 2848 32272 2854
rect 32220 2790 32272 2796
rect 29552 1964 29604 1970
rect 29552 1906 29604 1912
rect 29748 800 29776 2790
rect 30024 800 30052 2790
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 30300 800 30328 2382
rect 30576 800 30604 2790
rect 30840 2440 30892 2446
rect 30840 2382 30892 2388
rect 31116 2440 31168 2446
rect 31116 2382 31168 2388
rect 31392 2440 31444 2446
rect 31392 2382 31444 2388
rect 30852 800 30880 2382
rect 31128 800 31156 2382
rect 31404 800 31432 2382
rect 31680 800 31708 2790
rect 31944 2508 31996 2514
rect 31944 2450 31996 2456
rect 31956 800 31984 2450
rect 32232 800 32260 2790
rect 32496 2440 32548 2446
rect 32496 2382 32548 2388
rect 32508 800 32536 2382
rect 32784 800 32812 2926
rect 33876 2916 33928 2922
rect 33876 2858 33928 2864
rect 33324 2848 33376 2854
rect 33324 2790 33376 2796
rect 33048 2508 33100 2514
rect 33048 2450 33100 2456
rect 33060 800 33088 2450
rect 33336 800 33364 2790
rect 33600 2440 33652 2446
rect 33600 2382 33652 2388
rect 33612 800 33640 2382
rect 33888 800 33916 2858
rect 34428 2848 34480 2854
rect 34428 2790 34480 2796
rect 34152 2576 34204 2582
rect 34152 2518 34204 2524
rect 34164 800 34192 2518
rect 34440 800 34468 2790
rect 34716 800 34744 3470
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35360 1850 35388 3470
rect 35440 2848 35492 2854
rect 35440 2790 35492 2796
rect 34992 1822 35388 1850
rect 34992 800 35020 1822
rect 35452 1442 35480 2790
rect 35532 2508 35584 2514
rect 35532 2450 35584 2456
rect 35268 1414 35480 1442
rect 35268 800 35296 1414
rect 35544 800 35572 2450
rect 35728 2310 35756 56306
rect 40788 56302 40816 56646
rect 43812 56364 43864 56370
rect 43812 56306 43864 56312
rect 40776 56296 40828 56302
rect 40776 56238 40828 56244
rect 43824 37913 43852 56306
rect 44100 56234 44128 57394
rect 44192 56506 44220 57394
rect 47596 56506 47624 57394
rect 54956 57390 54984 59200
rect 56520 57882 56548 59200
rect 57518 57896 57574 57905
rect 56520 57854 56640 57882
rect 56612 57458 56640 57854
rect 57518 57831 57574 57840
rect 56600 57452 56652 57458
rect 56600 57394 56652 57400
rect 54944 57384 54996 57390
rect 54944 57326 54996 57332
rect 57532 57050 57560 57831
rect 58084 57458 58112 59200
rect 58438 59191 58494 59200
rect 58072 57452 58124 57458
rect 58072 57394 58124 57400
rect 57520 57044 57572 57050
rect 57520 56986 57572 56992
rect 57888 56840 57940 56846
rect 57888 56782 57940 56788
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 57900 56545 57928 56782
rect 57886 56536 57942 56545
rect 44180 56500 44232 56506
rect 44180 56442 44232 56448
rect 47584 56500 47636 56506
rect 57886 56471 57942 56480
rect 47584 56442 47636 56448
rect 58452 56370 58480 59191
rect 46756 56364 46808 56370
rect 46756 56306 46808 56312
rect 58440 56364 58492 56370
rect 58440 56306 58492 56312
rect 44088 56228 44140 56234
rect 44088 56170 44140 56176
rect 46768 56166 46796 56306
rect 46756 56160 46808 56166
rect 46756 56102 46808 56108
rect 43810 37904 43866 37913
rect 43810 37839 43866 37848
rect 36452 35556 36504 35562
rect 36452 35498 36504 35504
rect 35808 34536 35860 34542
rect 35808 34478 35860 34484
rect 35820 32910 35848 34478
rect 36084 33448 36136 33454
rect 36084 33390 36136 33396
rect 36096 32910 36124 33390
rect 35808 32904 35860 32910
rect 35808 32846 35860 32852
rect 36084 32904 36136 32910
rect 36084 32846 36136 32852
rect 35992 31816 36044 31822
rect 35992 31758 36044 31764
rect 36176 31816 36228 31822
rect 36176 31758 36228 31764
rect 35808 31340 35860 31346
rect 35808 31282 35860 31288
rect 35820 30190 35848 31282
rect 36004 30734 36032 31758
rect 36188 31482 36216 31758
rect 36268 31680 36320 31686
rect 36268 31622 36320 31628
rect 36176 31476 36228 31482
rect 36176 31418 36228 31424
rect 36280 30870 36308 31622
rect 36268 30864 36320 30870
rect 36268 30806 36320 30812
rect 35992 30728 36044 30734
rect 35992 30670 36044 30676
rect 35900 30252 35952 30258
rect 36004 30240 36032 30670
rect 35952 30212 36032 30240
rect 36280 30308 36308 30806
rect 36360 30320 36412 30326
rect 36280 30280 36360 30308
rect 35900 30194 35952 30200
rect 35808 30184 35860 30190
rect 35808 30126 35860 30132
rect 35820 29578 35848 30126
rect 35808 29572 35860 29578
rect 35808 29514 35860 29520
rect 35900 29572 35952 29578
rect 35900 29514 35952 29520
rect 35820 29034 35848 29514
rect 35808 29028 35860 29034
rect 35808 28970 35860 28976
rect 35820 28762 35848 28970
rect 35808 28756 35860 28762
rect 35808 28698 35860 28704
rect 35912 28626 35940 29514
rect 36084 29504 36136 29510
rect 36084 29446 36136 29452
rect 36096 28626 36124 29446
rect 36280 29102 36308 30280
rect 36360 30262 36412 30268
rect 36464 29306 36492 35498
rect 38936 32904 38988 32910
rect 38936 32846 38988 32852
rect 36636 32428 36688 32434
rect 36636 32370 36688 32376
rect 36648 32026 36676 32370
rect 38948 32366 38976 32846
rect 38936 32360 38988 32366
rect 38936 32302 38988 32308
rect 37280 32224 37332 32230
rect 37280 32166 37332 32172
rect 36636 32020 36688 32026
rect 36636 31962 36688 31968
rect 37292 31346 37320 32166
rect 37648 31680 37700 31686
rect 37648 31622 37700 31628
rect 37660 31346 37688 31622
rect 37280 31340 37332 31346
rect 37280 31282 37332 31288
rect 37648 31340 37700 31346
rect 37648 31282 37700 31288
rect 37660 30394 37688 31282
rect 38948 31142 38976 32302
rect 38936 31136 38988 31142
rect 38936 31078 38988 31084
rect 38948 30734 38976 31078
rect 37924 30728 37976 30734
rect 37924 30670 37976 30676
rect 38568 30728 38620 30734
rect 38568 30670 38620 30676
rect 38936 30728 38988 30734
rect 38936 30670 38988 30676
rect 37648 30388 37700 30394
rect 37648 30330 37700 30336
rect 36544 30048 36596 30054
rect 36544 29990 36596 29996
rect 36556 29646 36584 29990
rect 36544 29640 36596 29646
rect 36544 29582 36596 29588
rect 36636 29572 36688 29578
rect 36636 29514 36688 29520
rect 36648 29306 36676 29514
rect 36452 29300 36504 29306
rect 36452 29242 36504 29248
rect 36636 29300 36688 29306
rect 36636 29242 36688 29248
rect 36268 29096 36320 29102
rect 36268 29038 36320 29044
rect 36280 28694 36308 29038
rect 36268 28688 36320 28694
rect 36188 28648 36268 28676
rect 35900 28620 35952 28626
rect 35900 28562 35952 28568
rect 36084 28620 36136 28626
rect 36084 28562 36136 28568
rect 35992 28552 36044 28558
rect 35992 28494 36044 28500
rect 36004 28082 36032 28494
rect 36188 28150 36216 28648
rect 36268 28630 36320 28636
rect 36464 28558 36492 29242
rect 36452 28552 36504 28558
rect 36452 28494 36504 28500
rect 37280 28484 37332 28490
rect 37280 28426 37332 28432
rect 36176 28144 36228 28150
rect 36176 28086 36228 28092
rect 35992 28076 36044 28082
rect 35992 28018 36044 28024
rect 36004 26450 36032 28018
rect 37292 27946 37320 28426
rect 37464 28416 37516 28422
rect 37464 28358 37516 28364
rect 37476 28014 37504 28358
rect 37464 28008 37516 28014
rect 37464 27950 37516 27956
rect 37280 27940 37332 27946
rect 37280 27882 37332 27888
rect 36268 26784 36320 26790
rect 36268 26726 36320 26732
rect 35992 26444 36044 26450
rect 35992 26386 36044 26392
rect 36084 26308 36136 26314
rect 36084 26250 36136 26256
rect 36096 25974 36124 26250
rect 36084 25968 36136 25974
rect 36084 25910 36136 25916
rect 35992 25152 36044 25158
rect 35992 25094 36044 25100
rect 36004 24206 36032 25094
rect 35992 24200 36044 24206
rect 35992 24142 36044 24148
rect 35900 23724 35952 23730
rect 35900 23666 35952 23672
rect 35912 23186 35940 23666
rect 35900 23180 35952 23186
rect 35900 23122 35952 23128
rect 35912 22642 35940 23122
rect 36004 23118 36032 24142
rect 36176 23724 36228 23730
rect 36176 23666 36228 23672
rect 35992 23112 36044 23118
rect 35992 23054 36044 23060
rect 36188 22642 36216 23666
rect 36280 22642 36308 26726
rect 37556 26308 37608 26314
rect 37556 26250 37608 26256
rect 36360 25832 36412 25838
rect 36360 25774 36412 25780
rect 36372 25294 36400 25774
rect 36360 25288 36412 25294
rect 36360 25230 36412 25236
rect 37280 25220 37332 25226
rect 37280 25162 37332 25168
rect 37292 24410 37320 25162
rect 37372 24608 37424 24614
rect 37372 24550 37424 24556
rect 37280 24404 37332 24410
rect 37280 24346 37332 24352
rect 37384 24206 37412 24550
rect 37372 24200 37424 24206
rect 37372 24142 37424 24148
rect 36360 23724 36412 23730
rect 36360 23666 36412 23672
rect 36372 23322 36400 23666
rect 37188 23588 37240 23594
rect 37188 23530 37240 23536
rect 37200 23322 37228 23530
rect 36360 23316 36412 23322
rect 36360 23258 36412 23264
rect 37188 23316 37240 23322
rect 37188 23258 37240 23264
rect 36372 22982 36400 23258
rect 37280 23044 37332 23050
rect 37280 22986 37332 22992
rect 36360 22976 36412 22982
rect 36360 22918 36412 22924
rect 37292 22778 37320 22986
rect 37280 22772 37332 22778
rect 37280 22714 37332 22720
rect 37384 22642 37412 24142
rect 37568 24070 37596 26250
rect 37660 25498 37688 30330
rect 37936 30122 37964 30670
rect 37924 30116 37976 30122
rect 37924 30058 37976 30064
rect 37936 29714 37964 30058
rect 37924 29708 37976 29714
rect 37924 29650 37976 29656
rect 37936 29102 37964 29650
rect 38580 29238 38608 30670
rect 38568 29232 38620 29238
rect 38568 29174 38620 29180
rect 38752 29232 38804 29238
rect 38752 29174 38804 29180
rect 38016 29164 38068 29170
rect 38016 29106 38068 29112
rect 37924 29096 37976 29102
rect 37924 29038 37976 29044
rect 38028 28762 38056 29106
rect 38016 28756 38068 28762
rect 38016 28698 38068 28704
rect 38764 28082 38792 29174
rect 38752 28076 38804 28082
rect 38752 28018 38804 28024
rect 40592 26988 40644 26994
rect 40592 26930 40644 26936
rect 38752 26784 38804 26790
rect 38752 26726 38804 26732
rect 39948 26784 40000 26790
rect 39948 26726 40000 26732
rect 38764 26382 38792 26726
rect 38752 26376 38804 26382
rect 38752 26318 38804 26324
rect 39960 26042 39988 26726
rect 40408 26240 40460 26246
rect 40408 26182 40460 26188
rect 40500 26240 40552 26246
rect 40500 26182 40552 26188
rect 39948 26036 40000 26042
rect 39948 25978 40000 25984
rect 40420 25974 40448 26182
rect 38660 25968 38712 25974
rect 38660 25910 38712 25916
rect 40408 25968 40460 25974
rect 40408 25910 40460 25916
rect 37648 25492 37700 25498
rect 37648 25434 37700 25440
rect 38292 25492 38344 25498
rect 38292 25434 38344 25440
rect 38304 24886 38332 25434
rect 38672 25294 38700 25910
rect 40040 25900 40092 25906
rect 40040 25842 40092 25848
rect 38844 25696 38896 25702
rect 38844 25638 38896 25644
rect 38660 25288 38712 25294
rect 38660 25230 38712 25236
rect 38292 24880 38344 24886
rect 38292 24822 38344 24828
rect 38672 24614 38700 25230
rect 38660 24608 38712 24614
rect 38660 24550 38712 24556
rect 38568 24200 38620 24206
rect 38568 24142 38620 24148
rect 37556 24064 37608 24070
rect 37556 24006 37608 24012
rect 37464 23588 37516 23594
rect 37464 23530 37516 23536
rect 37476 22710 37504 23530
rect 37464 22704 37516 22710
rect 37464 22646 37516 22652
rect 35900 22636 35952 22642
rect 35900 22578 35952 22584
rect 36176 22636 36228 22642
rect 36176 22578 36228 22584
rect 36268 22636 36320 22642
rect 36268 22578 36320 22584
rect 37372 22636 37424 22642
rect 37372 22578 37424 22584
rect 36188 20448 36216 22578
rect 36636 22568 36688 22574
rect 36636 22510 36688 22516
rect 36648 21894 36676 22510
rect 37384 22234 37412 22578
rect 37372 22228 37424 22234
rect 37372 22170 37424 22176
rect 36636 21888 36688 21894
rect 36636 21830 36688 21836
rect 36268 20460 36320 20466
rect 36188 20420 36268 20448
rect 36268 20402 36320 20408
rect 36084 20052 36136 20058
rect 36084 19994 36136 20000
rect 36096 19378 36124 19994
rect 36280 19786 36308 20402
rect 36268 19780 36320 19786
rect 36268 19722 36320 19728
rect 36280 19446 36308 19722
rect 36268 19440 36320 19446
rect 36268 19382 36320 19388
rect 35900 19372 35952 19378
rect 35900 19314 35952 19320
rect 36084 19372 36136 19378
rect 36084 19314 36136 19320
rect 35912 17746 35940 19314
rect 36452 18284 36504 18290
rect 36452 18226 36504 18232
rect 35900 17740 35952 17746
rect 35900 17682 35952 17688
rect 36360 17604 36412 17610
rect 36360 17546 36412 17552
rect 36372 17338 36400 17546
rect 36360 17332 36412 17338
rect 36360 17274 36412 17280
rect 36084 17196 36136 17202
rect 35912 17156 36084 17184
rect 35912 16454 35940 17156
rect 36084 17138 36136 17144
rect 36268 16788 36320 16794
rect 36268 16730 36320 16736
rect 35900 16448 35952 16454
rect 35900 16390 35952 16396
rect 35808 14952 35860 14958
rect 35808 14894 35860 14900
rect 35820 14482 35848 14894
rect 35808 14476 35860 14482
rect 35808 14418 35860 14424
rect 35912 12850 35940 16390
rect 36280 15026 36308 16730
rect 36268 15020 36320 15026
rect 36268 14962 36320 14968
rect 36464 14006 36492 18226
rect 36452 14000 36504 14006
rect 36452 13942 36504 13948
rect 36268 13932 36320 13938
rect 36268 13874 36320 13880
rect 36084 13728 36136 13734
rect 36084 13670 36136 13676
rect 36096 12850 36124 13670
rect 36280 12850 36308 13874
rect 36464 13190 36492 13942
rect 36452 13184 36504 13190
rect 36452 13126 36504 13132
rect 35900 12844 35952 12850
rect 35900 12786 35952 12792
rect 36084 12844 36136 12850
rect 36084 12786 36136 12792
rect 36268 12844 36320 12850
rect 36268 12786 36320 12792
rect 35912 12102 35940 12786
rect 35900 12096 35952 12102
rect 35900 12038 35952 12044
rect 35808 9036 35860 9042
rect 35808 8978 35860 8984
rect 35820 8566 35848 8978
rect 36280 8974 36308 12786
rect 36544 11892 36596 11898
rect 36544 11834 36596 11840
rect 36556 11150 36584 11834
rect 36648 11830 36676 21830
rect 37568 20942 37596 24006
rect 38580 23594 38608 24142
rect 38672 23798 38700 24550
rect 38752 24268 38804 24274
rect 38752 24210 38804 24216
rect 38764 23866 38792 24210
rect 38752 23860 38804 23866
rect 38752 23802 38804 23808
rect 38660 23792 38712 23798
rect 38660 23734 38712 23740
rect 38568 23588 38620 23594
rect 38568 23530 38620 23536
rect 37740 23520 37792 23526
rect 37740 23462 37792 23468
rect 37752 22642 37780 23462
rect 38672 23118 38700 23734
rect 38660 23112 38712 23118
rect 38660 23054 38712 23060
rect 37740 22636 37792 22642
rect 37740 22578 37792 22584
rect 38764 22506 38792 23802
rect 38856 23662 38884 25638
rect 40052 25498 40080 25842
rect 40040 25492 40092 25498
rect 40040 25434 40092 25440
rect 40512 25294 40540 26182
rect 40604 26042 40632 26930
rect 41052 26308 41104 26314
rect 41052 26250 41104 26256
rect 40592 26036 40644 26042
rect 40592 25978 40644 25984
rect 40868 25900 40920 25906
rect 40868 25842 40920 25848
rect 40592 25832 40644 25838
rect 40592 25774 40644 25780
rect 40500 25288 40552 25294
rect 40500 25230 40552 25236
rect 40604 25226 40632 25774
rect 40592 25220 40644 25226
rect 40592 25162 40644 25168
rect 39212 25152 39264 25158
rect 39212 25094 39264 25100
rect 38844 23656 38896 23662
rect 38844 23598 38896 23604
rect 39224 23322 39252 25094
rect 39580 24132 39632 24138
rect 39580 24074 39632 24080
rect 39856 24132 39908 24138
rect 39856 24074 39908 24080
rect 39592 23730 39620 24074
rect 39764 23792 39816 23798
rect 39764 23734 39816 23740
rect 39580 23724 39632 23730
rect 39580 23666 39632 23672
rect 39212 23316 39264 23322
rect 39212 23258 39264 23264
rect 39776 22710 39804 23734
rect 39764 22704 39816 22710
rect 39764 22646 39816 22652
rect 38752 22500 38804 22506
rect 38752 22442 38804 22448
rect 39396 21548 39448 21554
rect 39396 21490 39448 21496
rect 38568 21344 38620 21350
rect 38568 21286 38620 21292
rect 38580 21146 38608 21286
rect 38568 21140 38620 21146
rect 38568 21082 38620 21088
rect 39408 20942 39436 21490
rect 37004 20936 37056 20942
rect 37004 20878 37056 20884
rect 37556 20936 37608 20942
rect 37556 20878 37608 20884
rect 38200 20936 38252 20942
rect 38200 20878 38252 20884
rect 39396 20936 39448 20942
rect 39396 20878 39448 20884
rect 37016 19854 37044 20878
rect 37188 20868 37240 20874
rect 37188 20810 37240 20816
rect 37200 20398 37228 20810
rect 37188 20392 37240 20398
rect 37188 20334 37240 20340
rect 37004 19848 37056 19854
rect 37004 19790 37056 19796
rect 37016 18766 37044 19790
rect 37004 18760 37056 18766
rect 37004 18702 37056 18708
rect 37016 18222 37044 18702
rect 37200 18698 37228 20334
rect 37832 19984 37884 19990
rect 37832 19926 37884 19932
rect 37372 19712 37424 19718
rect 37372 19654 37424 19660
rect 37280 19372 37332 19378
rect 37280 19314 37332 19320
rect 37188 18692 37240 18698
rect 37188 18634 37240 18640
rect 37200 18358 37228 18634
rect 37188 18352 37240 18358
rect 37188 18294 37240 18300
rect 37004 18216 37056 18222
rect 37004 18158 37056 18164
rect 37016 16590 37044 18158
rect 37004 16584 37056 16590
rect 36818 16552 36874 16561
rect 37004 16526 37056 16532
rect 36818 16487 36874 16496
rect 36832 16454 36860 16487
rect 36820 16448 36872 16454
rect 36820 16390 36872 16396
rect 37016 15570 37044 16526
rect 37200 16522 37228 18294
rect 37188 16516 37240 16522
rect 37188 16458 37240 16464
rect 37200 16114 37228 16458
rect 37188 16108 37240 16114
rect 37188 16050 37240 16056
rect 37004 15564 37056 15570
rect 37004 15506 37056 15512
rect 37292 14550 37320 19314
rect 37280 14544 37332 14550
rect 37280 14486 37332 14492
rect 36728 14272 36780 14278
rect 36728 14214 36780 14220
rect 36740 13938 36768 14214
rect 36728 13932 36780 13938
rect 36728 13874 36780 13880
rect 37280 12300 37332 12306
rect 37280 12242 37332 12248
rect 37292 11898 37320 12242
rect 37280 11892 37332 11898
rect 37280 11834 37332 11840
rect 36636 11824 36688 11830
rect 36636 11766 36688 11772
rect 36648 11150 36676 11766
rect 36544 11144 36596 11150
rect 36544 11086 36596 11092
rect 36636 11144 36688 11150
rect 36636 11086 36688 11092
rect 36556 10810 36584 11086
rect 36544 10804 36596 10810
rect 36544 10746 36596 10752
rect 36648 10266 36676 11086
rect 36636 10260 36688 10266
rect 36636 10202 36688 10208
rect 37096 10056 37148 10062
rect 37096 9998 37148 10004
rect 36268 8968 36320 8974
rect 36268 8910 36320 8916
rect 37004 8968 37056 8974
rect 37004 8910 37056 8916
rect 35808 8560 35860 8566
rect 35808 8502 35860 8508
rect 35820 6730 35848 8502
rect 36280 8498 36308 8910
rect 37016 8634 37044 8910
rect 37004 8628 37056 8634
rect 37004 8570 37056 8576
rect 36268 8492 36320 8498
rect 36268 8434 36320 8440
rect 36176 7404 36228 7410
rect 36176 7346 36228 7352
rect 35900 6792 35952 6798
rect 35900 6734 35952 6740
rect 35808 6724 35860 6730
rect 35808 6666 35860 6672
rect 35820 6390 35848 6666
rect 35808 6384 35860 6390
rect 35808 6326 35860 6332
rect 35912 6322 35940 6734
rect 36188 6322 36216 7346
rect 36280 6798 36308 8434
rect 37108 7546 37136 9998
rect 37280 9988 37332 9994
rect 37280 9930 37332 9936
rect 37292 8974 37320 9930
rect 37384 9518 37412 19654
rect 37648 19372 37700 19378
rect 37648 19314 37700 19320
rect 37556 18352 37608 18358
rect 37556 18294 37608 18300
rect 37464 18284 37516 18290
rect 37464 18226 37516 18232
rect 37476 17882 37504 18226
rect 37464 17876 37516 17882
rect 37464 17818 37516 17824
rect 37476 17270 37504 17818
rect 37464 17264 37516 17270
rect 37464 17206 37516 17212
rect 37568 17202 37596 18294
rect 37556 17196 37608 17202
rect 37556 17138 37608 17144
rect 37568 14958 37596 17138
rect 37556 14952 37608 14958
rect 37556 14894 37608 14900
rect 37568 14618 37596 14894
rect 37556 14612 37608 14618
rect 37556 14554 37608 14560
rect 37464 14408 37516 14414
rect 37516 14368 37596 14396
rect 37464 14350 37516 14356
rect 37464 13932 37516 13938
rect 37464 13874 37516 13880
rect 37476 12306 37504 13874
rect 37568 12322 37596 14368
rect 37660 14006 37688 19314
rect 37740 15496 37792 15502
rect 37740 15438 37792 15444
rect 37752 15162 37780 15438
rect 37740 15156 37792 15162
rect 37740 15098 37792 15104
rect 37752 14414 37780 15098
rect 37740 14408 37792 14414
rect 37740 14350 37792 14356
rect 37648 14000 37700 14006
rect 37648 13942 37700 13948
rect 37660 13530 37688 13942
rect 37648 13524 37700 13530
rect 37648 13466 37700 13472
rect 37660 12442 37688 13466
rect 37648 12436 37700 12442
rect 37648 12378 37700 12384
rect 37464 12300 37516 12306
rect 37568 12294 37780 12322
rect 37464 12242 37516 12248
rect 37556 12232 37608 12238
rect 37556 12174 37608 12180
rect 37568 11082 37596 12174
rect 37556 11076 37608 11082
rect 37556 11018 37608 11024
rect 37568 9586 37596 11018
rect 37556 9580 37608 9586
rect 37556 9522 37608 9528
rect 37372 9512 37424 9518
rect 37372 9454 37424 9460
rect 37568 9466 37596 9522
rect 37568 9438 37688 9466
rect 37752 9450 37780 12294
rect 37280 8968 37332 8974
rect 37280 8910 37332 8916
rect 37292 8430 37320 8910
rect 37280 8424 37332 8430
rect 37280 8366 37332 8372
rect 37188 7812 37240 7818
rect 37188 7754 37240 7760
rect 36636 7540 36688 7546
rect 36636 7482 36688 7488
rect 37096 7540 37148 7546
rect 37096 7482 37148 7488
rect 36648 6798 36676 7482
rect 36268 6792 36320 6798
rect 36268 6734 36320 6740
rect 36636 6792 36688 6798
rect 36636 6734 36688 6740
rect 36820 6792 36872 6798
rect 36820 6734 36872 6740
rect 37004 6792 37056 6798
rect 37004 6734 37056 6740
rect 36832 6458 36860 6734
rect 36820 6452 36872 6458
rect 36820 6394 36872 6400
rect 35900 6316 35952 6322
rect 35900 6258 35952 6264
rect 36176 6316 36228 6322
rect 36176 6258 36228 6264
rect 35808 6112 35860 6118
rect 35808 6054 35860 6060
rect 35820 5710 35848 6054
rect 35808 5704 35860 5710
rect 35808 5646 35860 5652
rect 35900 5636 35952 5642
rect 35900 5578 35952 5584
rect 35912 4214 35940 5578
rect 35900 4208 35952 4214
rect 35900 4150 35952 4156
rect 36188 4010 36216 6258
rect 37016 6186 37044 6734
rect 37200 6390 37228 7754
rect 37660 7410 37688 9438
rect 37740 9444 37792 9450
rect 37740 9386 37792 9392
rect 37752 8498 37780 9386
rect 37844 9178 37872 19926
rect 37924 19712 37976 19718
rect 37924 19654 37976 19660
rect 37936 18834 37964 19654
rect 38108 19440 38160 19446
rect 38108 19382 38160 19388
rect 37924 18828 37976 18834
rect 37924 18770 37976 18776
rect 37924 17672 37976 17678
rect 37924 17614 37976 17620
rect 37936 17270 37964 17614
rect 37924 17264 37976 17270
rect 37924 17206 37976 17212
rect 37936 15502 37964 17206
rect 37924 15496 37976 15502
rect 37924 15438 37976 15444
rect 37924 15360 37976 15366
rect 37924 15302 37976 15308
rect 37936 15026 37964 15302
rect 37924 15020 37976 15026
rect 37924 14962 37976 14968
rect 37924 12436 37976 12442
rect 38120 12434 38148 19382
rect 38212 17746 38240 20878
rect 39304 19848 39356 19854
rect 39408 19836 39436 20878
rect 39868 19854 39896 24074
rect 40604 24070 40632 25162
rect 40880 25158 40908 25842
rect 40960 25764 41012 25770
rect 40960 25706 41012 25712
rect 40972 25294 41000 25706
rect 41064 25702 41092 26250
rect 41052 25696 41104 25702
rect 41052 25638 41104 25644
rect 40960 25288 41012 25294
rect 40960 25230 41012 25236
rect 40868 25152 40920 25158
rect 40868 25094 40920 25100
rect 40880 24410 40908 25094
rect 40868 24404 40920 24410
rect 40868 24346 40920 24352
rect 40592 24064 40644 24070
rect 40592 24006 40644 24012
rect 40040 22976 40092 22982
rect 40040 22918 40092 22924
rect 40052 22642 40080 22918
rect 40040 22636 40092 22642
rect 40040 22578 40092 22584
rect 40604 21486 40632 24006
rect 40880 23866 40908 24346
rect 40972 24342 41000 25230
rect 40960 24336 41012 24342
rect 40960 24278 41012 24284
rect 40868 23860 40920 23866
rect 40868 23802 40920 23808
rect 40880 23730 40908 23802
rect 40868 23724 40920 23730
rect 40868 23666 40920 23672
rect 40776 23656 40828 23662
rect 40776 23598 40828 23604
rect 40788 22982 40816 23598
rect 40776 22976 40828 22982
rect 40776 22918 40828 22924
rect 40788 22778 40816 22918
rect 40776 22772 40828 22778
rect 40776 22714 40828 22720
rect 40684 21888 40736 21894
rect 40684 21830 40736 21836
rect 40696 21554 40724 21830
rect 40684 21548 40736 21554
rect 40684 21490 40736 21496
rect 40592 21480 40644 21486
rect 40592 21422 40644 21428
rect 40500 21412 40552 21418
rect 40500 21354 40552 21360
rect 40132 20868 40184 20874
rect 40132 20810 40184 20816
rect 40144 20602 40172 20810
rect 40408 20800 40460 20806
rect 40408 20742 40460 20748
rect 40132 20596 40184 20602
rect 40132 20538 40184 20544
rect 40420 19854 40448 20742
rect 39356 19808 39436 19836
rect 39856 19848 39908 19854
rect 39304 19790 39356 19796
rect 39856 19790 39908 19796
rect 40408 19848 40460 19854
rect 40408 19790 40460 19796
rect 39316 19514 39344 19790
rect 39304 19508 39356 19514
rect 39304 19450 39356 19456
rect 38936 18760 38988 18766
rect 38936 18702 38988 18708
rect 38752 18692 38804 18698
rect 38752 18634 38804 18640
rect 38200 17740 38252 17746
rect 38200 17682 38252 17688
rect 38764 17202 38792 18634
rect 38948 18086 38976 18702
rect 39316 18358 39344 19450
rect 39868 18698 39896 19790
rect 40132 19780 40184 19786
rect 40132 19722 40184 19728
rect 40144 19514 40172 19722
rect 40512 19666 40540 21354
rect 40420 19638 40540 19666
rect 40132 19508 40184 19514
rect 40132 19450 40184 19456
rect 39856 18692 39908 18698
rect 39856 18634 39908 18640
rect 39304 18352 39356 18358
rect 39304 18294 39356 18300
rect 38936 18080 38988 18086
rect 38936 18022 38988 18028
rect 38948 17678 38976 18022
rect 38936 17672 38988 17678
rect 38936 17614 38988 17620
rect 38752 17196 38804 17202
rect 38752 17138 38804 17144
rect 38660 16584 38712 16590
rect 38660 16526 38712 16532
rect 38200 16448 38252 16454
rect 38200 16390 38252 16396
rect 38212 13938 38240 16390
rect 38292 16176 38344 16182
rect 38292 16118 38344 16124
rect 38304 15706 38332 16118
rect 38292 15700 38344 15706
rect 38292 15642 38344 15648
rect 38304 15502 38332 15642
rect 38292 15496 38344 15502
rect 38292 15438 38344 15444
rect 38304 15026 38332 15438
rect 38672 15434 38700 16526
rect 39212 16516 39264 16522
rect 39212 16458 39264 16464
rect 39224 15570 39252 16458
rect 39316 16182 39344 18294
rect 39856 17128 39908 17134
rect 39856 17070 39908 17076
rect 39868 16522 39896 17070
rect 40224 16584 40276 16590
rect 40224 16526 40276 16532
rect 39856 16516 39908 16522
rect 39856 16458 39908 16464
rect 40236 16250 40264 16526
rect 40316 16448 40368 16454
rect 40316 16390 40368 16396
rect 40224 16244 40276 16250
rect 40224 16186 40276 16192
rect 39304 16176 39356 16182
rect 39304 16118 39356 16124
rect 39856 16108 39908 16114
rect 39856 16050 39908 16056
rect 39868 15706 39896 16050
rect 39856 15700 39908 15706
rect 39856 15642 39908 15648
rect 39212 15564 39264 15570
rect 39212 15506 39264 15512
rect 38660 15428 38712 15434
rect 38660 15370 38712 15376
rect 38672 15162 38700 15370
rect 38752 15360 38804 15366
rect 38752 15302 38804 15308
rect 38568 15156 38620 15162
rect 38568 15098 38620 15104
rect 38660 15156 38712 15162
rect 38660 15098 38712 15104
rect 38580 15026 38608 15098
rect 38764 15026 38792 15302
rect 38292 15020 38344 15026
rect 38292 14962 38344 14968
rect 38568 15020 38620 15026
rect 38568 14962 38620 14968
rect 38752 15020 38804 15026
rect 38752 14962 38804 14968
rect 38660 14952 38712 14958
rect 38660 14894 38712 14900
rect 38384 14408 38436 14414
rect 38384 14350 38436 14356
rect 38200 13932 38252 13938
rect 38200 13874 38252 13880
rect 38396 12986 38424 14350
rect 38568 14272 38620 14278
rect 38568 14214 38620 14220
rect 38580 13326 38608 14214
rect 38672 13734 38700 14894
rect 39028 14340 39080 14346
rect 39028 14282 39080 14288
rect 38660 13728 38712 13734
rect 38660 13670 38712 13676
rect 38568 13320 38620 13326
rect 38568 13262 38620 13268
rect 38672 13190 38700 13670
rect 39040 13394 39068 14282
rect 38844 13388 38896 13394
rect 38844 13330 38896 13336
rect 39028 13388 39080 13394
rect 39028 13330 39080 13336
rect 38752 13320 38804 13326
rect 38752 13262 38804 13268
rect 38660 13184 38712 13190
rect 38660 13126 38712 13132
rect 38384 12980 38436 12986
rect 38384 12922 38436 12928
rect 38672 12850 38700 13126
rect 38660 12844 38712 12850
rect 38660 12786 38712 12792
rect 37924 12378 37976 12384
rect 38028 12406 38148 12434
rect 37936 10742 37964 12378
rect 38028 11082 38056 12406
rect 38764 11898 38792 13262
rect 38752 11892 38804 11898
rect 38752 11834 38804 11840
rect 38764 11082 38792 11834
rect 38016 11076 38068 11082
rect 38016 11018 38068 11024
rect 38752 11076 38804 11082
rect 38752 11018 38804 11024
rect 38028 10810 38056 11018
rect 38016 10804 38068 10810
rect 38016 10746 38068 10752
rect 37924 10736 37976 10742
rect 37924 10678 37976 10684
rect 37936 10266 37964 10678
rect 37924 10260 37976 10266
rect 37924 10202 37976 10208
rect 38108 10056 38160 10062
rect 38856 10010 38884 13330
rect 39028 13184 39080 13190
rect 39028 13126 39080 13132
rect 39040 12918 39068 13126
rect 39028 12912 39080 12918
rect 39028 12854 39080 12860
rect 39224 12850 39252 15506
rect 40328 15502 40356 16390
rect 40316 15496 40368 15502
rect 40316 15438 40368 15444
rect 40316 15020 40368 15026
rect 40316 14962 40368 14968
rect 40328 14346 40356 14962
rect 40316 14340 40368 14346
rect 40316 14282 40368 14288
rect 40328 13870 40356 14282
rect 40420 14278 40448 19638
rect 40604 18426 40632 21422
rect 40696 20534 40724 21490
rect 40788 20602 40816 22714
rect 40868 21548 40920 21554
rect 40868 21490 40920 21496
rect 40880 21146 40908 21490
rect 40972 21418 41000 24278
rect 41052 24064 41104 24070
rect 41052 24006 41104 24012
rect 41512 24064 41564 24070
rect 41512 24006 41564 24012
rect 41064 23730 41092 24006
rect 41052 23724 41104 23730
rect 41052 23666 41104 23672
rect 41236 23724 41288 23730
rect 41236 23666 41288 23672
rect 41248 23118 41276 23666
rect 41524 23186 41552 24006
rect 41512 23180 41564 23186
rect 41512 23122 41564 23128
rect 41236 23112 41288 23118
rect 41236 23054 41288 23060
rect 40960 21412 41012 21418
rect 40960 21354 41012 21360
rect 40868 21140 40920 21146
rect 40868 21082 40920 21088
rect 40776 20596 40828 20602
rect 40776 20538 40828 20544
rect 40684 20528 40736 20534
rect 40684 20470 40736 20476
rect 40788 19938 40816 20538
rect 41248 20466 41276 23054
rect 40960 20460 41012 20466
rect 40960 20402 41012 20408
rect 41236 20460 41288 20466
rect 41236 20402 41288 20408
rect 40972 20058 41000 20402
rect 40960 20052 41012 20058
rect 40960 19994 41012 20000
rect 40696 19910 40816 19938
rect 40696 19446 40724 19910
rect 40684 19440 40736 19446
rect 40684 19382 40736 19388
rect 40592 18420 40644 18426
rect 40592 18362 40644 18368
rect 40696 16794 40724 19382
rect 41248 19378 41276 20402
rect 40868 19372 40920 19378
rect 40868 19314 40920 19320
rect 41052 19372 41104 19378
rect 41052 19314 41104 19320
rect 41236 19372 41288 19378
rect 41236 19314 41288 19320
rect 40880 18630 40908 19314
rect 41064 18970 41092 19314
rect 41052 18964 41104 18970
rect 41052 18906 41104 18912
rect 40868 18624 40920 18630
rect 40868 18566 40920 18572
rect 41052 18624 41104 18630
rect 41052 18566 41104 18572
rect 41064 18290 41092 18566
rect 41248 18442 41276 19314
rect 41328 18624 41380 18630
rect 41328 18566 41380 18572
rect 41156 18414 41276 18442
rect 41052 18284 41104 18290
rect 41052 18226 41104 18232
rect 41064 17746 41092 18226
rect 41052 17740 41104 17746
rect 41052 17682 41104 17688
rect 40684 16788 40736 16794
rect 40684 16730 40736 16736
rect 41156 16114 41184 18414
rect 41236 18284 41288 18290
rect 41236 18226 41288 18232
rect 41248 17882 41276 18226
rect 41340 18222 41368 18566
rect 41328 18216 41380 18222
rect 41328 18158 41380 18164
rect 41236 17876 41288 17882
rect 41236 17818 41288 17824
rect 41144 16108 41196 16114
rect 41144 16050 41196 16056
rect 40684 16040 40736 16046
rect 40684 15982 40736 15988
rect 40696 15026 40724 15982
rect 41156 15502 41184 16050
rect 41144 15496 41196 15502
rect 41144 15438 41196 15444
rect 41340 15094 41368 18158
rect 41328 15088 41380 15094
rect 41328 15030 41380 15036
rect 40684 15020 40736 15026
rect 40684 14962 40736 14968
rect 40408 14272 40460 14278
rect 40408 14214 40460 14220
rect 40316 13864 40368 13870
rect 40316 13806 40368 13812
rect 40420 13462 40448 14214
rect 40408 13456 40460 13462
rect 40408 13398 40460 13404
rect 39212 12844 39264 12850
rect 39212 12786 39264 12792
rect 39224 11762 39252 12786
rect 39212 11756 39264 11762
rect 39212 11698 39264 11704
rect 39028 11688 39080 11694
rect 39028 11630 39080 11636
rect 39040 11286 39068 11630
rect 39028 11280 39080 11286
rect 39028 11222 39080 11228
rect 38936 10464 38988 10470
rect 38936 10406 38988 10412
rect 38108 9998 38160 10004
rect 38120 9722 38148 9998
rect 38764 9982 38884 10010
rect 38108 9716 38160 9722
rect 38108 9658 38160 9664
rect 37832 9172 37884 9178
rect 37832 9114 37884 9120
rect 37844 8566 37872 9114
rect 38764 8974 38792 9982
rect 38844 9920 38896 9926
rect 38844 9862 38896 9868
rect 38856 9586 38884 9862
rect 38948 9654 38976 10406
rect 39040 10130 39068 11222
rect 40132 11076 40184 11082
rect 40132 11018 40184 11024
rect 40144 10742 40172 11018
rect 40132 10736 40184 10742
rect 40132 10678 40184 10684
rect 39028 10124 39080 10130
rect 39028 10066 39080 10072
rect 38936 9648 38988 9654
rect 38936 9590 38988 9596
rect 38844 9580 38896 9586
rect 38844 9522 38896 9528
rect 38948 9178 38976 9590
rect 38936 9172 38988 9178
rect 38936 9114 38988 9120
rect 38752 8968 38804 8974
rect 38752 8910 38804 8916
rect 37832 8560 37884 8566
rect 37832 8502 37884 8508
rect 37740 8492 37792 8498
rect 37740 8434 37792 8440
rect 39040 7698 39068 10066
rect 38948 7670 39068 7698
rect 37648 7404 37700 7410
rect 37648 7346 37700 7352
rect 37280 6656 37332 6662
rect 37280 6598 37332 6604
rect 37188 6384 37240 6390
rect 37188 6326 37240 6332
rect 37004 6180 37056 6186
rect 37004 6122 37056 6128
rect 37292 5302 37320 6598
rect 37660 6390 37688 7346
rect 38844 7200 38896 7206
rect 38844 7142 38896 7148
rect 38856 6798 38884 7142
rect 38844 6792 38896 6798
rect 38844 6734 38896 6740
rect 38948 6730 38976 7670
rect 39028 7540 39080 7546
rect 39028 7482 39080 7488
rect 39040 6798 39068 7482
rect 39672 7336 39724 7342
rect 39672 7278 39724 7284
rect 39028 6792 39080 6798
rect 39028 6734 39080 6740
rect 38936 6724 38988 6730
rect 38936 6666 38988 6672
rect 38384 6656 38436 6662
rect 38384 6598 38436 6604
rect 38396 6390 38424 6598
rect 39684 6458 39712 7278
rect 38752 6452 38804 6458
rect 38752 6394 38804 6400
rect 39672 6452 39724 6458
rect 39672 6394 39724 6400
rect 37648 6384 37700 6390
rect 37648 6326 37700 6332
rect 38384 6384 38436 6390
rect 38384 6326 38436 6332
rect 38292 6248 38344 6254
rect 38292 6190 38344 6196
rect 38304 5574 38332 6190
rect 37372 5568 37424 5574
rect 37372 5510 37424 5516
rect 38292 5568 38344 5574
rect 38292 5510 38344 5516
rect 37280 5296 37332 5302
rect 37280 5238 37332 5244
rect 37384 5234 37412 5510
rect 38764 5370 38792 6394
rect 38752 5364 38804 5370
rect 38752 5306 38804 5312
rect 37372 5228 37424 5234
rect 37372 5170 37424 5176
rect 36176 4004 36228 4010
rect 36176 3946 36228 3952
rect 46296 3664 46348 3670
rect 46296 3606 46348 3612
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 36636 3528 36688 3534
rect 36636 3470 36688 3476
rect 37464 3528 37516 3534
rect 37464 3470 37516 3476
rect 38568 3528 38620 3534
rect 38568 3470 38620 3476
rect 39948 3528 40000 3534
rect 39948 3470 40000 3476
rect 40500 3528 40552 3534
rect 40500 3470 40552 3476
rect 41052 3528 41104 3534
rect 41052 3470 41104 3476
rect 42432 3528 42484 3534
rect 42432 3470 42484 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 44364 3528 44416 3534
rect 44364 3470 44416 3476
rect 45192 3528 45244 3534
rect 45192 3470 45244 3476
rect 46020 3528 46072 3534
rect 46020 3470 46072 3476
rect 35716 2304 35768 2310
rect 35716 2246 35768 2252
rect 35820 800 35848 3470
rect 36360 2848 36412 2854
rect 36360 2790 36412 2796
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 36096 800 36124 2382
rect 36372 800 36400 2790
rect 36648 800 36676 3470
rect 37188 2916 37240 2922
rect 37188 2858 37240 2864
rect 36912 2372 36964 2378
rect 36912 2314 36964 2320
rect 36924 800 36952 2314
rect 37200 800 37228 2858
rect 37476 800 37504 3470
rect 38292 2984 38344 2990
rect 38292 2926 38344 2932
rect 37740 2848 37792 2854
rect 37740 2790 37792 2796
rect 37752 800 37780 2790
rect 38016 2576 38068 2582
rect 38016 2518 38068 2524
rect 38028 800 38056 2518
rect 38304 800 38332 2926
rect 38580 800 38608 3470
rect 39120 2916 39172 2922
rect 39120 2858 39172 2864
rect 38844 2508 38896 2514
rect 38844 2450 38896 2456
rect 38856 800 38884 2450
rect 39132 800 39160 2858
rect 39672 2848 39724 2854
rect 39672 2790 39724 2796
rect 39396 2440 39448 2446
rect 39396 2382 39448 2388
rect 39408 800 39436 2382
rect 39684 800 39712 2790
rect 39960 800 39988 3470
rect 40224 2916 40276 2922
rect 40224 2858 40276 2864
rect 40236 800 40264 2858
rect 40512 800 40540 3470
rect 40776 2508 40828 2514
rect 40776 2450 40828 2456
rect 40788 800 40816 2450
rect 41064 800 41092 3470
rect 42156 2984 42208 2990
rect 42156 2926 42208 2932
rect 41604 2848 41656 2854
rect 41604 2790 41656 2796
rect 41328 2440 41380 2446
rect 41328 2382 41380 2388
rect 41340 800 41368 2382
rect 41616 800 41644 2790
rect 41880 2576 41932 2582
rect 41880 2518 41932 2524
rect 41892 800 41920 2518
rect 42168 800 42196 2926
rect 42444 800 42472 3470
rect 42720 800 42748 3470
rect 42984 2916 43036 2922
rect 42984 2858 43036 2864
rect 44088 2916 44140 2922
rect 44088 2858 44140 2864
rect 42996 800 43024 2858
rect 43536 2848 43588 2854
rect 43536 2790 43588 2796
rect 43260 2508 43312 2514
rect 43260 2450 43312 2456
rect 43272 800 43300 2450
rect 43548 800 43576 2790
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 43824 800 43852 2382
rect 44100 800 44128 2858
rect 44376 800 44404 3470
rect 44916 2848 44968 2854
rect 44916 2790 44968 2796
rect 44640 2372 44692 2378
rect 44640 2314 44692 2320
rect 44652 800 44680 2314
rect 44928 800 44956 2790
rect 45204 800 45232 3470
rect 45468 2848 45520 2854
rect 45468 2790 45520 2796
rect 45480 800 45508 2790
rect 45744 2576 45796 2582
rect 45744 2518 45796 2524
rect 45756 800 45784 2518
rect 46032 800 46060 3470
rect 46308 800 46336 3606
rect 46572 2508 46624 2514
rect 46572 2450 46624 2456
rect 46584 800 46612 2450
rect 46768 2310 46796 56102
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 58162 55176 58218 55185
rect 58162 55111 58164 55120
rect 58216 55111 58218 55120
rect 58164 55082 58216 55088
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 57888 53984 57940 53990
rect 57888 53926 57940 53932
rect 57900 53825 57928 53926
rect 57886 53816 57942 53825
rect 57886 53751 57942 53760
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 57888 52488 57940 52494
rect 57886 52456 57888 52465
rect 57940 52456 57942 52465
rect 57886 52391 57942 52400
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 58164 51400 58216 51406
rect 58164 51342 58216 51348
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 58176 51105 58204 51342
rect 58162 51096 58218 51105
rect 58162 51031 58218 51040
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 58164 49768 58216 49774
rect 58162 49736 58164 49745
rect 58216 49736 58218 49745
rect 58162 49671 58218 49680
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 58164 48544 58216 48550
rect 58164 48486 58216 48492
rect 58176 48385 58204 48486
rect 58162 48376 58218 48385
rect 58162 48311 58218 48320
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 58164 47048 58216 47054
rect 58162 47016 58164 47025
rect 58216 47016 58218 47025
rect 58162 46951 58218 46960
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 58164 45960 58216 45966
rect 58164 45902 58216 45908
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 58176 45665 58204 45902
rect 58162 45656 58218 45665
rect 58162 45591 58218 45600
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 58162 44296 58218 44305
rect 58162 44231 58164 44240
rect 58216 44231 58218 44240
rect 58164 44202 58216 44208
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 58164 43104 58216 43110
rect 58164 43046 58216 43052
rect 58176 42945 58204 43046
rect 58162 42936 58218 42945
rect 58162 42871 58218 42880
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 58164 41608 58216 41614
rect 58162 41576 58164 41585
rect 58216 41576 58218 41585
rect 58162 41511 58218 41520
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 58164 40520 58216 40526
rect 58164 40462 58216 40468
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 58176 40225 58204 40462
rect 58162 40216 58218 40225
rect 58162 40151 58218 40160
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 58162 38856 58218 38865
rect 58162 38791 58164 38800
rect 58216 38791 58218 38800
rect 58164 38762 58216 38768
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 58164 37664 58216 37670
rect 58164 37606 58216 37612
rect 58176 37505 58204 37606
rect 58162 37496 58218 37505
rect 58162 37431 58218 37440
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 58164 36168 58216 36174
rect 58162 36136 58164 36145
rect 58216 36136 58218 36145
rect 58162 36071 58218 36080
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 58164 35080 58216 35086
rect 58164 35022 58216 35028
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 58176 34785 58204 35022
rect 58162 34776 58218 34785
rect 58162 34711 58218 34720
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 58162 33416 58218 33425
rect 58162 33351 58164 33360
rect 58216 33351 58218 33360
rect 58164 33322 58216 33328
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 58164 32224 58216 32230
rect 58164 32166 58216 32172
rect 58176 32065 58204 32166
rect 58162 32056 58218 32065
rect 58162 31991 58218 32000
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 58164 30728 58216 30734
rect 58162 30696 58164 30705
rect 58216 30696 58218 30705
rect 58162 30631 58218 30640
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 58164 29640 58216 29646
rect 58164 29582 58216 29588
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 58176 29345 58204 29582
rect 58162 29336 58218 29345
rect 58162 29271 58218 29280
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 58162 27976 58218 27985
rect 58162 27911 58164 27920
rect 58216 27911 58218 27920
rect 58164 27882 58216 27888
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 58164 26784 58216 26790
rect 58164 26726 58216 26732
rect 58176 26625 58204 26726
rect 58162 26616 58218 26625
rect 58162 26551 58218 26560
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 58164 25288 58216 25294
rect 58162 25256 58164 25265
rect 58216 25256 58218 25265
rect 58162 25191 58218 25200
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 58164 24200 58216 24206
rect 58164 24142 58216 24148
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 58176 23905 58204 24142
rect 58162 23896 58218 23905
rect 58162 23831 58218 23840
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 58162 22536 58218 22545
rect 58162 22471 58164 22480
rect 58216 22471 58218 22480
rect 58164 22442 58216 22448
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 58164 21344 58216 21350
rect 58164 21286 58216 21292
rect 58176 21185 58204 21286
rect 58162 21176 58218 21185
rect 58162 21111 58218 21120
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 58164 19848 58216 19854
rect 58162 19816 58164 19825
rect 58216 19816 58218 19825
rect 58162 19751 58218 19760
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 58164 18760 58216 18766
rect 58164 18702 58216 18708
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 58176 18465 58204 18702
rect 58162 18456 58218 18465
rect 58162 18391 58218 18400
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 58162 17096 58218 17105
rect 58162 17031 58164 17040
rect 58216 17031 58218 17040
rect 58164 17002 58216 17008
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 58164 15904 58216 15910
rect 58164 15846 58216 15852
rect 58176 15745 58204 15846
rect 58162 15736 58218 15745
rect 58162 15671 58218 15680
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 58164 14408 58216 14414
rect 58162 14376 58164 14385
rect 58216 14376 58218 14385
rect 58162 14311 58218 14320
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 58164 13320 58216 13326
rect 58164 13262 58216 13268
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 58176 13025 58204 13262
rect 58162 13016 58218 13025
rect 58162 12951 58218 12960
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 58162 11656 58218 11665
rect 58162 11591 58164 11600
rect 58216 11591 58218 11600
rect 58164 11562 58216 11568
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 58164 10464 58216 10470
rect 58164 10406 58216 10412
rect 58176 10305 58204 10406
rect 58162 10296 58218 10305
rect 58162 10231 58218 10240
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 58164 8968 58216 8974
rect 58162 8936 58164 8945
rect 58216 8936 58218 8945
rect 58162 8871 58218 8880
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 58164 7880 58216 7886
rect 58164 7822 58216 7828
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 58176 7585 58204 7822
rect 58162 7576 58218 7585
rect 58162 7511 58218 7520
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 58162 6216 58218 6225
rect 58162 6151 58164 6160
rect 58216 6151 58218 6160
rect 58164 6122 58216 6128
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 53748 5160 53800 5166
rect 53748 5102 53800 5108
rect 53656 5024 53708 5030
rect 53656 4966 53708 4972
rect 52184 4752 52236 4758
rect 52184 4694 52236 4700
rect 52092 4616 52144 4622
rect 52092 4558 52144 4564
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 51816 4072 51868 4078
rect 51816 4014 51868 4020
rect 51080 3936 51132 3942
rect 51080 3878 51132 3884
rect 51356 3936 51408 3942
rect 51356 3878 51408 3884
rect 50804 3596 50856 3602
rect 50804 3538 50856 3544
rect 47676 3528 47728 3534
rect 47676 3470 47728 3476
rect 48228 3528 48280 3534
rect 48228 3470 48280 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50620 3528 50672 3534
rect 50620 3470 50672 3476
rect 47400 2916 47452 2922
rect 47400 2858 47452 2864
rect 46848 2848 46900 2854
rect 46848 2790 46900 2796
rect 46756 2304 46808 2310
rect 46756 2246 46808 2252
rect 46860 800 46888 2790
rect 47124 2440 47176 2446
rect 47124 2382 47176 2388
rect 47136 800 47164 2382
rect 47412 800 47440 2858
rect 47688 800 47716 3470
rect 47952 2848 48004 2854
rect 47952 2790 48004 2796
rect 47964 800 47992 2790
rect 48240 800 48268 3470
rect 48780 2916 48832 2922
rect 48780 2858 48832 2864
rect 49884 2916 49936 2922
rect 49884 2858 49936 2864
rect 48504 2508 48556 2514
rect 48504 2450 48556 2456
rect 48516 800 48544 2450
rect 48792 800 48820 2858
rect 49332 2848 49384 2854
rect 49332 2790 49384 2796
rect 49056 2440 49108 2446
rect 49056 2382 49108 2388
rect 49068 800 49096 2382
rect 49344 800 49372 2790
rect 49608 2576 49660 2582
rect 49608 2518 49660 2524
rect 49620 800 49648 2518
rect 49896 800 49924 2858
rect 50172 800 50200 3470
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50632 1850 50660 3470
rect 50712 2848 50764 2854
rect 50712 2790 50764 2796
rect 50448 1822 50660 1850
rect 50448 800 50476 1822
rect 50724 1442 50752 2790
rect 50632 1414 50752 1442
rect 50632 800 50660 1414
rect 50816 1306 50844 3538
rect 50988 2916 51040 2922
rect 50988 2858 51040 2864
rect 50896 2440 50948 2446
rect 50896 2382 50948 2388
rect 50724 1278 50844 1306
rect 50724 800 50752 1278
rect 50908 1170 50936 2382
rect 50816 1142 50936 1170
rect 50816 800 50844 1142
rect 51000 1034 51028 2858
rect 50908 1006 51028 1034
rect 50908 800 50936 1006
rect 50988 944 51040 950
rect 50988 886 51040 892
rect 51000 800 51028 886
rect 51092 800 51120 3878
rect 51172 3528 51224 3534
rect 51172 3470 51224 3476
rect 51184 800 51212 3470
rect 51264 2304 51316 2310
rect 51264 2246 51316 2252
rect 51276 800 51304 2246
rect 51368 800 51396 3878
rect 51448 3664 51500 3670
rect 51448 3606 51500 3612
rect 51460 800 51488 3606
rect 51632 3596 51684 3602
rect 51632 3538 51684 3544
rect 51540 2848 51592 2854
rect 51540 2790 51592 2796
rect 51552 800 51580 2790
rect 51644 800 51672 3538
rect 51724 3052 51776 3058
rect 51724 2994 51776 3000
rect 51736 800 51764 2994
rect 51828 800 51856 4014
rect 51908 3120 51960 3126
rect 51908 3062 51960 3068
rect 51920 800 51948 3062
rect 52000 2644 52052 2650
rect 52000 2586 52052 2592
rect 52012 800 52040 2586
rect 52104 800 52132 4558
rect 52196 800 52224 4694
rect 53196 4684 53248 4690
rect 53196 4626 53248 4632
rect 52644 4616 52696 4622
rect 52644 4558 52696 4564
rect 52460 3936 52512 3942
rect 52460 3878 52512 3884
rect 52276 3528 52328 3534
rect 52276 3470 52328 3476
rect 52288 800 52316 3470
rect 52368 2100 52420 2106
rect 52368 2042 52420 2048
rect 52380 800 52408 2042
rect 52472 800 52500 3878
rect 52552 2440 52604 2446
rect 52552 2382 52604 2388
rect 52564 1154 52592 2382
rect 52552 1148 52604 1154
rect 52552 1090 52604 1096
rect 52552 944 52604 950
rect 52552 886 52604 892
rect 52564 800 52592 886
rect 52656 800 52684 4558
rect 53012 4140 53064 4146
rect 53012 4082 53064 4088
rect 52828 4004 52880 4010
rect 52828 3946 52880 3952
rect 52736 3732 52788 3738
rect 52736 3674 52788 3680
rect 52748 1426 52776 3674
rect 52736 1420 52788 1426
rect 52736 1362 52788 1368
rect 52840 1170 52868 3946
rect 53024 2774 53052 4082
rect 53104 2984 53156 2990
rect 53104 2926 53156 2932
rect 52748 1142 52868 1170
rect 52932 2746 53052 2774
rect 52748 800 52776 1142
rect 52932 1034 52960 2746
rect 53012 1420 53064 1426
rect 53012 1362 53064 1368
rect 52840 1006 52960 1034
rect 52840 800 52868 1006
rect 52920 944 52972 950
rect 52920 886 52972 892
rect 52932 800 52960 886
rect 53024 800 53052 1362
rect 53116 800 53144 2926
rect 53208 800 53236 4626
rect 53288 3460 53340 3466
rect 53288 3402 53340 3408
rect 53300 800 53328 3402
rect 53378 2952 53434 2961
rect 53378 2887 53434 2896
rect 53392 800 53420 2887
rect 53470 2816 53526 2825
rect 53470 2751 53526 2760
rect 53484 800 53512 2751
rect 53564 2032 53616 2038
rect 53564 1974 53616 1980
rect 53576 800 53604 1974
rect 53668 800 53696 4966
rect 53760 800 53788 5102
rect 54116 5092 54168 5098
rect 54116 5034 54168 5040
rect 53932 4752 53984 4758
rect 53932 4694 53984 4700
rect 53840 3596 53892 3602
rect 53840 3538 53892 3544
rect 53852 800 53880 3538
rect 53944 800 53972 4694
rect 54024 4072 54076 4078
rect 54024 4014 54076 4020
rect 54036 800 54064 4014
rect 54128 800 54156 5034
rect 58164 5024 58216 5030
rect 58164 4966 58216 4972
rect 58176 4865 58204 4966
rect 58162 4856 58218 4865
rect 58162 4791 58218 4800
rect 54300 4684 54352 4690
rect 54300 4626 54352 4632
rect 54208 2916 54260 2922
rect 54208 2858 54260 2864
rect 54220 800 54248 2858
rect 54312 800 54340 4626
rect 55312 3936 55364 3942
rect 55312 3878 55364 3884
rect 58440 3936 58492 3942
rect 58440 3878 58492 3884
rect 54760 3052 54812 3058
rect 54760 2994 54812 3000
rect 54772 882 54800 2994
rect 55324 2825 55352 3878
rect 57520 3528 57572 3534
rect 58164 3528 58216 3534
rect 57520 3470 57572 3476
rect 58162 3496 58164 3505
rect 58216 3496 58218 3505
rect 56600 2984 56652 2990
rect 56598 2952 56600 2961
rect 56652 2952 56654 2961
rect 56598 2887 56654 2896
rect 55310 2816 55366 2825
rect 55310 2751 55366 2760
rect 55956 2440 56008 2446
rect 55956 2382 56008 2388
rect 56600 2440 56652 2446
rect 56600 2382 56652 2388
rect 55968 2106 55996 2382
rect 55956 2100 56008 2106
rect 55956 2042 56008 2048
rect 56612 1426 56640 2382
rect 57532 2145 57560 3470
rect 58162 3431 58218 3440
rect 57888 2508 57940 2514
rect 57888 2450 57940 2456
rect 57518 2136 57574 2145
rect 57518 2071 57574 2080
rect 57900 2038 57928 2450
rect 57888 2032 57940 2038
rect 57888 1974 57940 1980
rect 56600 1420 56652 1426
rect 56600 1362 56652 1368
rect 54760 876 54812 882
rect 54760 818 54812 824
rect 5538 0 5594 800
rect 5630 0 5686 800
rect 5722 0 5778 800
rect 5814 0 5870 800
rect 5906 0 5962 800
rect 5998 0 6054 800
rect 6090 0 6146 800
rect 6182 0 6238 800
rect 6274 0 6330 800
rect 6366 0 6422 800
rect 6458 0 6514 800
rect 6550 0 6606 800
rect 6642 0 6698 800
rect 6734 0 6790 800
rect 6826 0 6882 800
rect 6918 0 6974 800
rect 7010 0 7066 800
rect 7102 0 7158 800
rect 7194 0 7250 800
rect 7286 0 7342 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8298 0 8354 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10506 0 10562 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48778 0 48834 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50066 0 50122 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50342 0 50398 800
rect 50434 0 50490 800
rect 50526 0 50582 800
rect 50618 0 50674 800
rect 50710 0 50766 800
rect 50802 0 50858 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51078 0 51134 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51354 0 51410 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51630 0 51686 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51906 0 51962 800
rect 51998 0 52054 800
rect 52090 0 52146 800
rect 52182 0 52238 800
rect 52274 0 52330 800
rect 52366 0 52422 800
rect 52458 0 52514 800
rect 52550 0 52606 800
rect 52642 0 52698 800
rect 52734 0 52790 800
rect 52826 0 52882 800
rect 52918 0 52974 800
rect 53010 0 53066 800
rect 53102 0 53158 800
rect 53194 0 53250 800
rect 53286 0 53342 800
rect 53378 0 53434 800
rect 53470 0 53526 800
rect 53562 0 53618 800
rect 53654 0 53710 800
rect 53746 0 53802 800
rect 53838 0 53894 800
rect 53930 0 53986 800
rect 54022 0 54078 800
rect 54114 0 54170 800
rect 54206 0 54262 800
rect 54298 0 54354 800
rect 58452 785 58480 3878
rect 58438 776 58494 785
rect 58438 711 58494 720
<< via2 >>
rect 58438 59200 58494 59256
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 1398 56616 1454 56672
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 14186 56108 14188 56128
rect 14188 56108 14240 56128
rect 14240 56108 14242 56128
rect 14186 56072 14242 56108
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 1398 55528 1454 55584
rect 17038 55564 17040 55584
rect 17040 55564 17092 55584
rect 17092 55564 17094 55584
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 1398 54440 1454 54496
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 1398 53352 1454 53408
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 1398 52264 1454 52320
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 1398 51176 1454 51232
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 1398 50088 1454 50144
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 1398 49000 1454 49056
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 1398 47912 1454 47968
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4894 38292 4896 38312
rect 4896 38292 4948 38312
rect 4948 38292 4950 38312
rect 4894 38256 4950 38292
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 6734 38292 6736 38312
rect 6736 38292 6788 38312
rect 6788 38292 6790 38312
rect 6734 38256 6790 38292
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 5630 31592 5686 31648
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4618 19216 4674 19272
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4158 18572 4160 18592
rect 4160 18572 4212 18592
rect 4212 18572 4214 18592
rect 4158 18536 4214 18572
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 2042 8608 2098 8664
rect 1858 5616 1914 5672
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 5538 13812 5540 13832
rect 5540 13812 5592 13832
rect 5592 13812 5594 13832
rect 5538 13776 5594 13812
rect 8298 31476 8354 31512
rect 8298 31456 8300 31476
rect 8300 31456 8352 31476
rect 8352 31456 8354 31476
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 2134 3032 2190 3088
rect 2594 3984 2650 4040
rect 2594 3032 2650 3088
rect 2502 2896 2558 2952
rect 3514 7928 3570 7984
rect 3882 9560 3938 9616
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 3974 7692 3976 7712
rect 3976 7692 4028 7712
rect 4028 7692 4030 7712
rect 3974 7656 4030 7692
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4894 3848 4950 3904
rect 4894 3732 4950 3768
rect 5078 4528 5134 4584
rect 4894 3712 4896 3732
rect 4896 3712 4948 3732
rect 4948 3712 4950 3732
rect 4894 3168 4950 3224
rect 5262 4664 5318 4720
rect 5262 3848 5318 3904
rect 5170 2760 5226 2816
rect 5538 5480 5594 5536
rect 5538 4276 5594 4312
rect 5538 4256 5540 4276
rect 5540 4256 5592 4276
rect 5592 4256 5594 4276
rect 5538 3984 5594 4040
rect 6090 8608 6146 8664
rect 5814 4120 5870 4176
rect 5998 3848 6054 3904
rect 6366 8744 6422 8800
rect 6734 11212 6790 11248
rect 6734 11192 6736 11212
rect 6736 11192 6788 11212
rect 6788 11192 6790 11212
rect 7378 15136 7434 15192
rect 7286 11212 7342 11248
rect 7286 11192 7288 11212
rect 7288 11192 7340 11212
rect 7340 11192 7342 11212
rect 6366 2896 6422 2952
rect 6550 2644 6606 2680
rect 6550 2624 6552 2644
rect 6552 2624 6604 2644
rect 6604 2624 6606 2644
rect 6918 3032 6974 3088
rect 7102 4120 7158 4176
rect 7654 4276 7710 4312
rect 7654 4256 7656 4276
rect 7656 4256 7708 4276
rect 7708 4256 7710 4276
rect 8022 3032 8078 3088
rect 7746 2760 7802 2816
rect 8574 8372 8576 8392
rect 8576 8372 8628 8392
rect 8628 8372 8630 8392
rect 8574 8336 8630 8372
rect 8206 3188 8262 3224
rect 8206 3168 8208 3188
rect 8208 3168 8260 3188
rect 8260 3168 8262 3188
rect 8850 14764 8852 14784
rect 8852 14764 8904 14784
rect 8904 14764 8906 14784
rect 8850 14728 8906 14764
rect 9586 34176 9642 34232
rect 10414 37984 10470 38040
rect 9862 24132 9918 24168
rect 9862 24112 9864 24132
rect 9864 24112 9916 24132
rect 9916 24112 9918 24132
rect 11334 31592 11390 31648
rect 8666 4020 8668 4040
rect 8668 4020 8720 4040
rect 8720 4020 8722 4040
rect 8666 3984 8722 4020
rect 8758 3712 8814 3768
rect 10690 19116 10692 19136
rect 10692 19116 10744 19136
rect 10744 19116 10746 19136
rect 10690 19080 10746 19116
rect 9770 11056 9826 11112
rect 13542 37032 13598 37088
rect 11702 19080 11758 19136
rect 10966 15408 11022 15464
rect 10230 10412 10232 10432
rect 10232 10412 10284 10432
rect 10284 10412 10286 10432
rect 10230 10376 10286 10412
rect 9586 8472 9642 8528
rect 9770 8508 9772 8528
rect 9772 8508 9824 8528
rect 9824 8508 9826 8528
rect 9770 8472 9826 8508
rect 9586 8084 9642 8120
rect 9586 8064 9588 8084
rect 9588 8064 9640 8084
rect 9640 8064 9642 8084
rect 9586 7112 9642 7168
rect 9494 6976 9550 7032
rect 9402 5072 9458 5128
rect 8666 3052 8722 3088
rect 8666 3032 8668 3052
rect 8668 3032 8720 3052
rect 8720 3032 8722 3052
rect 8942 3052 8998 3088
rect 8942 3032 8944 3052
rect 8944 3032 8996 3052
rect 8996 3032 8998 3052
rect 9494 4004 9550 4040
rect 9494 3984 9496 4004
rect 9496 3984 9548 4004
rect 9548 3984 9550 4004
rect 9862 3304 9918 3360
rect 10322 4664 10378 4720
rect 10414 2644 10470 2680
rect 10414 2624 10416 2644
rect 10416 2624 10468 2644
rect 10468 2624 10470 2644
rect 10598 3576 10654 3632
rect 14554 34196 14610 34232
rect 14554 34176 14556 34196
rect 14556 34176 14608 34196
rect 14608 34176 14610 34196
rect 11886 9288 11942 9344
rect 11794 9016 11850 9072
rect 12254 8492 12310 8528
rect 12254 8472 12256 8492
rect 12256 8472 12308 8492
rect 12308 8472 12310 8492
rect 10966 2896 11022 2952
rect 12438 8200 12494 8256
rect 11518 3984 11574 4040
rect 12254 4684 12310 4720
rect 12254 4664 12256 4684
rect 12256 4664 12308 4684
rect 12308 4664 12310 4684
rect 13358 8628 13414 8664
rect 13358 8608 13360 8628
rect 13360 8608 13412 8628
rect 13412 8608 13414 8628
rect 14830 19796 14832 19816
rect 14832 19796 14884 19816
rect 14884 19796 14886 19816
rect 14830 19760 14886 19796
rect 14094 3168 14150 3224
rect 14738 8336 14794 8392
rect 14554 3188 14610 3224
rect 14554 3168 14556 3188
rect 14556 3168 14608 3188
rect 14608 3168 14610 3188
rect 14554 2644 14610 2680
rect 14554 2624 14556 2644
rect 14556 2624 14608 2644
rect 14608 2624 14610 2644
rect 15566 9288 15622 9344
rect 15198 3188 15254 3224
rect 15198 3168 15200 3188
rect 15200 3168 15252 3188
rect 15252 3168 15254 3188
rect 15566 3032 15622 3088
rect 15842 4004 15898 4040
rect 15842 3984 15844 4004
rect 15844 3984 15896 4004
rect 15896 3984 15898 4004
rect 16118 3188 16174 3224
rect 16118 3168 16120 3188
rect 16120 3168 16172 3188
rect 16172 3168 16174 3188
rect 17038 55528 17094 55564
rect 17682 55528 17738 55584
rect 17774 55292 17776 55312
rect 17776 55292 17828 55312
rect 17828 55292 17830 55312
rect 17774 55256 17830 55292
rect 16762 37984 16818 38040
rect 17866 37032 17922 37088
rect 16854 31476 16910 31512
rect 16854 31456 16856 31476
rect 16856 31456 16908 31476
rect 16908 31456 16910 31476
rect 16762 26324 16764 26344
rect 16764 26324 16816 26344
rect 16816 26324 16818 26344
rect 16762 26288 16818 26324
rect 16670 24148 16672 24168
rect 16672 24148 16724 24168
rect 16724 24148 16726 24168
rect 16670 24112 16726 24148
rect 17038 26288 17094 26344
rect 16578 9016 16634 9072
rect 17222 26444 17278 26480
rect 17222 26424 17224 26444
rect 17224 26424 17276 26444
rect 17276 26424 17278 26444
rect 17958 32428 18014 32464
rect 17958 32408 17960 32428
rect 17960 32408 18012 32428
rect 18012 32408 18014 32428
rect 17682 20460 17738 20496
rect 17682 20440 17684 20460
rect 17684 20440 17736 20460
rect 17736 20440 17738 20460
rect 18786 55292 18788 55312
rect 18788 55292 18840 55312
rect 18840 55292 18842 55312
rect 18786 55256 18842 55292
rect 18510 23704 18566 23760
rect 17314 5616 17370 5672
rect 17406 3188 17462 3224
rect 17406 3168 17408 3188
rect 17408 3168 17460 3188
rect 17460 3168 17462 3188
rect 17498 2524 17500 2544
rect 17500 2524 17552 2544
rect 17552 2524 17554 2544
rect 17498 2488 17554 2524
rect 17682 2624 17738 2680
rect 18878 26444 18934 26480
rect 18878 26424 18880 26444
rect 18880 26424 18932 26444
rect 18932 26424 18934 26444
rect 20166 56788 20168 56808
rect 20168 56788 20220 56808
rect 20220 56788 20222 56808
rect 20166 56752 20222 56788
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 19798 55292 19800 55312
rect 19800 55292 19852 55312
rect 19852 55292 19854 55312
rect 19798 55256 19854 55292
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19982 41656 20038 41712
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19246 19896 19302 19952
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 20258 55564 20260 55584
rect 20260 55564 20312 55584
rect 20312 55564 20314 55584
rect 20258 55528 20314 55564
rect 21730 55564 21732 55584
rect 21732 55564 21784 55584
rect 21784 55564 21786 55584
rect 21730 55528 21786 55564
rect 23018 55564 23020 55584
rect 23020 55564 23072 55584
rect 23072 55564 23074 55584
rect 23018 55528 23074 55564
rect 23754 55564 23756 55584
rect 23756 55564 23808 55584
rect 23808 55564 23810 55584
rect 23754 55528 23810 55564
rect 20166 29824 20222 29880
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19890 29144 19946 29200
rect 20074 29416 20130 29472
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 20166 29008 20222 29064
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 20534 29144 20590 29200
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19890 15000 19946 15056
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 18786 3304 18842 3360
rect 18786 2624 18842 2680
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19430 8336 19486 8392
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 20626 28952 20682 29008
rect 20626 24520 20682 24576
rect 20810 15444 20812 15464
rect 20812 15444 20864 15464
rect 20864 15444 20866 15464
rect 20810 15408 20866 15444
rect 20534 13524 20590 13560
rect 20534 13504 20536 13524
rect 20536 13504 20588 13524
rect 20588 13504 20590 13524
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19890 3032 19946 3088
rect 19798 2796 19800 2816
rect 19800 2796 19852 2816
rect 19852 2796 19854 2816
rect 19798 2760 19854 2796
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20258 3732 20314 3768
rect 20258 3712 20260 3732
rect 20260 3712 20312 3732
rect 20312 3712 20314 3732
rect 20442 3032 20498 3088
rect 21914 29280 21970 29336
rect 21914 29008 21970 29064
rect 22190 29416 22246 29472
rect 22190 24520 22246 24576
rect 21914 17176 21970 17232
rect 22190 14884 22246 14920
rect 22190 14864 22192 14884
rect 22192 14864 22244 14884
rect 22244 14864 22246 14884
rect 24766 32408 24822 32464
rect 24490 29280 24546 29336
rect 24674 29824 24730 29880
rect 24214 23704 24270 23760
rect 24490 23740 24492 23760
rect 24492 23740 24544 23760
rect 24544 23740 24546 23760
rect 24490 23704 24546 23740
rect 21362 7404 21418 7440
rect 21362 7384 21364 7404
rect 21364 7384 21416 7404
rect 21416 7384 21418 7404
rect 20994 3168 21050 3224
rect 21270 2624 21326 2680
rect 22926 5480 22982 5536
rect 22374 3168 22430 3224
rect 23018 3188 23074 3224
rect 23018 3168 23020 3188
rect 23020 3168 23072 3188
rect 23072 3168 23074 3188
rect 23662 7520 23718 7576
rect 25042 16532 25044 16552
rect 25044 16532 25096 16552
rect 25096 16532 25098 16552
rect 25042 16496 25098 16532
rect 24674 6840 24730 6896
rect 26790 55256 26846 55312
rect 29918 56228 29974 56264
rect 29918 56208 29920 56228
rect 29920 56208 29972 56228
rect 29972 56208 29974 56228
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 32126 53080 32182 53136
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 30930 50224 30986 50280
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 29182 47504 29238 47560
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 27986 44784 28042 44840
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 26146 29164 26202 29200
rect 26146 29144 26148 29164
rect 26148 29144 26200 29164
rect 26200 29144 26202 29164
rect 25410 23704 25466 23760
rect 25778 7520 25834 7576
rect 26606 17212 26608 17232
rect 26608 17212 26660 17232
rect 26660 17212 26662 17232
rect 26606 17176 26662 17212
rect 26974 19760 27030 19816
rect 28262 32000 28318 32056
rect 28538 32000 28594 32056
rect 27250 15000 27306 15056
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 29274 26288 29330 26344
rect 28262 15000 28318 15056
rect 28170 13504 28226 13560
rect 28170 7404 28226 7440
rect 28170 7384 28172 7404
rect 28172 7384 28224 7404
rect 28224 7384 28226 7404
rect 26330 2896 26386 2952
rect 29550 5616 29606 5672
rect 29366 2352 29422 2408
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 30654 20440 30710 20496
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 29918 5616 29974 5672
rect 30654 5652 30656 5672
rect 30656 5652 30708 5672
rect 30708 5652 30710 5672
rect 30654 5616 30710 5652
rect 29642 5108 29644 5128
rect 29644 5108 29696 5128
rect 29696 5108 29698 5128
rect 29642 5072 29698 5108
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 35346 14900 35348 14920
rect 35348 14900 35400 14920
rect 35400 14900 35402 14920
rect 35346 14864 35402 14900
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 57518 57840 57574 57896
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 57886 56480 57942 56536
rect 43810 37848 43866 37904
rect 36818 16496 36874 16552
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 58162 55140 58218 55176
rect 58162 55120 58164 55140
rect 58164 55120 58216 55140
rect 58216 55120 58218 55140
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 57886 53760 57942 53816
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 57886 52436 57888 52456
rect 57888 52436 57940 52456
rect 57940 52436 57942 52456
rect 57886 52400 57942 52436
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 58162 51040 58218 51096
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 58162 49716 58164 49736
rect 58164 49716 58216 49736
rect 58216 49716 58218 49736
rect 58162 49680 58218 49716
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 58162 48320 58218 48376
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 58162 46996 58164 47016
rect 58164 46996 58216 47016
rect 58216 46996 58218 47016
rect 58162 46960 58218 46996
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 58162 45600 58218 45656
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 58162 44260 58218 44296
rect 58162 44240 58164 44260
rect 58164 44240 58216 44260
rect 58216 44240 58218 44260
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 58162 42880 58218 42936
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 58162 41556 58164 41576
rect 58164 41556 58216 41576
rect 58216 41556 58218 41576
rect 58162 41520 58218 41556
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 58162 40160 58218 40216
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 58162 38820 58218 38856
rect 58162 38800 58164 38820
rect 58164 38800 58216 38820
rect 58216 38800 58218 38820
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 58162 37440 58218 37496
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 58162 36116 58164 36136
rect 58164 36116 58216 36136
rect 58216 36116 58218 36136
rect 58162 36080 58218 36116
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 58162 34720 58218 34776
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 58162 33380 58218 33416
rect 58162 33360 58164 33380
rect 58164 33360 58216 33380
rect 58216 33360 58218 33380
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 58162 32000 58218 32056
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 58162 30676 58164 30696
rect 58164 30676 58216 30696
rect 58216 30676 58218 30696
rect 58162 30640 58218 30676
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 58162 29280 58218 29336
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 58162 27940 58218 27976
rect 58162 27920 58164 27940
rect 58164 27920 58216 27940
rect 58216 27920 58218 27940
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 58162 26560 58218 26616
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 58162 25236 58164 25256
rect 58164 25236 58216 25256
rect 58216 25236 58218 25256
rect 58162 25200 58218 25236
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 58162 23840 58218 23896
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 58162 22500 58218 22536
rect 58162 22480 58164 22500
rect 58164 22480 58216 22500
rect 58216 22480 58218 22500
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 58162 21120 58218 21176
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 58162 19796 58164 19816
rect 58164 19796 58216 19816
rect 58216 19796 58218 19816
rect 58162 19760 58218 19796
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 58162 18400 58218 18456
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 58162 17060 58218 17096
rect 58162 17040 58164 17060
rect 58164 17040 58216 17060
rect 58216 17040 58218 17060
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 58162 15680 58218 15736
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 58162 14356 58164 14376
rect 58164 14356 58216 14376
rect 58216 14356 58218 14376
rect 58162 14320 58218 14356
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 58162 12960 58218 13016
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 58162 11620 58218 11656
rect 58162 11600 58164 11620
rect 58164 11600 58216 11620
rect 58216 11600 58218 11620
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 58162 10240 58218 10296
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 58162 8916 58164 8936
rect 58164 8916 58216 8936
rect 58216 8916 58218 8936
rect 58162 8880 58218 8916
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 58162 7520 58218 7576
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 58162 6180 58218 6216
rect 58162 6160 58164 6180
rect 58164 6160 58216 6180
rect 58216 6160 58218 6180
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 53378 2896 53434 2952
rect 53470 2760 53526 2816
rect 58162 4800 58218 4856
rect 58162 3476 58164 3496
rect 58164 3476 58216 3496
rect 58216 3476 58218 3496
rect 56598 2932 56600 2952
rect 56600 2932 56652 2952
rect 56652 2932 56654 2952
rect 56598 2896 56654 2932
rect 55310 2760 55366 2816
rect 58162 3440 58218 3476
rect 57518 2080 57574 2136
rect 58438 720 58494 776
<< metal3 >>
rect 58433 59258 58499 59261
rect 59200 59258 60000 59288
rect 58433 59256 60000 59258
rect 58433 59200 58438 59256
rect 58494 59200 60000 59256
rect 58433 59198 60000 59200
rect 58433 59195 58499 59198
rect 59200 59168 60000 59198
rect 57513 57898 57579 57901
rect 59200 57898 60000 57928
rect 57513 57896 60000 57898
rect 57513 57840 57518 57896
rect 57574 57840 60000 57896
rect 57513 57838 60000 57840
rect 57513 57835 57579 57838
rect 59200 57808 60000 57838
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 18638 56748 18644 56812
rect 18708 56810 18714 56812
rect 20161 56810 20227 56813
rect 18708 56808 20227 56810
rect 18708 56752 20166 56808
rect 20222 56752 20227 56808
rect 18708 56750 20227 56752
rect 18708 56748 18714 56750
rect 20161 56747 20227 56750
rect 0 56674 800 56704
rect 1393 56674 1459 56677
rect 0 56672 1459 56674
rect 0 56616 1398 56672
rect 1454 56616 1459 56672
rect 0 56614 1459 56616
rect 0 56584 800 56614
rect 1393 56611 1459 56614
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 57881 56538 57947 56541
rect 59200 56538 60000 56568
rect 57881 56536 60000 56538
rect 57881 56480 57886 56536
rect 57942 56480 60000 56536
rect 57881 56478 60000 56480
rect 57881 56475 57947 56478
rect 59200 56448 60000 56478
rect 23974 56204 23980 56268
rect 24044 56266 24050 56268
rect 29913 56266 29979 56269
rect 24044 56264 29979 56266
rect 24044 56208 29918 56264
rect 29974 56208 29979 56264
rect 24044 56206 29979 56208
rect 24044 56204 24050 56206
rect 29913 56203 29979 56206
rect 14181 56132 14247 56133
rect 14181 56130 14228 56132
rect 14136 56128 14228 56130
rect 14136 56072 14186 56128
rect 14136 56070 14228 56072
rect 14181 56068 14228 56070
rect 14292 56068 14298 56132
rect 14181 56067 14247 56068
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 0 55586 800 55616
rect 1393 55586 1459 55589
rect 0 55584 1459 55586
rect 0 55528 1398 55584
rect 1454 55528 1459 55584
rect 0 55526 1459 55528
rect 0 55496 800 55526
rect 1393 55523 1459 55526
rect 17033 55586 17099 55589
rect 17677 55588 17743 55589
rect 20253 55588 20319 55589
rect 17677 55586 17724 55588
rect 17033 55584 17724 55586
rect 17033 55528 17038 55584
rect 17094 55528 17682 55584
rect 17033 55526 17724 55528
rect 17033 55523 17099 55526
rect 17677 55524 17724 55526
rect 17788 55524 17794 55588
rect 20253 55586 20300 55588
rect 20208 55584 20300 55586
rect 20208 55528 20258 55584
rect 20208 55526 20300 55528
rect 20253 55524 20300 55526
rect 20364 55524 20370 55588
rect 21214 55524 21220 55588
rect 21284 55586 21290 55588
rect 21725 55586 21791 55589
rect 21284 55584 21791 55586
rect 21284 55528 21730 55584
rect 21786 55528 21791 55584
rect 21284 55526 21791 55528
rect 21284 55524 21290 55526
rect 17677 55523 17743 55524
rect 20253 55523 20319 55524
rect 21725 55523 21791 55526
rect 22318 55524 22324 55588
rect 22388 55586 22394 55588
rect 23013 55586 23079 55589
rect 23749 55588 23815 55589
rect 23749 55586 23796 55588
rect 22388 55584 23079 55586
rect 22388 55528 23018 55584
rect 23074 55528 23079 55584
rect 22388 55526 23079 55528
rect 23704 55584 23796 55586
rect 23704 55528 23754 55584
rect 23704 55526 23796 55528
rect 22388 55524 22394 55526
rect 23013 55523 23079 55526
rect 23749 55524 23796 55526
rect 23860 55524 23866 55588
rect 23749 55523 23815 55524
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 17534 55252 17540 55316
rect 17604 55314 17610 55316
rect 17769 55314 17835 55317
rect 18781 55316 18847 55317
rect 18781 55314 18828 55316
rect 17604 55312 17835 55314
rect 17604 55256 17774 55312
rect 17830 55256 17835 55312
rect 17604 55254 17835 55256
rect 18736 55312 18828 55314
rect 18736 55256 18786 55312
rect 18736 55254 18828 55256
rect 17604 55252 17610 55254
rect 17769 55251 17835 55254
rect 18781 55252 18828 55254
rect 18892 55252 18898 55316
rect 19793 55314 19859 55317
rect 20110 55314 20116 55316
rect 19793 55312 20116 55314
rect 19793 55256 19798 55312
rect 19854 55256 20116 55312
rect 19793 55254 20116 55256
rect 18781 55251 18847 55252
rect 19793 55251 19859 55254
rect 20110 55252 20116 55254
rect 20180 55252 20186 55316
rect 21398 55252 21404 55316
rect 21468 55314 21474 55316
rect 26785 55314 26851 55317
rect 21468 55312 26851 55314
rect 21468 55256 26790 55312
rect 26846 55256 26851 55312
rect 21468 55254 26851 55256
rect 21468 55252 21474 55254
rect 26785 55251 26851 55254
rect 58157 55178 58223 55181
rect 59200 55178 60000 55208
rect 58157 55176 60000 55178
rect 58157 55120 58162 55176
rect 58218 55120 60000 55176
rect 58157 55118 60000 55120
rect 58157 55115 58223 55118
rect 59200 55088 60000 55118
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 0 54498 800 54528
rect 1393 54498 1459 54501
rect 0 54496 1459 54498
rect 0 54440 1398 54496
rect 1454 54440 1459 54496
rect 0 54438 1459 54440
rect 0 54408 800 54438
rect 1393 54435 1459 54438
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 57881 53818 57947 53821
rect 59200 53818 60000 53848
rect 57881 53816 60000 53818
rect 57881 53760 57886 53816
rect 57942 53760 60000 53816
rect 57881 53758 60000 53760
rect 57881 53755 57947 53758
rect 59200 53728 60000 53758
rect 0 53410 800 53440
rect 1393 53410 1459 53413
rect 0 53408 1459 53410
rect 0 53352 1398 53408
rect 1454 53352 1459 53408
rect 0 53350 1459 53352
rect 0 53320 800 53350
rect 1393 53347 1459 53350
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 14590 53076 14596 53140
rect 14660 53138 14666 53140
rect 32121 53138 32187 53141
rect 14660 53136 32187 53138
rect 14660 53080 32126 53136
rect 32182 53080 32187 53136
rect 14660 53078 32187 53080
rect 14660 53076 14666 53078
rect 32121 53075 32187 53078
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 57881 52458 57947 52461
rect 59200 52458 60000 52488
rect 57881 52456 60000 52458
rect 57881 52400 57886 52456
rect 57942 52400 60000 52456
rect 57881 52398 60000 52400
rect 57881 52395 57947 52398
rect 59200 52368 60000 52398
rect 0 52322 800 52352
rect 1393 52322 1459 52325
rect 0 52320 1459 52322
rect 0 52264 1398 52320
rect 1454 52264 1459 52320
rect 0 52262 1459 52264
rect 0 52232 800 52262
rect 1393 52259 1459 52262
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 0 51234 800 51264
rect 1393 51234 1459 51237
rect 0 51232 1459 51234
rect 0 51176 1398 51232
rect 1454 51176 1459 51232
rect 0 51174 1459 51176
rect 0 51144 800 51174
rect 1393 51171 1459 51174
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 58157 51098 58223 51101
rect 59200 51098 60000 51128
rect 58157 51096 60000 51098
rect 58157 51040 58162 51096
rect 58218 51040 60000 51096
rect 58157 51038 60000 51040
rect 58157 51035 58223 51038
rect 59200 51008 60000 51038
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 14774 50220 14780 50284
rect 14844 50282 14850 50284
rect 30925 50282 30991 50285
rect 14844 50280 30991 50282
rect 14844 50224 30930 50280
rect 30986 50224 30991 50280
rect 14844 50222 30991 50224
rect 14844 50220 14850 50222
rect 30925 50219 30991 50222
rect 0 50146 800 50176
rect 1393 50146 1459 50149
rect 0 50144 1459 50146
rect 0 50088 1398 50144
rect 1454 50088 1459 50144
rect 0 50086 1459 50088
rect 0 50056 800 50086
rect 1393 50083 1459 50086
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 58157 49738 58223 49741
rect 59200 49738 60000 49768
rect 58157 49736 60000 49738
rect 58157 49680 58162 49736
rect 58218 49680 60000 49736
rect 58157 49678 60000 49680
rect 58157 49675 58223 49678
rect 59200 49648 60000 49678
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 0 49058 800 49088
rect 1393 49058 1459 49061
rect 0 49056 1459 49058
rect 0 49000 1398 49056
rect 1454 49000 1459 49056
rect 0 48998 1459 49000
rect 0 48968 800 48998
rect 1393 48995 1459 48998
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 58157 48378 58223 48381
rect 59200 48378 60000 48408
rect 58157 48376 60000 48378
rect 58157 48320 58162 48376
rect 58218 48320 60000 48376
rect 58157 48318 60000 48320
rect 58157 48315 58223 48318
rect 59200 48288 60000 48318
rect 0 47970 800 48000
rect 1393 47970 1459 47973
rect 0 47968 1459 47970
rect 0 47912 1398 47968
rect 1454 47912 1459 47968
rect 0 47910 1459 47912
rect 0 47880 800 47910
rect 1393 47907 1459 47910
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 15878 47500 15884 47564
rect 15948 47562 15954 47564
rect 29177 47562 29243 47565
rect 15948 47560 29243 47562
rect 15948 47504 29182 47560
rect 29238 47504 29243 47560
rect 15948 47502 29243 47504
rect 15948 47500 15954 47502
rect 29177 47499 29243 47502
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 58157 47018 58223 47021
rect 59200 47018 60000 47048
rect 58157 47016 60000 47018
rect 58157 46960 58162 47016
rect 58218 46960 60000 47016
rect 58157 46958 60000 46960
rect 58157 46955 58223 46958
rect 59200 46928 60000 46958
rect 0 46792 800 46912
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 0 45704 800 45824
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 58157 45658 58223 45661
rect 59200 45658 60000 45688
rect 58157 45656 60000 45658
rect 58157 45600 58162 45656
rect 58218 45600 60000 45656
rect 58157 45598 60000 45600
rect 58157 45595 58223 45598
rect 59200 45568 60000 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 15326 44780 15332 44844
rect 15396 44842 15402 44844
rect 27981 44842 28047 44845
rect 15396 44840 28047 44842
rect 15396 44784 27986 44840
rect 28042 44784 28047 44840
rect 15396 44782 28047 44784
rect 15396 44780 15402 44782
rect 27981 44779 28047 44782
rect 0 44616 800 44736
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 58157 44298 58223 44301
rect 59200 44298 60000 44328
rect 58157 44296 60000 44298
rect 58157 44240 58162 44296
rect 58218 44240 60000 44296
rect 58157 44238 60000 44240
rect 58157 44235 58223 44238
rect 59200 44208 60000 44238
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 0 43528 800 43648
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 58157 42938 58223 42941
rect 59200 42938 60000 42968
rect 58157 42936 60000 42938
rect 58157 42880 58162 42936
rect 58218 42880 60000 42936
rect 58157 42878 60000 42880
rect 58157 42875 58223 42878
rect 59200 42848 60000 42878
rect 0 42440 800 42560
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 17350 41652 17356 41716
rect 17420 41714 17426 41716
rect 19977 41714 20043 41717
rect 17420 41712 20043 41714
rect 17420 41656 19982 41712
rect 20038 41656 20043 41712
rect 17420 41654 20043 41656
rect 17420 41652 17426 41654
rect 19977 41651 20043 41654
rect 58157 41578 58223 41581
rect 59200 41578 60000 41608
rect 58157 41576 60000 41578
rect 58157 41520 58162 41576
rect 58218 41520 60000 41576
rect 58157 41518 60000 41520
rect 58157 41515 58223 41518
rect 59200 41488 60000 41518
rect 0 41352 800 41472
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 0 40264 800 40384
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 58157 40218 58223 40221
rect 59200 40218 60000 40248
rect 58157 40216 60000 40218
rect 58157 40160 58162 40216
rect 58218 40160 60000 40216
rect 58157 40158 60000 40160
rect 58157 40155 58223 40158
rect 59200 40128 60000 40158
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 0 39176 800 39296
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 58157 38858 58223 38861
rect 59200 38858 60000 38888
rect 58157 38856 60000 38858
rect 58157 38800 58162 38856
rect 58218 38800 60000 38856
rect 58157 38798 60000 38800
rect 58157 38795 58223 38798
rect 59200 38768 60000 38798
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 4889 38314 4955 38317
rect 6729 38314 6795 38317
rect 4889 38312 6795 38314
rect 4889 38256 4894 38312
rect 4950 38256 6734 38312
rect 6790 38256 6795 38312
rect 4889 38254 6795 38256
rect 4889 38251 4955 38254
rect 6729 38251 6795 38254
rect 0 38088 800 38208
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 10409 38042 10475 38045
rect 16757 38042 16823 38045
rect 10409 38040 16823 38042
rect 10409 37984 10414 38040
rect 10470 37984 16762 38040
rect 16818 37984 16823 38040
rect 10409 37982 16823 37984
rect 10409 37979 10475 37982
rect 16757 37979 16823 37982
rect 23054 37844 23060 37908
rect 23124 37906 23130 37908
rect 43805 37906 43871 37909
rect 23124 37904 43871 37906
rect 23124 37848 43810 37904
rect 43866 37848 43871 37904
rect 23124 37846 43871 37848
rect 23124 37844 23130 37846
rect 43805 37843 43871 37846
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 58157 37498 58223 37501
rect 59200 37498 60000 37528
rect 58157 37496 60000 37498
rect 58157 37440 58162 37496
rect 58218 37440 60000 37496
rect 58157 37438 60000 37440
rect 58157 37435 58223 37438
rect 59200 37408 60000 37438
rect 0 37000 800 37120
rect 13537 37090 13603 37093
rect 17861 37090 17927 37093
rect 13537 37088 17927 37090
rect 13537 37032 13542 37088
rect 13598 37032 17866 37088
rect 17922 37032 17927 37088
rect 13537 37030 17927 37032
rect 13537 37027 13603 37030
rect 17861 37027 17927 37030
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 58157 36138 58223 36141
rect 59200 36138 60000 36168
rect 58157 36136 60000 36138
rect 58157 36080 58162 36136
rect 58218 36080 60000 36136
rect 58157 36078 60000 36080
rect 58157 36075 58223 36078
rect 59200 36048 60000 36078
rect 0 35912 800 36032
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 0 34824 800 34944
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 58157 34778 58223 34781
rect 59200 34778 60000 34808
rect 58157 34776 60000 34778
rect 58157 34720 58162 34776
rect 58218 34720 60000 34776
rect 58157 34718 60000 34720
rect 58157 34715 58223 34718
rect 59200 34688 60000 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 9581 34234 9647 34237
rect 14549 34234 14615 34237
rect 9581 34232 14615 34234
rect 9581 34176 9586 34232
rect 9642 34176 14554 34232
rect 14610 34176 14615 34232
rect 9581 34174 14615 34176
rect 9581 34171 9647 34174
rect 14549 34171 14615 34174
rect 0 33736 800 33856
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 58157 33418 58223 33421
rect 59200 33418 60000 33448
rect 58157 33416 60000 33418
rect 58157 33360 58162 33416
rect 58218 33360 60000 33416
rect 58157 33358 60000 33360
rect 58157 33355 58223 33358
rect 59200 33328 60000 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 0 32648 800 32768
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 17953 32466 18019 32469
rect 24761 32466 24827 32469
rect 17953 32464 24827 32466
rect 17953 32408 17958 32464
rect 18014 32408 24766 32464
rect 24822 32408 24827 32464
rect 17953 32406 24827 32408
rect 17953 32403 18019 32406
rect 24761 32403 24827 32406
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 28257 32058 28323 32061
rect 28533 32058 28599 32061
rect 28257 32056 28599 32058
rect 28257 32000 28262 32056
rect 28318 32000 28538 32056
rect 28594 32000 28599 32056
rect 28257 31998 28599 32000
rect 28257 31995 28323 31998
rect 28533 31995 28599 31998
rect 58157 32058 58223 32061
rect 59200 32058 60000 32088
rect 58157 32056 60000 32058
rect 58157 32000 58162 32056
rect 58218 32000 60000 32056
rect 58157 31998 60000 32000
rect 58157 31995 58223 31998
rect 59200 31968 60000 31998
rect 0 31560 800 31680
rect 5625 31650 5691 31653
rect 11329 31650 11395 31653
rect 5625 31648 11395 31650
rect 5625 31592 5630 31648
rect 5686 31592 11334 31648
rect 11390 31592 11395 31648
rect 5625 31590 11395 31592
rect 5625 31587 5691 31590
rect 11329 31587 11395 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 8293 31514 8359 31517
rect 16849 31514 16915 31517
rect 8293 31512 16915 31514
rect 8293 31456 8298 31512
rect 8354 31456 16854 31512
rect 16910 31456 16915 31512
rect 8293 31454 16915 31456
rect 8293 31451 8359 31454
rect 16849 31451 16915 31454
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 58157 30698 58223 30701
rect 59200 30698 60000 30728
rect 58157 30696 60000 30698
rect 58157 30640 58162 30696
rect 58218 30640 60000 30696
rect 58157 30638 60000 30640
rect 58157 30635 58223 30638
rect 59200 30608 60000 30638
rect 0 30472 800 30592
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 20161 29882 20227 29885
rect 24669 29882 24735 29885
rect 20161 29880 24735 29882
rect 20161 29824 20166 29880
rect 20222 29824 24674 29880
rect 24730 29824 24735 29880
rect 20161 29822 24735 29824
rect 20161 29819 20227 29822
rect 24669 29819 24735 29822
rect 0 29384 800 29504
rect 20069 29474 20135 29477
rect 22185 29474 22251 29477
rect 20069 29472 22251 29474
rect 20069 29416 20074 29472
rect 20130 29416 22190 29472
rect 22246 29416 22251 29472
rect 20069 29414 22251 29416
rect 20069 29411 20135 29414
rect 22185 29411 22251 29414
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 21909 29338 21975 29341
rect 24485 29338 24551 29341
rect 20302 29278 21834 29338
rect 19885 29202 19951 29205
rect 20302 29202 20362 29278
rect 20529 29202 20595 29205
rect 19885 29200 20362 29202
rect 19885 29144 19890 29200
rect 19946 29144 20362 29200
rect 19885 29142 20362 29144
rect 20486 29200 20595 29202
rect 20486 29144 20534 29200
rect 20590 29144 20595 29200
rect 19885 29139 19951 29142
rect 20486 29139 20595 29144
rect 21774 29202 21834 29278
rect 21909 29336 24551 29338
rect 21909 29280 21914 29336
rect 21970 29280 24490 29336
rect 24546 29280 24551 29336
rect 21909 29278 24551 29280
rect 21909 29275 21975 29278
rect 24485 29275 24551 29278
rect 58157 29338 58223 29341
rect 59200 29338 60000 29368
rect 58157 29336 60000 29338
rect 58157 29280 58162 29336
rect 58218 29280 60000 29336
rect 58157 29278 60000 29280
rect 58157 29275 58223 29278
rect 59200 29248 60000 29278
rect 26141 29202 26207 29205
rect 21774 29200 26207 29202
rect 21774 29144 26146 29200
rect 26202 29144 26207 29200
rect 21774 29142 26207 29144
rect 26141 29139 26207 29142
rect 20161 29066 20227 29069
rect 20486 29066 20546 29139
rect 21909 29066 21975 29069
rect 20161 29064 20546 29066
rect 20161 29008 20166 29064
rect 20222 29008 20546 29064
rect 20670 29064 21975 29066
rect 20670 29013 21914 29064
rect 20161 29006 20546 29008
rect 20621 29008 21914 29013
rect 21970 29008 21975 29064
rect 20161 29003 20227 29006
rect 20621 28952 20626 29008
rect 20682 29006 21975 29008
rect 20682 28952 20730 29006
rect 21909 29003 21975 29006
rect 20621 28950 20730 28952
rect 20621 28947 20687 28950
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 0 28296 800 28416
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 58157 27978 58223 27981
rect 59200 27978 60000 28008
rect 58157 27976 60000 27978
rect 58157 27920 58162 27976
rect 58218 27920 60000 27976
rect 58157 27918 60000 27920
rect 58157 27915 58223 27918
rect 59200 27888 60000 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 0 27208 800 27328
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 58157 26618 58223 26621
rect 59200 26618 60000 26648
rect 58157 26616 60000 26618
rect 58157 26560 58162 26616
rect 58218 26560 60000 26616
rect 58157 26558 60000 26560
rect 58157 26555 58223 26558
rect 59200 26528 60000 26558
rect 17217 26482 17283 26485
rect 18873 26482 18939 26485
rect 17217 26480 18939 26482
rect 17217 26424 17222 26480
rect 17278 26424 18878 26480
rect 18934 26424 18939 26480
rect 17217 26422 18939 26424
rect 17217 26419 17283 26422
rect 18873 26419 18939 26422
rect 16757 26346 16823 26349
rect 17033 26346 17099 26349
rect 29269 26346 29335 26349
rect 16757 26344 29335 26346
rect 16757 26288 16762 26344
rect 16818 26288 17038 26344
rect 17094 26288 29274 26344
rect 29330 26288 29335 26344
rect 16757 26286 29335 26288
rect 16757 26283 16823 26286
rect 17033 26283 17099 26286
rect 29269 26283 29335 26286
rect 0 26120 800 26240
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 58157 25258 58223 25261
rect 59200 25258 60000 25288
rect 58157 25256 60000 25258
rect 58157 25200 58162 25256
rect 58218 25200 60000 25256
rect 58157 25198 60000 25200
rect 58157 25195 58223 25198
rect 59200 25168 60000 25198
rect 0 25032 800 25152
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 20621 24578 20687 24581
rect 22185 24578 22251 24581
rect 20621 24576 22251 24578
rect 20621 24520 20626 24576
rect 20682 24520 22190 24576
rect 22246 24520 22251 24576
rect 20621 24518 22251 24520
rect 20621 24515 20687 24518
rect 22185 24515 22251 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 9857 24170 9923 24173
rect 16665 24170 16731 24173
rect 9857 24168 16731 24170
rect 9857 24112 9862 24168
rect 9918 24112 16670 24168
rect 16726 24112 16731 24168
rect 9857 24110 16731 24112
rect 9857 24107 9923 24110
rect 16665 24107 16731 24110
rect 0 23944 800 24064
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 58157 23898 58223 23901
rect 59200 23898 60000 23928
rect 58157 23896 60000 23898
rect 58157 23840 58162 23896
rect 58218 23840 60000 23896
rect 58157 23838 60000 23840
rect 58157 23835 58223 23838
rect 59200 23808 60000 23838
rect 18505 23762 18571 23765
rect 24209 23762 24275 23765
rect 24485 23762 24551 23765
rect 25405 23762 25471 23765
rect 18505 23760 25471 23762
rect 18505 23704 18510 23760
rect 18566 23704 24214 23760
rect 24270 23704 24490 23760
rect 24546 23704 25410 23760
rect 25466 23704 25471 23760
rect 18505 23702 25471 23704
rect 18505 23699 18571 23702
rect 24209 23699 24275 23702
rect 24485 23699 24551 23702
rect 25405 23699 25471 23702
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 0 22856 800 22976
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 58157 22538 58223 22541
rect 59200 22538 60000 22568
rect 58157 22536 60000 22538
rect 58157 22480 58162 22536
rect 58218 22480 60000 22536
rect 58157 22478 60000 22480
rect 58157 22475 58223 22478
rect 59200 22448 60000 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 0 21768 800 21888
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 58157 21178 58223 21181
rect 59200 21178 60000 21208
rect 58157 21176 60000 21178
rect 58157 21120 58162 21176
rect 58218 21120 60000 21176
rect 58157 21118 60000 21120
rect 58157 21115 58223 21118
rect 59200 21088 60000 21118
rect 0 20680 800 20800
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 17677 20498 17743 20501
rect 30649 20498 30715 20501
rect 17677 20496 30715 20498
rect 17677 20440 17682 20496
rect 17738 20440 30654 20496
rect 30710 20440 30715 20496
rect 17677 20438 30715 20440
rect 17677 20435 17743 20438
rect 30649 20435 30715 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 6678 19892 6684 19956
rect 6748 19954 6754 19956
rect 19241 19954 19307 19957
rect 6748 19952 19307 19954
rect 6748 19896 19246 19952
rect 19302 19896 19307 19952
rect 6748 19894 19307 19896
rect 6748 19892 6754 19894
rect 19241 19891 19307 19894
rect 14825 19818 14891 19821
rect 26969 19818 27035 19821
rect 14825 19816 27035 19818
rect 14825 19760 14830 19816
rect 14886 19760 26974 19816
rect 27030 19760 27035 19816
rect 14825 19758 27035 19760
rect 14825 19755 14891 19758
rect 26969 19755 27035 19758
rect 58157 19818 58223 19821
rect 59200 19818 60000 19848
rect 58157 19816 60000 19818
rect 58157 19760 58162 19816
rect 58218 19760 60000 19816
rect 58157 19758 60000 19760
rect 58157 19755 58223 19758
rect 59200 19728 60000 19758
rect 0 19592 800 19712
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 4613 19276 4679 19277
rect 4613 19274 4660 19276
rect 4568 19272 4660 19274
rect 4568 19216 4618 19272
rect 4568 19214 4660 19216
rect 4613 19212 4660 19214
rect 4724 19212 4730 19276
rect 4613 19211 4679 19212
rect 10685 19138 10751 19141
rect 11697 19138 11763 19141
rect 10685 19136 11763 19138
rect 10685 19080 10690 19136
rect 10746 19080 11702 19136
rect 11758 19080 11763 19136
rect 10685 19078 11763 19080
rect 10685 19075 10751 19078
rect 11697 19075 11763 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 0 18504 800 18624
rect 4153 18594 4219 18597
rect 4654 18594 4660 18596
rect 4153 18592 4660 18594
rect 4153 18536 4158 18592
rect 4214 18536 4660 18592
rect 4153 18534 4660 18536
rect 4153 18531 4219 18534
rect 4654 18532 4660 18534
rect 4724 18532 4730 18596
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 58157 18458 58223 18461
rect 59200 18458 60000 18488
rect 58157 18456 60000 18458
rect 58157 18400 58162 18456
rect 58218 18400 60000 18456
rect 58157 18398 60000 18400
rect 58157 18395 58223 18398
rect 59200 18368 60000 18398
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 0 17416 800 17536
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 21909 17234 21975 17237
rect 26601 17234 26667 17237
rect 21909 17232 26667 17234
rect 21909 17176 21914 17232
rect 21970 17176 26606 17232
rect 26662 17176 26667 17232
rect 21909 17174 26667 17176
rect 21909 17171 21975 17174
rect 26601 17171 26667 17174
rect 58157 17098 58223 17101
rect 59200 17098 60000 17128
rect 58157 17096 60000 17098
rect 58157 17040 58162 17096
rect 58218 17040 60000 17096
rect 58157 17038 60000 17040
rect 58157 17035 58223 17038
rect 59200 17008 60000 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 25037 16554 25103 16557
rect 36813 16554 36879 16557
rect 25037 16552 36879 16554
rect 25037 16496 25042 16552
rect 25098 16496 36818 16552
rect 36874 16496 36879 16552
rect 25037 16494 36879 16496
rect 25037 16491 25103 16494
rect 36813 16491 36879 16494
rect 0 16328 800 16448
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 58157 15738 58223 15741
rect 59200 15738 60000 15768
rect 58157 15736 60000 15738
rect 58157 15680 58162 15736
rect 58218 15680 60000 15736
rect 58157 15678 60000 15680
rect 58157 15675 58223 15678
rect 59200 15648 60000 15678
rect 10961 15466 11027 15469
rect 20805 15466 20871 15469
rect 10961 15464 20871 15466
rect 10961 15408 10966 15464
rect 11022 15408 20810 15464
rect 20866 15408 20871 15464
rect 10961 15406 20871 15408
rect 10961 15403 11027 15406
rect 20805 15403 20871 15406
rect 0 15240 800 15360
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 5574 15132 5580 15196
rect 5644 15194 5650 15196
rect 7373 15194 7439 15197
rect 5644 15192 7439 15194
rect 5644 15136 7378 15192
rect 7434 15136 7439 15192
rect 5644 15134 7439 15136
rect 5644 15132 5650 15134
rect 7373 15131 7439 15134
rect 19885 15058 19951 15061
rect 27245 15058 27311 15061
rect 28257 15058 28323 15061
rect 19885 15056 28323 15058
rect 19885 15000 19890 15056
rect 19946 15000 27250 15056
rect 27306 15000 28262 15056
rect 28318 15000 28323 15056
rect 19885 14998 28323 15000
rect 19885 14995 19951 14998
rect 27245 14995 27311 14998
rect 28257 14995 28323 14998
rect 22185 14922 22251 14925
rect 35341 14922 35407 14925
rect 22185 14920 35407 14922
rect 22185 14864 22190 14920
rect 22246 14864 35346 14920
rect 35402 14864 35407 14920
rect 22185 14862 35407 14864
rect 22185 14859 22251 14862
rect 35341 14859 35407 14862
rect 8702 14724 8708 14788
rect 8772 14786 8778 14788
rect 8845 14786 8911 14789
rect 8772 14784 8911 14786
rect 8772 14728 8850 14784
rect 8906 14728 8911 14784
rect 8772 14726 8911 14728
rect 8772 14724 8778 14726
rect 8845 14723 8911 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 58157 14378 58223 14381
rect 59200 14378 60000 14408
rect 58157 14376 60000 14378
rect 58157 14320 58162 14376
rect 58218 14320 60000 14376
rect 58157 14318 60000 14320
rect 58157 14315 58223 14318
rect 59200 14288 60000 14318
rect 0 14152 800 14272
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 5533 13834 5599 13837
rect 6494 13834 6500 13836
rect 5533 13832 6500 13834
rect 5533 13776 5538 13832
rect 5594 13776 6500 13832
rect 5533 13774 6500 13776
rect 5533 13771 5599 13774
rect 6494 13772 6500 13774
rect 6564 13772 6570 13836
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 20529 13562 20595 13565
rect 28165 13562 28231 13565
rect 20529 13560 28231 13562
rect 20529 13504 20534 13560
rect 20590 13504 28170 13560
rect 28226 13504 28231 13560
rect 20529 13502 28231 13504
rect 20529 13499 20595 13502
rect 28165 13499 28231 13502
rect 0 13064 800 13184
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 58157 13018 58223 13021
rect 59200 13018 60000 13048
rect 58157 13016 60000 13018
rect 58157 12960 58162 13016
rect 58218 12960 60000 13016
rect 58157 12958 60000 12960
rect 58157 12955 58223 12958
rect 59200 12928 60000 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 0 11976 800 12096
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 58157 11658 58223 11661
rect 59200 11658 60000 11688
rect 58157 11656 60000 11658
rect 58157 11600 58162 11656
rect 58218 11600 60000 11656
rect 58157 11598 60000 11600
rect 58157 11595 58223 11598
rect 59200 11568 60000 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 6729 11250 6795 11253
rect 7281 11250 7347 11253
rect 6729 11248 7347 11250
rect 6729 11192 6734 11248
rect 6790 11192 7286 11248
rect 7342 11192 7347 11248
rect 6729 11190 7347 11192
rect 6729 11187 6795 11190
rect 7281 11187 7347 11190
rect 9765 11114 9831 11117
rect 11094 11114 11100 11116
rect 9765 11112 11100 11114
rect 9765 11056 9770 11112
rect 9826 11056 11100 11112
rect 9765 11054 11100 11056
rect 9765 11051 9831 11054
rect 11094 11052 11100 11054
rect 11164 11052 11170 11116
rect 0 10888 800 11008
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 10225 10434 10291 10437
rect 10358 10434 10364 10436
rect 10225 10432 10364 10434
rect 10225 10376 10230 10432
rect 10286 10376 10364 10432
rect 10225 10374 10364 10376
rect 10225 10371 10291 10374
rect 10358 10372 10364 10374
rect 10428 10372 10434 10436
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 58157 10298 58223 10301
rect 59200 10298 60000 10328
rect 58157 10296 60000 10298
rect 58157 10240 58162 10296
rect 58218 10240 60000 10296
rect 58157 10238 60000 10240
rect 58157 10235 58223 10238
rect 59200 10208 60000 10238
rect 16246 9964 16252 10028
rect 16316 10026 16322 10028
rect 21398 10026 21404 10028
rect 16316 9966 21404 10026
rect 16316 9964 16322 9966
rect 21398 9964 21404 9966
rect 21468 9964 21474 10028
rect 0 9800 800 9920
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 20110 9692 20116 9756
rect 20180 9754 20186 9756
rect 20846 9754 20852 9756
rect 20180 9694 20852 9754
rect 20180 9692 20186 9694
rect 20846 9692 20852 9694
rect 20916 9692 20922 9756
rect 3877 9618 3943 9621
rect 8334 9618 8340 9620
rect 3877 9616 8340 9618
rect 3877 9560 3882 9616
rect 3938 9560 8340 9616
rect 3877 9558 8340 9560
rect 3877 9555 3943 9558
rect 8334 9556 8340 9558
rect 8404 9556 8410 9620
rect 11881 9346 11947 9349
rect 15561 9346 15627 9349
rect 11881 9344 15627 9346
rect 11881 9288 11886 9344
rect 11942 9288 15566 9344
rect 15622 9288 15627 9344
rect 11881 9286 15627 9288
rect 11881 9283 11947 9286
rect 15561 9283 15627 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 11789 9074 11855 9077
rect 16573 9074 16639 9077
rect 11789 9072 16639 9074
rect 11789 9016 11794 9072
rect 11850 9016 16578 9072
rect 16634 9016 16639 9072
rect 11789 9014 16639 9016
rect 11789 9011 11855 9014
rect 16573 9011 16639 9014
rect 58157 8938 58223 8941
rect 59200 8938 60000 8968
rect 58157 8936 60000 8938
rect 58157 8880 58162 8936
rect 58218 8880 60000 8936
rect 58157 8878 60000 8880
rect 58157 8875 58223 8878
rect 59200 8848 60000 8878
rect 0 8712 800 8832
rect 2630 8740 2636 8804
rect 2700 8802 2706 8804
rect 6361 8802 6427 8805
rect 2700 8800 6427 8802
rect 2700 8744 6366 8800
rect 6422 8744 6427 8800
rect 2700 8742 6427 8744
rect 2700 8740 2706 8742
rect 6361 8739 6427 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 2037 8666 2103 8669
rect 6085 8666 6151 8669
rect 13353 8666 13419 8669
rect 2037 8664 13419 8666
rect 2037 8608 2042 8664
rect 2098 8608 6090 8664
rect 6146 8608 13358 8664
rect 13414 8608 13419 8664
rect 2037 8606 13419 8608
rect 2037 8603 2103 8606
rect 6085 8603 6151 8606
rect 13353 8603 13419 8606
rect 9438 8468 9444 8532
rect 9508 8530 9514 8532
rect 9581 8530 9647 8533
rect 9508 8528 9647 8530
rect 9508 8472 9586 8528
rect 9642 8472 9647 8528
rect 9508 8470 9647 8472
rect 9508 8468 9514 8470
rect 9581 8467 9647 8470
rect 9765 8530 9831 8533
rect 12249 8530 12315 8533
rect 9765 8528 12315 8530
rect 9765 8472 9770 8528
rect 9826 8472 12254 8528
rect 12310 8472 12315 8528
rect 9765 8470 12315 8472
rect 9765 8467 9831 8470
rect 12249 8467 12315 8470
rect 8150 8332 8156 8396
rect 8220 8394 8226 8396
rect 8569 8394 8635 8397
rect 14733 8394 14799 8397
rect 8220 8392 14799 8394
rect 8220 8336 8574 8392
rect 8630 8336 14738 8392
rect 14794 8336 14799 8392
rect 8220 8334 14799 8336
rect 8220 8332 8226 8334
rect 8569 8331 8635 8334
rect 14733 8331 14799 8334
rect 18822 8332 18828 8396
rect 18892 8394 18898 8396
rect 19425 8394 19491 8397
rect 18892 8392 19491 8394
rect 18892 8336 19430 8392
rect 19486 8336 19491 8392
rect 18892 8334 19491 8336
rect 18892 8332 18898 8334
rect 19425 8331 19491 8334
rect 10910 8196 10916 8260
rect 10980 8258 10986 8260
rect 12433 8258 12499 8261
rect 10980 8256 12499 8258
rect 10980 8200 12438 8256
rect 12494 8200 12499 8256
rect 10980 8198 12499 8200
rect 10980 8196 10986 8198
rect 12433 8195 12499 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 9581 8122 9647 8125
rect 4662 8120 9647 8122
rect 4662 8064 9586 8120
rect 9642 8064 9647 8120
rect 4662 8062 9647 8064
rect 3509 7986 3575 7989
rect 4662 7986 4722 8062
rect 9581 8059 9647 8062
rect 3509 7984 4722 7986
rect 3509 7928 3514 7984
rect 3570 7928 4722 7984
rect 3509 7926 4722 7928
rect 3509 7923 3575 7926
rect 0 7624 800 7744
rect 3969 7714 4035 7717
rect 9990 7714 9996 7716
rect 3969 7712 9996 7714
rect 3969 7656 3974 7712
rect 4030 7656 9996 7712
rect 3969 7654 9996 7656
rect 3969 7651 4035 7654
rect 9990 7652 9996 7654
rect 10060 7652 10066 7716
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 23657 7578 23723 7581
rect 25773 7578 25839 7581
rect 23657 7576 25839 7578
rect 23657 7520 23662 7576
rect 23718 7520 25778 7576
rect 25834 7520 25839 7576
rect 23657 7518 25839 7520
rect 23657 7515 23723 7518
rect 25773 7515 25839 7518
rect 58157 7578 58223 7581
rect 59200 7578 60000 7608
rect 58157 7576 60000 7578
rect 58157 7520 58162 7576
rect 58218 7520 60000 7576
rect 58157 7518 60000 7520
rect 58157 7515 58223 7518
rect 59200 7488 60000 7518
rect 21357 7442 21423 7445
rect 28165 7442 28231 7445
rect 21357 7440 28231 7442
rect 21357 7384 21362 7440
rect 21418 7384 28170 7440
rect 28226 7384 28231 7440
rect 21357 7382 28231 7384
rect 21357 7379 21423 7382
rect 28165 7379 28231 7382
rect 9438 7108 9444 7172
rect 9508 7170 9514 7172
rect 9581 7170 9647 7173
rect 9508 7168 9647 7170
rect 9508 7112 9586 7168
rect 9642 7112 9647 7168
rect 9508 7110 9647 7112
rect 9508 7108 9514 7110
rect 9581 7107 9647 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 9489 7036 9555 7037
rect 9438 7034 9444 7036
rect 9398 6974 9444 7034
rect 9508 7032 9555 7036
rect 9550 6976 9555 7032
rect 9438 6972 9444 6974
rect 9508 6972 9555 6976
rect 9489 6971 9555 6972
rect 9990 6836 9996 6900
rect 10060 6898 10066 6900
rect 24669 6898 24735 6901
rect 10060 6896 24735 6898
rect 10060 6840 24674 6896
rect 24730 6840 24735 6896
rect 10060 6838 24735 6840
rect 10060 6836 10066 6838
rect 24669 6835 24735 6838
rect 0 6536 800 6656
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 58157 6218 58223 6221
rect 59200 6218 60000 6248
rect 58157 6216 60000 6218
rect 58157 6160 58162 6216
rect 58218 6160 60000 6216
rect 58157 6158 60000 6160
rect 58157 6155 58223 6158
rect 59200 6128 60000 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 1853 5674 1919 5677
rect 2446 5674 2452 5676
rect 1853 5672 2452 5674
rect 1853 5616 1858 5672
rect 1914 5616 2452 5672
rect 1853 5614 2452 5616
rect 1853 5611 1919 5614
rect 2446 5612 2452 5614
rect 2516 5612 2522 5676
rect 4654 5612 4660 5676
rect 4724 5674 4730 5676
rect 17309 5674 17375 5677
rect 4724 5672 17375 5674
rect 4724 5616 17314 5672
rect 17370 5616 17375 5672
rect 4724 5614 17375 5616
rect 4724 5612 4730 5614
rect 17309 5611 17375 5614
rect 29545 5674 29611 5677
rect 29913 5674 29979 5677
rect 30649 5674 30715 5677
rect 29545 5672 30715 5674
rect 29545 5616 29550 5672
rect 29606 5616 29918 5672
rect 29974 5616 30654 5672
rect 30710 5616 30715 5672
rect 29545 5614 30715 5616
rect 29545 5611 29611 5614
rect 29913 5611 29979 5614
rect 30649 5611 30715 5614
rect 0 5448 800 5568
rect 5533 5540 5599 5541
rect 5533 5536 5580 5540
rect 5644 5538 5650 5540
rect 22921 5538 22987 5541
rect 23974 5538 23980 5540
rect 5533 5480 5538 5536
rect 5533 5476 5580 5480
rect 5644 5478 5690 5538
rect 22921 5536 23980 5538
rect 22921 5480 22926 5536
rect 22982 5480 23980 5536
rect 22921 5478 23980 5480
rect 5644 5476 5650 5478
rect 5533 5475 5599 5476
rect 22921 5475 22987 5478
rect 23974 5476 23980 5478
rect 24044 5476 24050 5540
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 8334 5068 8340 5132
rect 8404 5130 8410 5132
rect 9397 5130 9463 5133
rect 29637 5130 29703 5133
rect 8404 5128 29703 5130
rect 8404 5072 9402 5128
rect 9458 5072 29642 5128
rect 29698 5072 29703 5128
rect 8404 5070 29703 5072
rect 8404 5068 8410 5070
rect 9397 5067 9463 5070
rect 29637 5067 29703 5070
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 58157 4858 58223 4861
rect 59200 4858 60000 4888
rect 58157 4856 60000 4858
rect 58157 4800 58162 4856
rect 58218 4800 60000 4856
rect 58157 4798 60000 4800
rect 58157 4795 58223 4798
rect 59200 4768 60000 4798
rect 5257 4722 5323 4725
rect 5214 4720 5323 4722
rect 5214 4664 5262 4720
rect 5318 4664 5323 4720
rect 5214 4659 5323 4664
rect 10317 4722 10383 4725
rect 12249 4722 12315 4725
rect 10317 4720 12315 4722
rect 10317 4664 10322 4720
rect 10378 4664 12254 4720
rect 12310 4664 12315 4720
rect 10317 4662 12315 4664
rect 10317 4659 10383 4662
rect 12249 4659 12315 4662
rect 5073 4586 5139 4589
rect 5214 4586 5274 4659
rect 5073 4584 5274 4586
rect 5073 4528 5078 4584
rect 5134 4528 5274 4584
rect 5073 4526 5274 4528
rect 5073 4523 5139 4526
rect 0 4360 800 4480
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 5533 4314 5599 4317
rect 7649 4314 7715 4317
rect 5533 4312 7715 4314
rect 5533 4256 5538 4312
rect 5594 4256 7654 4312
rect 7710 4256 7715 4312
rect 5533 4254 7715 4256
rect 5533 4251 5599 4254
rect 7649 4251 7715 4254
rect 5809 4178 5875 4181
rect 5398 4176 5875 4178
rect 5398 4120 5814 4176
rect 5870 4120 5875 4176
rect 5398 4118 5875 4120
rect 2589 4044 2655 4045
rect 2589 4040 2636 4044
rect 2700 4042 2706 4044
rect 5398 4042 5458 4118
rect 5809 4115 5875 4118
rect 7097 4178 7163 4181
rect 8150 4178 8156 4180
rect 7097 4176 8156 4178
rect 7097 4120 7102 4176
rect 7158 4120 8156 4176
rect 7097 4118 8156 4120
rect 7097 4115 7163 4118
rect 8150 4116 8156 4118
rect 8220 4116 8226 4180
rect 2589 3984 2594 4040
rect 2589 3980 2636 3984
rect 2700 3982 2746 4042
rect 5030 3982 5458 4042
rect 5533 4042 5599 4045
rect 8661 4044 8727 4045
rect 9489 4044 9555 4045
rect 6678 4042 6684 4044
rect 5533 4040 6684 4042
rect 5533 3984 5538 4040
rect 5594 3984 6684 4040
rect 5533 3982 6684 3984
rect 2700 3980 2706 3982
rect 2589 3979 2655 3980
rect 4889 3906 4955 3909
rect 5030 3906 5090 3982
rect 5533 3979 5599 3982
rect 6678 3980 6684 3982
rect 6748 3980 6754 4044
rect 8661 4040 8708 4044
rect 8772 4042 8778 4044
rect 8661 3984 8666 4040
rect 8661 3980 8708 3984
rect 8772 3982 8818 4042
rect 8772 3980 8778 3982
rect 9438 3980 9444 4044
rect 9508 4042 9555 4044
rect 9508 4040 9600 4042
rect 9550 3984 9600 4040
rect 9508 3982 9600 3984
rect 9508 3980 9555 3982
rect 11094 3980 11100 4044
rect 11164 4042 11170 4044
rect 11513 4042 11579 4045
rect 15837 4044 15903 4045
rect 15837 4042 15884 4044
rect 11164 4040 11579 4042
rect 11164 3984 11518 4040
rect 11574 3984 11579 4040
rect 11164 3982 11579 3984
rect 15792 4040 15884 4042
rect 15792 3984 15842 4040
rect 15792 3982 15884 3984
rect 11164 3980 11170 3982
rect 8661 3979 8727 3980
rect 9489 3979 9555 3980
rect 11513 3979 11579 3982
rect 15837 3980 15884 3982
rect 15948 3980 15954 4044
rect 15837 3979 15903 3980
rect 4662 3904 5090 3906
rect 4662 3848 4894 3904
rect 4950 3848 5090 3904
rect 4662 3846 5090 3848
rect 5257 3906 5323 3909
rect 5993 3906 6059 3909
rect 5257 3904 6059 3906
rect 5257 3848 5262 3904
rect 5318 3848 5998 3904
rect 6054 3848 6059 3904
rect 5257 3846 6059 3848
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 4662 3634 4722 3846
rect 4889 3843 4955 3846
rect 5257 3843 5323 3846
rect 5993 3843 6059 3846
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 4889 3770 4955 3773
rect 8753 3770 8819 3773
rect 20253 3772 20319 3773
rect 20253 3770 20300 3772
rect 4889 3768 8819 3770
rect 4889 3712 4894 3768
rect 4950 3712 8758 3768
rect 8814 3712 8819 3768
rect 4889 3710 8819 3712
rect 20208 3768 20300 3770
rect 20208 3712 20258 3768
rect 20208 3710 20300 3712
rect 4889 3707 4955 3710
rect 8753 3707 8819 3710
rect 20253 3708 20300 3710
rect 20364 3708 20370 3772
rect 20253 3707 20319 3708
rect 10593 3634 10659 3637
rect 2730 3632 10659 3634
rect 2730 3576 10598 3632
rect 10654 3576 10659 3632
rect 2730 3574 10659 3576
rect 2446 3436 2452 3500
rect 2516 3498 2522 3500
rect 2730 3498 2790 3574
rect 10593 3571 10659 3574
rect 2516 3438 2790 3498
rect 58157 3498 58223 3501
rect 59200 3498 60000 3528
rect 58157 3496 60000 3498
rect 58157 3440 58162 3496
rect 58218 3440 60000 3496
rect 58157 3438 60000 3440
rect 2516 3436 2522 3438
rect 58157 3435 58223 3438
rect 59200 3408 60000 3438
rect 0 3272 800 3392
rect 9857 3362 9923 3365
rect 9990 3362 9996 3364
rect 9857 3360 9996 3362
rect 9857 3304 9862 3360
rect 9918 3304 9996 3360
rect 9857 3302 9996 3304
rect 9857 3299 9923 3302
rect 9990 3300 9996 3302
rect 10060 3300 10066 3364
rect 17534 3300 17540 3364
rect 17604 3362 17610 3364
rect 18781 3362 18847 3365
rect 17604 3360 18847 3362
rect 17604 3304 18786 3360
rect 18842 3304 18847 3360
rect 17604 3302 18847 3304
rect 17604 3300 17610 3302
rect 18781 3299 18847 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 4654 3164 4660 3228
rect 4724 3226 4730 3228
rect 4889 3226 4955 3229
rect 4724 3224 4955 3226
rect 4724 3168 4894 3224
rect 4950 3168 4955 3224
rect 4724 3166 4955 3168
rect 4724 3164 4730 3166
rect 4889 3163 4955 3166
rect 8201 3226 8267 3229
rect 14089 3226 14155 3229
rect 14549 3228 14615 3229
rect 14549 3226 14596 3228
rect 8201 3224 14155 3226
rect 8201 3168 8206 3224
rect 8262 3168 14094 3224
rect 14150 3168 14155 3224
rect 8201 3166 14155 3168
rect 14504 3224 14596 3226
rect 14504 3168 14554 3224
rect 14504 3166 14596 3168
rect 8201 3163 8267 3166
rect 14089 3163 14155 3166
rect 14549 3164 14596 3166
rect 14660 3164 14666 3228
rect 15193 3226 15259 3229
rect 15326 3226 15332 3228
rect 15193 3224 15332 3226
rect 15193 3168 15198 3224
rect 15254 3168 15332 3224
rect 15193 3166 15332 3168
rect 14549 3163 14615 3164
rect 15193 3163 15259 3166
rect 15326 3164 15332 3166
rect 15396 3164 15402 3228
rect 16113 3226 16179 3229
rect 17401 3228 17467 3229
rect 16246 3226 16252 3228
rect 16113 3224 16252 3226
rect 16113 3168 16118 3224
rect 16174 3168 16252 3224
rect 16113 3166 16252 3168
rect 16113 3163 16179 3166
rect 16246 3164 16252 3166
rect 16316 3164 16322 3228
rect 17350 3164 17356 3228
rect 17420 3226 17467 3228
rect 17420 3224 17512 3226
rect 17462 3168 17512 3224
rect 17420 3166 17512 3168
rect 17420 3164 17467 3166
rect 20846 3164 20852 3228
rect 20916 3226 20922 3228
rect 20989 3226 21055 3229
rect 22369 3228 22435 3229
rect 20916 3224 21055 3226
rect 20916 3168 20994 3224
rect 21050 3168 21055 3224
rect 20916 3166 21055 3168
rect 20916 3164 20922 3166
rect 17401 3163 17467 3164
rect 20989 3163 21055 3166
rect 22318 3164 22324 3228
rect 22388 3226 22435 3228
rect 23013 3228 23079 3229
rect 23013 3226 23060 3228
rect 22388 3224 22480 3226
rect 22430 3168 22480 3224
rect 22388 3166 22480 3168
rect 22968 3224 23060 3226
rect 22968 3168 23018 3224
rect 22968 3166 23060 3168
rect 22388 3164 22435 3166
rect 22369 3163 22435 3164
rect 23013 3164 23060 3166
rect 23124 3164 23130 3228
rect 23013 3163 23079 3164
rect 2129 3090 2195 3093
rect 2589 3090 2655 3093
rect 6913 3090 6979 3093
rect 2129 3088 6979 3090
rect 2129 3032 2134 3088
rect 2190 3032 2594 3088
rect 2650 3032 6918 3088
rect 6974 3032 6979 3088
rect 2129 3030 6979 3032
rect 2129 3027 2195 3030
rect 2589 3027 2655 3030
rect 6913 3027 6979 3030
rect 8017 3090 8083 3093
rect 8661 3090 8727 3093
rect 8017 3088 8727 3090
rect 8017 3032 8022 3088
rect 8078 3032 8666 3088
rect 8722 3032 8727 3088
rect 8017 3030 8727 3032
rect 8017 3027 8083 3030
rect 8661 3027 8727 3030
rect 8937 3090 9003 3093
rect 15561 3090 15627 3093
rect 8937 3088 15627 3090
rect 8937 3032 8942 3088
rect 8998 3032 15566 3088
rect 15622 3032 15627 3088
rect 8937 3030 15627 3032
rect 8937 3027 9003 3030
rect 15561 3027 15627 3030
rect 19885 3090 19951 3093
rect 20437 3090 20503 3093
rect 19885 3088 20503 3090
rect 19885 3032 19890 3088
rect 19946 3032 20442 3088
rect 20498 3032 20503 3088
rect 19885 3030 20503 3032
rect 19885 3027 19951 3030
rect 20437 3027 20503 3030
rect 2497 2954 2563 2957
rect 6361 2954 6427 2957
rect 10961 2956 11027 2957
rect 10910 2954 10916 2956
rect 2497 2952 6427 2954
rect 2497 2896 2502 2952
rect 2558 2896 6366 2952
rect 6422 2896 6427 2952
rect 2497 2894 6427 2896
rect 10834 2894 10916 2954
rect 10980 2954 11027 2956
rect 26325 2954 26391 2957
rect 10980 2952 26391 2954
rect 11022 2896 26330 2952
rect 26386 2896 26391 2952
rect 2497 2891 2563 2894
rect 6361 2891 6427 2894
rect 10910 2892 10916 2894
rect 10980 2894 26391 2896
rect 10980 2892 11027 2894
rect 10961 2891 11027 2892
rect 26325 2891 26391 2894
rect 53373 2954 53439 2957
rect 56593 2954 56659 2957
rect 53373 2952 56659 2954
rect 53373 2896 53378 2952
rect 53434 2896 56598 2952
rect 56654 2896 56659 2952
rect 53373 2894 56659 2896
rect 53373 2891 53439 2894
rect 56593 2891 56659 2894
rect 5165 2818 5231 2821
rect 7741 2818 7807 2821
rect 5165 2816 7807 2818
rect 5165 2760 5170 2816
rect 5226 2760 7746 2816
rect 7802 2760 7807 2816
rect 5165 2758 7807 2760
rect 5165 2755 5231 2758
rect 7741 2755 7807 2758
rect 14222 2756 14228 2820
rect 14292 2818 14298 2820
rect 19793 2818 19859 2821
rect 14292 2816 19859 2818
rect 14292 2760 19798 2816
rect 19854 2760 19859 2816
rect 14292 2758 19859 2760
rect 14292 2756 14298 2758
rect 19793 2755 19859 2758
rect 53465 2818 53531 2821
rect 55305 2818 55371 2821
rect 53465 2816 55371 2818
rect 53465 2760 53470 2816
rect 53526 2760 55310 2816
rect 55366 2760 55371 2816
rect 53465 2758 55371 2760
rect 53465 2755 53531 2758
rect 55305 2755 55371 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 6545 2684 6611 2685
rect 10409 2684 10475 2685
rect 6494 2620 6500 2684
rect 6564 2682 6611 2684
rect 6564 2680 6656 2682
rect 6606 2624 6656 2680
rect 6564 2622 6656 2624
rect 6564 2620 6611 2622
rect 10358 2620 10364 2684
rect 10428 2682 10475 2684
rect 14549 2682 14615 2685
rect 17677 2684 17743 2685
rect 14774 2682 14780 2684
rect 10428 2680 10520 2682
rect 10470 2624 10520 2680
rect 10428 2622 10520 2624
rect 14549 2680 14780 2682
rect 14549 2624 14554 2680
rect 14610 2624 14780 2680
rect 14549 2622 14780 2624
rect 10428 2620 10475 2622
rect 6545 2619 6611 2620
rect 10409 2619 10475 2620
rect 14549 2619 14615 2622
rect 14774 2620 14780 2622
rect 14844 2620 14850 2684
rect 17677 2682 17724 2684
rect 17632 2680 17724 2682
rect 17632 2624 17682 2680
rect 17632 2622 17724 2624
rect 17677 2620 17724 2622
rect 17788 2620 17794 2684
rect 18638 2620 18644 2684
rect 18708 2682 18714 2684
rect 18781 2682 18847 2685
rect 21265 2684 21331 2685
rect 18708 2680 18847 2682
rect 18708 2624 18786 2680
rect 18842 2624 18847 2680
rect 18708 2622 18847 2624
rect 18708 2620 18714 2622
rect 17677 2619 17743 2620
rect 18781 2619 18847 2622
rect 21214 2620 21220 2684
rect 21284 2682 21331 2684
rect 21284 2680 21376 2682
rect 21326 2624 21376 2680
rect 21284 2622 21376 2624
rect 21284 2620 21331 2622
rect 21265 2619 21331 2620
rect 17493 2546 17559 2549
rect 23790 2546 23796 2548
rect 17493 2544 23796 2546
rect 17493 2488 17498 2544
rect 17554 2488 23796 2544
rect 17493 2486 23796 2488
rect 17493 2483 17559 2486
rect 23790 2484 23796 2486
rect 23860 2484 23866 2548
rect 6494 2348 6500 2412
rect 6564 2410 6570 2412
rect 29361 2410 29427 2413
rect 6564 2408 29427 2410
rect 6564 2352 29366 2408
rect 29422 2352 29427 2408
rect 6564 2350 29427 2352
rect 6564 2348 6570 2350
rect 29361 2347 29427 2350
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 57513 2138 57579 2141
rect 59200 2138 60000 2168
rect 57513 2136 60000 2138
rect 57513 2080 57518 2136
rect 57574 2080 60000 2136
rect 57513 2078 60000 2080
rect 57513 2075 57579 2078
rect 59200 2048 60000 2078
rect 58433 778 58499 781
rect 59200 778 60000 808
rect 58433 776 60000 778
rect 58433 720 58438 776
rect 58494 720 60000 776
rect 58433 718 60000 720
rect 58433 715 58499 718
rect 59200 688 60000 718
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 18644 56748 18708 56812
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 23980 56204 24044 56268
rect 14228 56128 14292 56132
rect 14228 56072 14242 56128
rect 14242 56072 14292 56128
rect 14228 56068 14292 56072
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 17724 55584 17788 55588
rect 17724 55528 17738 55584
rect 17738 55528 17788 55584
rect 17724 55524 17788 55528
rect 20300 55584 20364 55588
rect 20300 55528 20314 55584
rect 20314 55528 20364 55584
rect 20300 55524 20364 55528
rect 21220 55524 21284 55588
rect 22324 55524 22388 55588
rect 23796 55584 23860 55588
rect 23796 55528 23810 55584
rect 23810 55528 23860 55584
rect 23796 55524 23860 55528
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 17540 55252 17604 55316
rect 18828 55312 18892 55316
rect 18828 55256 18842 55312
rect 18842 55256 18892 55312
rect 18828 55252 18892 55256
rect 20116 55252 20180 55316
rect 21404 55252 21468 55316
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 14596 53076 14660 53140
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 14780 50220 14844 50284
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 15884 47500 15948 47564
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 15332 44780 15396 44844
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 17356 41652 17420 41716
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 23060 37844 23124 37908
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 6684 19892 6748 19956
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4660 19272 4724 19276
rect 4660 19216 4674 19272
rect 4674 19216 4724 19272
rect 4660 19212 4724 19216
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 4660 18532 4724 18596
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 5580 15132 5644 15196
rect 8708 14724 8772 14788
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 6500 13772 6564 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 11100 11052 11164 11116
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 10364 10372 10428 10436
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 16252 9964 16316 10028
rect 21404 9964 21468 10028
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 20116 9692 20180 9756
rect 20852 9692 20916 9756
rect 8340 9556 8404 9620
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 2636 8740 2700 8804
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 9444 8468 9508 8532
rect 8156 8332 8220 8396
rect 18828 8332 18892 8396
rect 10916 8196 10980 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 9996 7652 10060 7716
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 9444 7108 9508 7172
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 9444 7032 9508 7036
rect 9444 6976 9494 7032
rect 9494 6976 9508 7032
rect 9444 6972 9508 6976
rect 9996 6836 10060 6900
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 2452 5612 2516 5676
rect 4660 5612 4724 5676
rect 5580 5536 5644 5540
rect 5580 5480 5594 5536
rect 5594 5480 5644 5536
rect 5580 5476 5644 5480
rect 23980 5476 24044 5540
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 8340 5068 8404 5132
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 2636 4040 2700 4044
rect 8156 4116 8220 4180
rect 2636 3984 2650 4040
rect 2650 3984 2700 4040
rect 2636 3980 2700 3984
rect 6684 3980 6748 4044
rect 8708 4040 8772 4044
rect 8708 3984 8722 4040
rect 8722 3984 8772 4040
rect 8708 3980 8772 3984
rect 9444 4040 9508 4044
rect 9444 3984 9494 4040
rect 9494 3984 9508 4040
rect 9444 3980 9508 3984
rect 11100 3980 11164 4044
rect 15884 4040 15948 4044
rect 15884 3984 15898 4040
rect 15898 3984 15948 4040
rect 15884 3980 15948 3984
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 20300 3768 20364 3772
rect 20300 3712 20314 3768
rect 20314 3712 20364 3768
rect 20300 3708 20364 3712
rect 2452 3436 2516 3500
rect 9996 3300 10060 3364
rect 17540 3300 17604 3364
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4660 3164 4724 3228
rect 14596 3224 14660 3228
rect 14596 3168 14610 3224
rect 14610 3168 14660 3224
rect 14596 3164 14660 3168
rect 15332 3164 15396 3228
rect 16252 3164 16316 3228
rect 17356 3224 17420 3228
rect 17356 3168 17406 3224
rect 17406 3168 17420 3224
rect 17356 3164 17420 3168
rect 20852 3164 20916 3228
rect 22324 3224 22388 3228
rect 22324 3168 22374 3224
rect 22374 3168 22388 3224
rect 22324 3164 22388 3168
rect 23060 3224 23124 3228
rect 23060 3168 23074 3224
rect 23074 3168 23124 3224
rect 23060 3164 23124 3168
rect 10916 2952 10980 2956
rect 10916 2896 10966 2952
rect 10966 2896 10980 2952
rect 10916 2892 10980 2896
rect 14228 2756 14292 2820
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 6500 2680 6564 2684
rect 6500 2624 6550 2680
rect 6550 2624 6564 2680
rect 6500 2620 6564 2624
rect 10364 2680 10428 2684
rect 10364 2624 10414 2680
rect 10414 2624 10428 2680
rect 10364 2620 10428 2624
rect 14780 2620 14844 2684
rect 17724 2680 17788 2684
rect 17724 2624 17738 2680
rect 17738 2624 17788 2680
rect 17724 2620 17788 2624
rect 18644 2620 18708 2684
rect 21220 2680 21284 2684
rect 21220 2624 21270 2680
rect 21270 2624 21284 2680
rect 21220 2620 21284 2624
rect 23796 2484 23860 2548
rect 6500 2348 6564 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 18643 56812 18709 56813
rect 18643 56748 18644 56812
rect 18708 56748 18709 56812
rect 18643 56747 18709 56748
rect 14227 56132 14293 56133
rect 14227 56068 14228 56132
rect 14292 56068 14293 56132
rect 14227 56067 14293 56068
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 6683 19956 6749 19957
rect 6683 19892 6684 19956
rect 6748 19892 6749 19956
rect 6683 19891 6749 19892
rect 4659 19276 4725 19277
rect 4659 19212 4660 19276
rect 4724 19212 4725 19276
rect 4659 19211 4725 19212
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4662 18597 4722 19211
rect 4659 18596 4725 18597
rect 4659 18532 4660 18596
rect 4724 18532 4725 18596
rect 4659 18531 4725 18532
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 2635 8804 2701 8805
rect 2635 8740 2636 8804
rect 2700 8740 2701 8804
rect 2635 8739 2701 8740
rect 2451 5676 2517 5677
rect 2451 5612 2452 5676
rect 2516 5612 2517 5676
rect 2451 5611 2517 5612
rect 2454 3501 2514 5611
rect 2638 4045 2698 8739
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4662 5677 4722 18531
rect 5579 15196 5645 15197
rect 5579 15132 5580 15196
rect 5644 15132 5645 15196
rect 5579 15131 5645 15132
rect 4659 5676 4725 5677
rect 4659 5612 4660 5676
rect 4724 5612 4725 5676
rect 4659 5611 4725 5612
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 2635 4044 2701 4045
rect 2635 3980 2636 4044
rect 2700 3980 2701 4044
rect 2635 3979 2701 3980
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 2451 3500 2517 3501
rect 2451 3436 2452 3500
rect 2516 3436 2517 3500
rect 2451 3435 2517 3436
rect 4208 2752 4528 3776
rect 4662 3229 4722 5611
rect 5582 5541 5642 15131
rect 6499 13836 6565 13837
rect 6499 13772 6500 13836
rect 6564 13772 6565 13836
rect 6499 13771 6565 13772
rect 5579 5540 5645 5541
rect 5579 5476 5580 5540
rect 5644 5476 5645 5540
rect 5579 5475 5645 5476
rect 4659 3228 4725 3229
rect 4659 3164 4660 3228
rect 4724 3164 4725 3228
rect 4659 3163 4725 3164
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 6502 2685 6562 13771
rect 6686 4045 6746 19891
rect 8707 14788 8773 14789
rect 8707 14724 8708 14788
rect 8772 14724 8773 14788
rect 8707 14723 8773 14724
rect 8339 9620 8405 9621
rect 8339 9556 8340 9620
rect 8404 9556 8405 9620
rect 8339 9555 8405 9556
rect 8155 8396 8221 8397
rect 8155 8332 8156 8396
rect 8220 8332 8221 8396
rect 8155 8331 8221 8332
rect 8158 4181 8218 8331
rect 8342 5133 8402 9555
rect 8339 5132 8405 5133
rect 8339 5068 8340 5132
rect 8404 5068 8405 5132
rect 8339 5067 8405 5068
rect 8155 4180 8221 4181
rect 8155 4116 8156 4180
rect 8220 4116 8221 4180
rect 8155 4115 8221 4116
rect 8710 4045 8770 14723
rect 11099 11116 11165 11117
rect 11099 11052 11100 11116
rect 11164 11052 11165 11116
rect 11099 11051 11165 11052
rect 10363 10436 10429 10437
rect 10363 10372 10364 10436
rect 10428 10372 10429 10436
rect 10363 10371 10429 10372
rect 9443 8532 9509 8533
rect 9443 8468 9444 8532
rect 9508 8468 9509 8532
rect 9443 8467 9509 8468
rect 9446 7173 9506 8467
rect 9995 7716 10061 7717
rect 9995 7652 9996 7716
rect 10060 7652 10061 7716
rect 9995 7651 10061 7652
rect 9443 7172 9509 7173
rect 9443 7108 9444 7172
rect 9508 7108 9509 7172
rect 9443 7107 9509 7108
rect 9443 7036 9509 7037
rect 9443 6972 9444 7036
rect 9508 6972 9509 7036
rect 9443 6971 9509 6972
rect 9446 4045 9506 6971
rect 9998 6901 10058 7651
rect 9995 6900 10061 6901
rect 9995 6836 9996 6900
rect 10060 6836 10061 6900
rect 9995 6835 10061 6836
rect 6683 4044 6749 4045
rect 6683 3980 6684 4044
rect 6748 3980 6749 4044
rect 6683 3979 6749 3980
rect 8707 4044 8773 4045
rect 8707 3980 8708 4044
rect 8772 3980 8773 4044
rect 8707 3979 8773 3980
rect 9443 4044 9509 4045
rect 9443 3980 9444 4044
rect 9508 3980 9509 4044
rect 9443 3979 9509 3980
rect 9998 3365 10058 6835
rect 9995 3364 10061 3365
rect 9995 3300 9996 3364
rect 10060 3300 10061 3364
rect 9995 3299 10061 3300
rect 10366 2685 10426 10371
rect 10915 8260 10981 8261
rect 10915 8196 10916 8260
rect 10980 8196 10981 8260
rect 10915 8195 10981 8196
rect 10918 2957 10978 8195
rect 11102 4045 11162 11051
rect 11099 4044 11165 4045
rect 11099 3980 11100 4044
rect 11164 3980 11165 4044
rect 11099 3979 11165 3980
rect 10915 2956 10981 2957
rect 10915 2892 10916 2956
rect 10980 2892 10981 2956
rect 10915 2891 10981 2892
rect 14230 2821 14290 56067
rect 17723 55588 17789 55589
rect 17723 55524 17724 55588
rect 17788 55524 17789 55588
rect 17723 55523 17789 55524
rect 17539 55316 17605 55317
rect 17539 55252 17540 55316
rect 17604 55252 17605 55316
rect 17539 55251 17605 55252
rect 14595 53140 14661 53141
rect 14595 53076 14596 53140
rect 14660 53076 14661 53140
rect 14595 53075 14661 53076
rect 14598 3229 14658 53075
rect 14779 50284 14845 50285
rect 14779 50220 14780 50284
rect 14844 50220 14845 50284
rect 14779 50219 14845 50220
rect 14595 3228 14661 3229
rect 14595 3164 14596 3228
rect 14660 3164 14661 3228
rect 14595 3163 14661 3164
rect 14227 2820 14293 2821
rect 14227 2756 14228 2820
rect 14292 2756 14293 2820
rect 14227 2755 14293 2756
rect 14782 2685 14842 50219
rect 15883 47564 15949 47565
rect 15883 47500 15884 47564
rect 15948 47500 15949 47564
rect 15883 47499 15949 47500
rect 15331 44844 15397 44845
rect 15331 44780 15332 44844
rect 15396 44780 15397 44844
rect 15331 44779 15397 44780
rect 15334 3229 15394 44779
rect 15886 4045 15946 47499
rect 17355 41716 17421 41717
rect 17355 41652 17356 41716
rect 17420 41652 17421 41716
rect 17355 41651 17421 41652
rect 16251 10028 16317 10029
rect 16251 9964 16252 10028
rect 16316 9964 16317 10028
rect 16251 9963 16317 9964
rect 15883 4044 15949 4045
rect 15883 3980 15884 4044
rect 15948 3980 15949 4044
rect 15883 3979 15949 3980
rect 16254 3229 16314 9963
rect 17358 3229 17418 41651
rect 17542 3365 17602 55251
rect 17539 3364 17605 3365
rect 17539 3300 17540 3364
rect 17604 3300 17605 3364
rect 17539 3299 17605 3300
rect 15331 3228 15397 3229
rect 15331 3164 15332 3228
rect 15396 3164 15397 3228
rect 15331 3163 15397 3164
rect 16251 3228 16317 3229
rect 16251 3164 16252 3228
rect 16316 3164 16317 3228
rect 16251 3163 16317 3164
rect 17355 3228 17421 3229
rect 17355 3164 17356 3228
rect 17420 3164 17421 3228
rect 17355 3163 17421 3164
rect 17726 2685 17786 55523
rect 18646 2685 18706 56747
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 23979 56268 24045 56269
rect 23979 56204 23980 56268
rect 24044 56204 24045 56268
rect 23979 56203 24045 56204
rect 20299 55588 20365 55589
rect 20299 55524 20300 55588
rect 20364 55524 20365 55588
rect 20299 55523 20365 55524
rect 21219 55588 21285 55589
rect 21219 55524 21220 55588
rect 21284 55524 21285 55588
rect 21219 55523 21285 55524
rect 22323 55588 22389 55589
rect 22323 55524 22324 55588
rect 22388 55524 22389 55588
rect 22323 55523 22389 55524
rect 23795 55588 23861 55589
rect 23795 55524 23796 55588
rect 23860 55524 23861 55588
rect 23795 55523 23861 55524
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 18827 55316 18893 55317
rect 18827 55252 18828 55316
rect 18892 55252 18893 55316
rect 18827 55251 18893 55252
rect 18830 8397 18890 55251
rect 19568 54432 19888 55456
rect 20115 55316 20181 55317
rect 20115 55252 20116 55316
rect 20180 55252 20181 55316
rect 20115 55251 20181 55252
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 20118 9757 20178 55251
rect 20115 9756 20181 9757
rect 20115 9692 20116 9756
rect 20180 9692 20181 9756
rect 20115 9691 20181 9692
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 18827 8396 18893 8397
rect 18827 8332 18828 8396
rect 18892 8332 18893 8396
rect 18827 8331 18893 8332
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 20302 3773 20362 55523
rect 20851 9756 20917 9757
rect 20851 9692 20852 9756
rect 20916 9692 20917 9756
rect 20851 9691 20917 9692
rect 20299 3772 20365 3773
rect 20299 3708 20300 3772
rect 20364 3708 20365 3772
rect 20299 3707 20365 3708
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 6499 2684 6565 2685
rect 6499 2620 6500 2684
rect 6564 2620 6565 2684
rect 6499 2619 6565 2620
rect 10363 2684 10429 2685
rect 10363 2620 10364 2684
rect 10428 2620 10429 2684
rect 10363 2619 10429 2620
rect 14779 2684 14845 2685
rect 14779 2620 14780 2684
rect 14844 2620 14845 2684
rect 14779 2619 14845 2620
rect 17723 2684 17789 2685
rect 17723 2620 17724 2684
rect 17788 2620 17789 2684
rect 17723 2619 17789 2620
rect 18643 2684 18709 2685
rect 18643 2620 18644 2684
rect 18708 2620 18709 2684
rect 18643 2619 18709 2620
rect 6502 2413 6562 2619
rect 6499 2412 6565 2413
rect 6499 2348 6500 2412
rect 6564 2348 6565 2412
rect 6499 2347 6565 2348
rect 19568 2208 19888 3232
rect 20854 3229 20914 9691
rect 20851 3228 20917 3229
rect 20851 3164 20852 3228
rect 20916 3164 20917 3228
rect 20851 3163 20917 3164
rect 21222 2685 21282 55523
rect 21403 55316 21469 55317
rect 21403 55252 21404 55316
rect 21468 55252 21469 55316
rect 21403 55251 21469 55252
rect 21406 10029 21466 55251
rect 21403 10028 21469 10029
rect 21403 9964 21404 10028
rect 21468 9964 21469 10028
rect 21403 9963 21469 9964
rect 22326 3229 22386 55523
rect 23059 37908 23125 37909
rect 23059 37844 23060 37908
rect 23124 37844 23125 37908
rect 23059 37843 23125 37844
rect 23062 3229 23122 37843
rect 22323 3228 22389 3229
rect 22323 3164 22324 3228
rect 22388 3164 22389 3228
rect 22323 3163 22389 3164
rect 23059 3228 23125 3229
rect 23059 3164 23060 3228
rect 23124 3164 23125 3228
rect 23059 3163 23125 3164
rect 21219 2684 21285 2685
rect 21219 2620 21220 2684
rect 21284 2620 21285 2684
rect 21219 2619 21285 2620
rect 23798 2549 23858 55523
rect 23982 5541 24042 56203
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 23979 5540 24045 5541
rect 23979 5476 23980 5540
rect 24044 5476 24045 5540
rect 23979 5475 24045 5476
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 23795 2548 23861 2549
rect 23795 2484 23796 2548
rect 23860 2484 23861 2548
rect 23795 2483 23861 2484
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10120 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__B
timestamp 1649977179
transform 1 0 9568 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A0
timestamp 1649977179
transform -1 0 4416 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A0
timestamp 1649977179
transform 1 0 4416 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A0
timestamp 1649977179
transform -1 0 1840 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A0
timestamp 1649977179
transform 1 0 4048 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A0
timestamp 1649977179
transform 1 0 4600 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A0
timestamp 1649977179
transform 1 0 5428 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__A0
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A0
timestamp 1649977179
transform 1 0 10120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A0
timestamp 1649977179
transform 1 0 3864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A0
timestamp 1649977179
transform 1 0 12420 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A0
timestamp 1649977179
transform 1 0 3312 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A0
timestamp 1649977179
transform 1 0 8648 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__A
timestamp 1649977179
transform 1 0 5704 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A
timestamp 1649977179
transform -1 0 7728 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A
timestamp 1649977179
transform -1 0 17572 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A
timestamp 1649977179
transform -1 0 13340 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__B
timestamp 1649977179
transform -1 0 12236 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A
timestamp 1649977179
transform 1 0 8372 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A
timestamp 1649977179
transform 1 0 11592 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A
timestamp 1649977179
transform 1 0 8556 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A1
timestamp 1649977179
transform -1 0 5060 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A
timestamp 1649977179
transform 1 0 4508 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A1
timestamp 1649977179
transform 1 0 5336 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A
timestamp 1649977179
transform 1 0 5704 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A1
timestamp 1649977179
transform 1 0 3864 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A
timestamp 1649977179
transform 1 0 8372 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A1
timestamp 1649977179
transform -1 0 7360 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A
timestamp 1649977179
transform 1 0 12144 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A1
timestamp 1649977179
transform 1 0 7452 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A
timestamp 1649977179
transform 1 0 24564 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A
timestamp 1649977179
transform -1 0 14812 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A1
timestamp 1649977179
transform -1 0 13616 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A
timestamp 1649977179
transform -1 0 26220 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A1
timestamp 1649977179
transform -1 0 17848 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__A
timestamp 1649977179
transform 1 0 23368 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A1
timestamp 1649977179
transform -1 0 16744 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A1
timestamp 1649977179
transform 1 0 15640 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A
timestamp 1649977179
transform 1 0 24196 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A1
timestamp 1649977179
transform -1 0 15364 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A
timestamp 1649977179
transform 1 0 16100 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A1
timestamp 1649977179
transform 1 0 15180 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__C1
timestamp 1649977179
transform 1 0 13892 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A1
timestamp 1649977179
transform 1 0 13800 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__C1
timestamp 1649977179
transform -1 0 12972 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__A
timestamp 1649977179
transform 1 0 20056 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__B
timestamp 1649977179
transform -1 0 20424 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__A
timestamp 1649977179
transform -1 0 29992 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A
timestamp 1649977179
transform 1 0 28888 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A
timestamp 1649977179
transform 1 0 29348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A1
timestamp 1649977179
transform -1 0 29716 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__C1
timestamp 1649977179
transform -1 0 29072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A1
timestamp 1649977179
transform 1 0 26956 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__C1
timestamp 1649977179
transform 1 0 27140 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A1
timestamp 1649977179
transform 1 0 26312 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__C1
timestamp 1649977179
transform 1 0 27600 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A
timestamp 1649977179
transform 1 0 28888 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A1
timestamp 1649977179
transform 1 0 28520 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A1
timestamp 1649977179
transform 1 0 29532 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A1
timestamp 1649977179
transform 1 0 35420 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A1
timestamp 1649977179
transform -1 0 37260 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A1
timestamp 1649977179
transform -1 0 37444 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A
timestamp 1649977179
transform 1 0 28888 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A1
timestamp 1649977179
transform -1 0 36616 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A1
timestamp 1649977179
transform -1 0 35696 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A1
timestamp 1649977179
transform -1 0 35972 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A1
timestamp 1649977179
transform -1 0 32752 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A
timestamp 1649977179
transform 1 0 19872 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__B
timestamp 1649977179
transform -1 0 20976 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A
timestamp 1649977179
transform -1 0 31648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A
timestamp 1649977179
transform -1 0 31188 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A
timestamp 1649977179
transform -1 0 32752 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A1
timestamp 1649977179
transform 1 0 27784 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A
timestamp 1649977179
transform 1 0 30360 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A1
timestamp 1649977179
transform 1 0 27048 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A1
timestamp 1649977179
transform 1 0 26956 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A1
timestamp 1649977179
transform -1 0 31556 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A1
timestamp 1649977179
transform 1 0 30268 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A1
timestamp 1649977179
transform 1 0 33212 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A
timestamp 1649977179
transform 1 0 31372 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A1
timestamp 1649977179
transform 1 0 33212 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A1
timestamp 1649977179
transform 1 0 33580 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A1
timestamp 1649977179
transform 1 0 34132 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A1
timestamp 1649977179
transform 1 0 34500 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A1
timestamp 1649977179
transform 1 0 32016 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A
timestamp 1649977179
transform 1 0 29716 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A1
timestamp 1649977179
transform 1 0 31832 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__C1
timestamp 1649977179
transform 1 0 31464 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A
timestamp 1649977179
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B
timestamp 1649977179
transform 1 0 8832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A
timestamp 1649977179
transform 1 0 7820 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A
timestamp 1649977179
transform 1 0 16836 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A1
timestamp 1649977179
transform 1 0 5520 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__C1
timestamp 1649977179
transform 1 0 5060 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__A1
timestamp 1649977179
transform 1 0 5244 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__C1
timestamp 1649977179
transform 1 0 5704 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A1
timestamp 1649977179
transform 1 0 5336 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__C1
timestamp 1649977179
transform 1 0 5520 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A1
timestamp 1649977179
transform 1 0 8188 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__C1
timestamp 1649977179
transform -1 0 7452 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A
timestamp 1649977179
transform 1 0 19872 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A1
timestamp 1649977179
transform 1 0 7820 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__C1
timestamp 1649977179
transform 1 0 8280 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A1
timestamp 1649977179
transform 1 0 20884 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__C1
timestamp 1649977179
transform 1 0 19228 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A1
timestamp 1649977179
transform 1 0 18492 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__C1
timestamp 1649977179
transform 1 0 18584 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A1
timestamp 1649977179
transform 1 0 20792 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__C1
timestamp 1649977179
transform -1 0 20240 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A1
timestamp 1649977179
transform 1 0 20700 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__C1
timestamp 1649977179
transform 1 0 19412 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__A
timestamp 1649977179
transform -1 0 17940 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A1
timestamp 1649977179
transform 1 0 17664 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A1
timestamp 1649977179
transform 1 0 15732 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A1
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A
timestamp 1649977179
transform -1 0 19412 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__B
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A
timestamp 1649977179
transform 1 0 17112 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1649977179
transform -1 0 16376 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A1
timestamp 1649977179
transform 1 0 10028 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A1
timestamp 1649977179
transform 1 0 9200 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A
timestamp 1649977179
transform 1 0 23276 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A1
timestamp 1649977179
transform 1 0 10856 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__C1
timestamp 1649977179
transform -1 0 11684 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__A1
timestamp 1649977179
transform 1 0 12052 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__C1
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A1
timestamp 1649977179
transform 1 0 13800 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__C1
timestamp 1649977179
transform -1 0 14536 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__A1
timestamp 1649977179
transform 1 0 25576 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__C1
timestamp 1649977179
transform -1 0 24564 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A1
timestamp 1649977179
transform 1 0 25484 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__C1
timestamp 1649977179
transform 1 0 23736 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__A
timestamp 1649977179
transform -1 0 25484 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__A1
timestamp 1649977179
transform 1 0 23828 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__A1
timestamp 1649977179
transform 1 0 25760 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A1
timestamp 1649977179
transform 1 0 24656 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__A1
timestamp 1649977179
transform 1 0 26220 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__A1
timestamp 1649977179
transform 1 0 23736 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__A
timestamp 1649977179
transform 1 0 14352 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__A
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A
timestamp 1649977179
transform 1 0 20884 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__B
timestamp 1649977179
transform 1 0 20700 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A
timestamp 1649977179
transform 1 0 23276 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A
timestamp 1649977179
transform 1 0 21252 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A
timestamp 1649977179
transform -1 0 25116 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A1
timestamp 1649977179
transform 1 0 23276 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__A
timestamp 1649977179
transform 1 0 15548 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__A1
timestamp 1649977179
transform -1 0 24564 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__A
timestamp 1649977179
transform 1 0 13432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__A1
timestamp 1649977179
transform -1 0 23736 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A
timestamp 1649977179
transform -1 0 19504 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__A1
timestamp 1649977179
transform -1 0 24288 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__A
timestamp 1649977179
transform 1 0 17756 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__A1
timestamp 1649977179
transform 1 0 23736 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A
timestamp 1649977179
transform 1 0 28520 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A
timestamp 1649977179
transform 1 0 32844 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__A1
timestamp 1649977179
transform 1 0 29808 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A
timestamp 1649977179
transform 1 0 29624 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__A1
timestamp 1649977179
transform -1 0 31648 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A
timestamp 1649977179
transform 1 0 28980 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A1
timestamp 1649977179
transform 1 0 30728 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A
timestamp 1649977179
transform 1 0 27232 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__A1
timestamp 1649977179
transform -1 0 33396 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__A
timestamp 1649977179
transform 1 0 26680 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__A1
timestamp 1649977179
transform -1 0 29992 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__A
timestamp 1649977179
transform 1 0 18584 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__A1
timestamp 1649977179
transform 1 0 21988 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__A
timestamp 1649977179
transform 1 0 18952 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__A1
timestamp 1649977179
transform -1 0 25208 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__A
timestamp 1649977179
transform 1 0 19596 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__B
timestamp 1649977179
transform 1 0 18308 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__A
timestamp 1649977179
transform 1 0 21160 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__A
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__A1
timestamp 1649977179
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A1
timestamp 1649977179
transform 1 0 15456 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__A1
timestamp 1649977179
transform 1 0 15272 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__A1
timestamp 1649977179
transform 1 0 19596 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__C1
timestamp 1649977179
transform 1 0 20424 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__A1
timestamp 1649977179
transform 1 0 19504 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__C1
timestamp 1649977179
transform -1 0 17664 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A1
timestamp 1649977179
transform -1 0 27968 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__C1
timestamp 1649977179
transform -1 0 27416 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__A1
timestamp 1649977179
transform 1 0 31188 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__C1
timestamp 1649977179
transform -1 0 29716 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A1
timestamp 1649977179
transform 1 0 30544 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__C1
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__A1
timestamp 1649977179
transform -1 0 27692 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__C1
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__A1
timestamp 1649977179
transform -1 0 25392 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__C1
timestamp 1649977179
transform 1 0 27416 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__A1
timestamp 1649977179
transform 1 0 21344 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__C1
timestamp 1649977179
transform 1 0 22632 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A1
timestamp 1649977179
transform 1 0 21160 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__C1
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__A
timestamp 1649977179
transform -1 0 24472 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__B
timestamp 1649977179
transform -1 0 23460 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__A
timestamp 1649977179
transform 1 0 34868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A
timestamp 1649977179
transform 1 0 33212 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__A1
timestamp 1649977179
transform 1 0 34592 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__C1
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__A1
timestamp 1649977179
transform -1 0 40020 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__C1
timestamp 1649977179
transform 1 0 37996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__A1
timestamp 1649977179
transform -1 0 37904 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__C1
timestamp 1649977179
transform -1 0 36432 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__A1
timestamp 1649977179
transform -1 0 39192 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__C1
timestamp 1649977179
transform 1 0 36800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__A1
timestamp 1649977179
transform 1 0 38180 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__C1
timestamp 1649977179
transform -1 0 40020 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__A1
timestamp 1649977179
transform 1 0 37444 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__C1
timestamp 1649977179
transform 1 0 36892 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__A
timestamp 1649977179
transform -1 0 34868 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__A1
timestamp 1649977179
transform 1 0 39192 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__A1
timestamp 1649977179
transform -1 0 41860 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__A1
timestamp 1649977179
transform 1 0 39928 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__A1
timestamp 1649977179
transform 1 0 40664 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__A1
timestamp 1649977179
transform -1 0 41124 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A1
timestamp 1649977179
transform 1 0 35420 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__A
timestamp 1649977179
transform 1 0 21160 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__B
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__A
timestamp 1649977179
transform 1 0 34500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__A
timestamp 1649977179
transform -1 0 36800 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__A1
timestamp 1649977179
transform -1 0 34592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__A1
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__A1
timestamp 1649977179
transform 1 0 33764 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A1
timestamp 1649977179
transform 1 0 36616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__A1
timestamp 1649977179
transform -1 0 40020 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__A1
timestamp 1649977179
transform -1 0 37444 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__A1
timestamp 1649977179
transform -1 0 39376 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__A1
timestamp 1649977179
transform 1 0 41124 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__A1
timestamp 1649977179
transform -1 0 40388 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__A1
timestamp 1649977179
transform -1 0 41400 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__C1
timestamp 1649977179
transform -1 0 41676 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A1
timestamp 1649977179
transform 1 0 38272 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__C1
timestamp 1649977179
transform 1 0 38824 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__A1
timestamp 1649977179
transform 1 0 35512 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__C1
timestamp 1649977179
transform 1 0 36248 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__A
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__B
timestamp 1649977179
transform -1 0 24564 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__A
timestamp 1649977179
transform -1 0 28152 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__A
timestamp 1649977179
transform 1 0 27232 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__A1
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__C1
timestamp 1649977179
transform 1 0 28060 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__A1
timestamp 1649977179
transform -1 0 26588 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__C1
timestamp 1649977179
transform -1 0 27876 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A1
timestamp 1649977179
transform 1 0 29072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__A1
timestamp 1649977179
transform 1 0 28336 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__A1
timestamp 1649977179
transform 1 0 29072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__A1
timestamp 1649977179
transform 1 0 33856 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1282__A1
timestamp 1649977179
transform 1 0 31464 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__A
timestamp 1649977179
transform 1 0 14352 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__A
timestamp 1649977179
transform 1 0 23736 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__A1
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__A1
timestamp 1649977179
transform 1 0 32292 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__A1
timestamp 1649977179
transform 1 0 31556 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__A1
timestamp 1649977179
transform 1 0 25484 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__A1
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__A
timestamp 1649977179
transform 1 0 5152 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__A
timestamp 1649977179
transform 1 0 20332 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__A
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__B
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__A
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__A
timestamp 1649977179
transform 1 0 7912 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__A
timestamp 1649977179
transform -1 0 16008 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__A
timestamp 1649977179
transform 1 0 7820 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__A
timestamp 1649977179
transform 1 0 7268 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__A1
timestamp 1649977179
transform 1 0 4784 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__A
timestamp 1649977179
transform 1 0 3128 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__A1
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__A
timestamp 1649977179
transform 1 0 4416 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__A1
timestamp 1649977179
transform 1 0 2944 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__A
timestamp 1649977179
transform 1 0 5704 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__A1
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__A
timestamp 1649977179
transform 1 0 5888 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__A1
timestamp 1649977179
transform 1 0 5704 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__A
timestamp 1649977179
transform -1 0 22172 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__A
timestamp 1649977179
transform 1 0 20884 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__A
timestamp 1649977179
transform -1 0 20424 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__A
timestamp 1649977179
transform -1 0 21620 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__A1
timestamp 1649977179
transform -1 0 22724 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__A
timestamp 1649977179
transform 1 0 25116 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__A1
timestamp 1649977179
transform 1 0 23184 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__A
timestamp 1649977179
transform 1 0 26128 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__A1
timestamp 1649977179
transform 1 0 23736 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__A
timestamp 1649977179
transform 1 0 15548 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__A1
timestamp 1649977179
transform 1 0 21712 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__A
timestamp 1649977179
transform -1 0 17020 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__A1
timestamp 1649977179
transform -1 0 22264 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__A
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__B
timestamp 1649977179
transform 1 0 19320 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__A
timestamp 1649977179
transform 1 0 17756 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__A1
timestamp 1649977179
transform 1 0 17388 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__A2
timestamp 1649977179
transform 1 0 17480 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__A
timestamp 1649977179
transform 1 0 8924 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1341__B
timestamp 1649977179
transform -1 0 21896 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__A1
timestamp 1649977179
transform 1 0 18768 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__A2
timestamp 1649977179
transform -1 0 19412 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__A
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__B
timestamp 1649977179
transform 1 0 21988 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__A
timestamp 1649977179
transform -1 0 22724 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__A
timestamp 1649977179
transform -1 0 22816 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__A1
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__A1
timestamp 1649977179
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__A1
timestamp 1649977179
transform 1 0 14812 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__A
timestamp 1649977179
transform 1 0 16652 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__A1
timestamp 1649977179
transform 1 0 15824 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__A1
timestamp 1649977179
transform 1 0 17480 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1365__A1
timestamp 1649977179
transform -1 0 24656 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__A1
timestamp 1649977179
transform -1 0 25208 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__A1
timestamp 1649977179
transform -1 0 27140 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__A
timestamp 1649977179
transform 1 0 12972 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__A1
timestamp 1649977179
transform 1 0 24196 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__C1
timestamp 1649977179
transform -1 0 24564 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__A1
timestamp 1649977179
transform 1 0 25576 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__C1
timestamp 1649977179
transform 1 0 26128 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__A1
timestamp 1649977179
transform 1 0 22632 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__C1
timestamp 1649977179
transform 1 0 23184 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__A1
timestamp 1649977179
transform -1 0 22264 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__C1
timestamp 1649977179
transform -1 0 22080 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__A
timestamp 1649977179
transform 1 0 10212 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__B
timestamp 1649977179
transform 1 0 9384 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__A
timestamp 1649977179
transform -1 0 9384 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__A
timestamp 1649977179
transform 1 0 12420 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__A1
timestamp 1649977179
transform 1 0 7176 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__C1
timestamp 1649977179
transform -1 0 8464 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__A1
timestamp 1649977179
transform 1 0 5244 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__C1
timestamp 1649977179
transform -1 0 4876 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__A1
timestamp 1649977179
transform 1 0 4508 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__C1
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__A1
timestamp 1649977179
transform 1 0 7176 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__C1
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__A1
timestamp 1649977179
transform 1 0 6164 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__C1
timestamp 1649977179
transform 1 0 7452 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__A1
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__C1
timestamp 1649977179
transform 1 0 13892 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__A1
timestamp 1649977179
transform 1 0 16192 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1406__A1
timestamp 1649977179
transform 1 0 18584 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1408__A1
timestamp 1649977179
transform 1 0 16008 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__A1
timestamp 1649977179
transform 1 0 18400 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__A1
timestamp 1649977179
transform 1 0 15364 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__A1
timestamp 1649977179
transform -1 0 10028 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__A
timestamp 1649977179
transform 1 0 10856 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__B
timestamp 1649977179
transform -1 0 10580 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1418__A
timestamp 1649977179
transform 1 0 9844 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1420__A
timestamp 1649977179
transform 1 0 11776 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__A1
timestamp 1649977179
transform 1 0 3588 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__A1
timestamp 1649977179
transform 1 0 2852 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__A1
timestamp 1649977179
transform 1 0 3220 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__A1
timestamp 1649977179
transform -1 0 5336 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__A1
timestamp 1649977179
transform -1 0 6624 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__A1
timestamp 1649977179
transform 1 0 12512 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__A1
timestamp 1649977179
transform -1 0 10488 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__A1
timestamp 1649977179
transform 1 0 11500 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__A1
timestamp 1649977179
transform 1 0 11500 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__A
timestamp 1649977179
transform -1 0 10304 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__A1
timestamp 1649977179
transform 1 0 12328 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__C1
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__A1
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__C1
timestamp 1649977179
transform 1 0 11040 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__A1
timestamp 1649977179
transform -1 0 9108 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__C1
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__A
timestamp 1649977179
transform 1 0 13892 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__B
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1453__A
timestamp 1649977179
transform -1 0 14812 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__A
timestamp 1649977179
transform 1 0 14812 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__A1
timestamp 1649977179
transform 1 0 9200 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__C1
timestamp 1649977179
transform -1 0 9936 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__A1
timestamp 1649977179
transform 1 0 10856 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__C1
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__A
timestamp 1649977179
transform 1 0 14076 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1464__A1
timestamp 1649977179
transform 1 0 12604 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1466__A1
timestamp 1649977179
transform -1 0 12788 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1468__A1
timestamp 1649977179
transform 1 0 11960 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__A1
timestamp 1649977179
transform -1 0 18860 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1474__A1
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1476__A
timestamp 1649977179
transform 1 0 19780 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1477__A1
timestamp 1649977179
transform -1 0 23828 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1479__A1
timestamp 1649977179
transform -1 0 21344 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__A1
timestamp 1649977179
transform 1 0 17664 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__A1
timestamp 1649977179
transform 1 0 16468 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__A1
timestamp 1649977179
transform 1 0 17664 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1487__A
timestamp 1649977179
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1489__A
timestamp 1649977179
transform 1 0 20608 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1491__A
timestamp 1649977179
transform -1 0 20516 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__A
timestamp 1649977179
transform 1 0 16468 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__A1
timestamp 1649977179
transform 1 0 14812 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__A1
timestamp 1649977179
transform 1 0 13432 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1499__A1
timestamp 1649977179
transform 1 0 14260 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1501__A1
timestamp 1649977179
transform 1 0 18032 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__A1
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1507__A
timestamp 1649977179
transform -1 0 26956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1508__A1
timestamp 1649977179
transform 1 0 29624 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1510__A1
timestamp 1649977179
transform 1 0 29624 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1512__A1
timestamp 1649977179
transform 1 0 29716 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1514__A1
timestamp 1649977179
transform 1 0 26864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1516__A1
timestamp 1649977179
transform 1 0 26312 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1519__A1
timestamp 1649977179
transform 1 0 17480 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1519__C1
timestamp 1649977179
transform 1 0 17112 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__A1
timestamp 1649977179
transform 1 0 16928 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__C1
timestamp 1649977179
transform 1 0 17480 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1535__D
timestamp 1649977179
transform -1 0 25484 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1541__C1
timestamp 1649977179
transform 1 0 6900 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1546__A
timestamp 1649977179
transform -1 0 23920 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1546__D
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1554__C1
timestamp 1649977179
transform 1 0 7452 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1559__D
timestamp 1649977179
transform -1 0 23736 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1567__C1
timestamp 1649977179
transform -1 0 7820 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1583__A
timestamp 1649977179
transform 1 0 30176 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1585__A
timestamp 1649977179
transform -1 0 32292 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1599__A2
timestamp 1649977179
transform -1 0 16836 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1599__B1
timestamp 1649977179
transform -1 0 15456 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1601__A
timestamp 1649977179
transform 1 0 9108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1604__A1
timestamp 1649977179
transform -1 0 8280 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1616__A2
timestamp 1649977179
transform 1 0 15548 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1616__B1
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1618__A
timestamp 1649977179
transform 1 0 10028 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1620__A1
timestamp 1649977179
transform -1 0 6624 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1629__A2
timestamp 1649977179
transform 1 0 22356 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1629__B1
timestamp 1649977179
transform 1 0 22908 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1633__B1
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1641__A2
timestamp 1649977179
transform 1 0 22080 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1641__B1
timestamp 1649977179
transform -1 0 23460 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1646__B1
timestamp 1649977179
transform 1 0 10396 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1654__A2
timestamp 1649977179
transform -1 0 22448 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1654__B1
timestamp 1649977179
transform -1 0 24564 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1659__B1
timestamp 1649977179
transform -1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1671__B1
timestamp 1649977179
transform -1 0 12880 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1688__D
timestamp 1649977179
transform -1 0 25116 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1695__B1
timestamp 1649977179
transform 1 0 5704 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1708__A
timestamp 1649977179
transform -1 0 1932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2176__A
timestamp 1649977179
transform -1 0 46920 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2177__A
timestamp 1649977179
transform 1 0 21712 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2178__A
timestamp 1649977179
transform -1 0 44620 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2179__A
timestamp 1649977179
transform -1 0 20148 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2180__A
timestamp 1649977179
transform 1 0 18768 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2181__A
timestamp 1649977179
transform -1 0 18768 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2182__A
timestamp 1649977179
transform -1 0 17112 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2183__A
timestamp 1649977179
transform 1 0 19688 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2184__A
timestamp 1649977179
transform -1 0 20792 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2185__A
timestamp 1649977179
transform 1 0 24380 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2186__A
timestamp 1649977179
transform -1 0 29716 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2187__A
timestamp 1649977179
transform -1 0 32936 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2188__A
timestamp 1649977179
transform 1 0 30912 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2189__A
timestamp 1649977179
transform 1 0 27968 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2190__A
timestamp 1649977179
transform 1 0 24932 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2191__A
timestamp 1649977179
transform 1 0 26772 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2192__A
timestamp 1649977179
transform 1 0 26036 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2193__A
timestamp 1649977179
transform 1 0 23644 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2194__A
timestamp 1649977179
transform 1 0 22356 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2195__A
timestamp 1649977179
transform 1 0 20884 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2196__A
timestamp 1649977179
transform -1 0 18124 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2197__A
timestamp 1649977179
transform -1 0 17572 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2198__A
timestamp 1649977179
transform -1 0 17112 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2199__A
timestamp 1649977179
transform 1 0 17756 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2200__A
timestamp 1649977179
transform 1 0 16008 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2201__A
timestamp 1649977179
transform 1 0 14168 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2202__A
timestamp 1649977179
transform -1 0 20424 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2203__A
timestamp 1649977179
transform 1 0 23000 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2204__A
timestamp 1649977179
transform 1 0 29900 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2205__A
timestamp 1649977179
transform -1 0 36340 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 20332 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_wb_clk_i_A
timestamp 1649977179
transform 1 0 12972 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_wb_clk_i_A
timestamp 1649977179
transform 1 0 10028 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_wb_clk_i_A
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_wb_clk_i_A
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_wb_clk_i_A
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_wb_clk_i_A
timestamp 1649977179
transform -1 0 12696 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_wb_clk_i_A
timestamp 1649977179
transform 1 0 14444 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_wb_clk_i_A
timestamp 1649977179
transform 1 0 8648 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_5_wb_clk_i_A
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_wb_clk_i_A
timestamp 1649977179
transform 1 0 8096 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_wb_clk_i_A
timestamp 1649977179
transform 1 0 5336 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_wb_clk_i_A
timestamp 1649977179
transform 1 0 9108 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_wb_clk_i_A
timestamp 1649977179
transform -1 0 17020 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_wb_clk_i_A
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_11_wb_clk_i_A
timestamp 1649977179
transform 1 0 23184 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_12_wb_clk_i_A
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_13_wb_clk_i_A
timestamp 1649977179
transform 1 0 25852 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_14_wb_clk_i_A
timestamp 1649977179
transform -1 0 29808 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_15_wb_clk_i_A
timestamp 1649977179
transform 1 0 32200 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_16_wb_clk_i_A
timestamp 1649977179
transform 1 0 37444 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_17_wb_clk_i_A
timestamp 1649977179
transform 1 0 38088 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_18_wb_clk_i_A
timestamp 1649977179
transform 1 0 30820 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_19_wb_clk_i_A
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_20_wb_clk_i_A
timestamp 1649977179
transform 1 0 32292 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_21_wb_clk_i_A
timestamp 1649977179
transform 1 0 37444 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_22_wb_clk_i_A
timestamp 1649977179
transform 1 0 37536 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_23_wb_clk_i_A
timestamp 1649977179
transform 1 0 37352 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_24_wb_clk_i_A
timestamp 1649977179
transform 1 0 36524 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_25_wb_clk_i_A
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_26_wb_clk_i_A
timestamp 1649977179
transform 1 0 26036 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_27_wb_clk_i_A
timestamp 1649977179
transform 1 0 25852 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_28_wb_clk_i_A
timestamp 1649977179
transform 1 0 16008 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_29_wb_clk_i_A
timestamp 1649977179
transform 1 0 16744 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_30_wb_clk_i_A
timestamp 1649977179
transform 1 0 13800 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_31_wb_clk_i_A
timestamp 1649977179
transform 1 0 4324 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 16928 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 17480 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 21160 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 26404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 19412 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 20608 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 20056 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 20240 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 25300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 20792 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 10304 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 18032 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 21344 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 21528 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 21988 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 22080 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 23184 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 23736 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 22632 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 27140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 24564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 13064 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 12512 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 15824 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 16376 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 16744 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 13616 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 25852 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 1840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 6532 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 11960 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 11408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 3312 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 13892 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 10120 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 7268 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 7820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 2116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 1748 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 9384 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 4508 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 1840 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 9936 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 5060 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 1564 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 2300 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 5612 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 1748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 7820 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 10856 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 10212 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 2024 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 10488 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 2852 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 4324 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 1840 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output61_A
timestamp 1649977179
transform 1 0 40756 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output68_A
timestamp 1649977179
transform 1 0 2576 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output87_A
timestamp 1649977179
transform 1 0 42320 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output96_A
timestamp 1649977179
transform 1 0 3128 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output97_A
timestamp 1649977179
transform -1 0 4232 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16
timestamp 1649977179
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1649977179
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1649977179
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1649977179
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_89 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103
timestamp 1649977179
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1649977179
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1649977179
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131
timestamp 1649977179
transform 1 0 13156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1649977179
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_148
timestamp 1649977179
transform 1 0 14720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1649977179
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1649977179
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_173
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_179
timestamp 1649977179
transform 1 0 17572 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_184
timestamp 1649977179
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1649977179
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_201
timestamp 1649977179
transform 1 0 19596 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_207
timestamp 1649977179
transform 1 0 20148 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_212
timestamp 1649977179
transform 1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1649977179
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1649977179
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_238
timestamp 1649977179
transform 1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_246
timestamp 1649977179
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_255
timestamp 1649977179
transform 1 0 24564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1649977179
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_269
timestamp 1649977179
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1649977179
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_283
timestamp 1649977179
transform 1 0 27140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_290
timestamp 1649977179
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_297
timestamp 1649977179
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1649977179
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_316
timestamp 1649977179
transform 1 0 30176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_323
timestamp 1649977179
transform 1 0 30820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1649977179
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_340
timestamp 1649977179
transform 1 0 32384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_347
timestamp 1649977179
transform 1 0 33028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_354
timestamp 1649977179
transform 1 0 33672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1649977179
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_368
timestamp 1649977179
transform 1 0 34960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_375
timestamp 1649977179
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_382
timestamp 1649977179
transform 1 0 36248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1649977179
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_396
timestamp 1649977179
transform 1 0 37536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1649977179
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_410
timestamp 1649977179
transform 1 0 38824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1649977179
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_424
timestamp 1649977179
transform 1 0 40112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_431
timestamp 1649977179
transform 1 0 40756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_438
timestamp 1649977179
transform 1 0 41400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1649977179
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_452
timestamp 1649977179
transform 1 0 42688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_459
timestamp 1649977179
transform 1 0 43332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_466
timestamp 1649977179
transform 1 0 43976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1649977179
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_480
timestamp 1649977179
transform 1 0 45264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_487
timestamp 1649977179
transform 1 0 45908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_494
timestamp 1649977179
transform 1 0 46552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1649977179
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_508
timestamp 1649977179
transform 1 0 47840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_515
timestamp 1649977179
transform 1 0 48484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_522
timestamp 1649977179
transform 1 0 49128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_530
timestamp 1649977179
transform 1 0 49864 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_536
timestamp 1649977179
transform 1 0 50416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_543
timestamp 1649977179
transform 1 0 51060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_550
timestamp 1649977179
transform 1 0 51704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_558
timestamp 1649977179
transform 1 0 52440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_564
timestamp 1649977179
transform 1 0 52992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_571
timestamp 1649977179
transform 1 0 53636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_578
timestamp 1649977179
transform 1 0 54280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_586
timestamp 1649977179
transform 1 0 55016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_592
timestamp 1649977179
transform 1 0 55568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_599
timestamp 1649977179
transform 1 0 56212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_606
timestamp 1649977179
transform 1 0 56856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 1649977179
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_620
timestamp 1649977179
transform 1 0 58144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_624
timestamp 1649977179
transform 1 0 58512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_10
timestamp 1649977179
transform 1 0 2024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_30
timestamp 1649977179
transform 1 0 3864 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_38
timestamp 1649977179
transform 1 0 4600 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_43
timestamp 1649977179
transform 1 0 5060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_71
timestamp 1649977179
transform 1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_86
timestamp 1649977179
transform 1 0 9016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1649977179
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106
timestamp 1649977179
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_117
timestamp 1649977179
transform 1 0 11868 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_129
timestamp 1649977179
transform 1 0 12972 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_136
timestamp 1649977179
transform 1 0 13616 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_148
timestamp 1649977179
transform 1 0 14720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_156
timestamp 1649977179
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1649977179
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1649977179
transform 1 0 16928 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1649977179
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1649977179
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_196
timestamp 1649977179
transform 1 0 19136 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_204
timestamp 1649977179
transform 1 0 19872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_212
timestamp 1649977179
transform 1 0 20608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_232
timestamp 1649977179
transform 1 0 22448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_240
timestamp 1649977179
transform 1 0 23184 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_244
timestamp 1649977179
transform 1 0 23552 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_248
timestamp 1649977179
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_255
timestamp 1649977179
transform 1 0 24564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_262
timestamp 1649977179
transform 1 0 25208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_269
timestamp 1649977179
transform 1 0 25852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1649977179
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_285
timestamp 1649977179
transform 1 0 27324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_289
timestamp 1649977179
transform 1 0 27692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_296
timestamp 1649977179
transform 1 0 28336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_303
timestamp 1649977179
transform 1 0 28980 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_310
timestamp 1649977179
transform 1 0 29624 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_317
timestamp 1649977179
transform 1 0 30268 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_324 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 30912 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_340
timestamp 1649977179
transform 1 0 32384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_347
timestamp 1649977179
transform 1 0 33028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_354
timestamp 1649977179
transform 1 0 33672 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_361
timestamp 1649977179
transform 1 0 34316 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_368
timestamp 1649977179
transform 1 0 34960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_375
timestamp 1649977179
transform 1 0 35604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_382
timestamp 1649977179
transform 1 0 36248 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1649977179
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_396
timestamp 1649977179
transform 1 0 37536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1649977179
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_410
timestamp 1649977179
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_417
timestamp 1649977179
transform 1 0 39468 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_424
timestamp 1649977179
transform 1 0 40112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_431
timestamp 1649977179
transform 1 0 40756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_438
timestamp 1649977179
transform 1 0 41400 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1649977179
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_452
timestamp 1649977179
transform 1 0 42688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_459
timestamp 1649977179
transform 1 0 43332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_466
timestamp 1649977179
transform 1 0 43976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_473
timestamp 1649977179
transform 1 0 44620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_480
timestamp 1649977179
transform 1 0 45264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_487
timestamp 1649977179
transform 1 0 45908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_494
timestamp 1649977179
transform 1 0 46552 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1649977179
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_508
timestamp 1649977179
transform 1 0 47840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_515
timestamp 1649977179
transform 1 0 48484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_522
timestamp 1649977179
transform 1 0 49128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_529
timestamp 1649977179
transform 1 0 49772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_536
timestamp 1649977179
transform 1 0 50416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_543
timestamp 1649977179
transform 1 0 51060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_550
timestamp 1649977179
transform 1 0 51704 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_558
timestamp 1649977179
transform 1 0 52440 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_564
timestamp 1649977179
transform 1 0 52992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_571
timestamp 1649977179
transform 1 0 53636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_578
timestamp 1649977179
transform 1 0 54280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_585
timestamp 1649977179
transform 1 0 54924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_592
timestamp 1649977179
transform 1 0 55568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_599
timestamp 1649977179
transform 1 0 56212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_606
timestamp 1649977179
transform 1 0 56856 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_614
timestamp 1649977179
transform 1 0 57592 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_620
timestamp 1649977179
transform 1 0 58144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_624
timestamp 1649977179
transform 1 0 58512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1649977179
transform 1 0 1748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1649977179
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_33
timestamp 1649977179
transform 1 0 4140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_50
timestamp 1649977179
transform 1 0 5704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_58
timestamp 1649977179
transform 1 0 6440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_69
timestamp 1649977179
transform 1 0 7452 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_75
timestamp 1649977179
transform 1 0 8004 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1649977179
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_95
timestamp 1649977179
transform 1 0 9844 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_107
timestamp 1649977179
transform 1 0 10948 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_115
timestamp 1649977179
transform 1 0 11684 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_122
timestamp 1649977179
transform 1 0 12328 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_129
timestamp 1649977179
transform 1 0 12972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1649977179
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_151
timestamp 1649977179
transform 1 0 14996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_158
timestamp 1649977179
transform 1 0 15640 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_178
timestamp 1649977179
transform 1 0 17480 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1649977179
transform 1 0 18032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1649977179
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1649977179
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_210
timestamp 1649977179
transform 1 0 20424 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_214
timestamp 1649977179
transform 1 0 20792 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_219
timestamp 1649977179
transform 1 0 21252 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_223
timestamp 1649977179
transform 1 0 21620 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_228
timestamp 1649977179
transform 1 0 22080 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1649977179
transform 1 0 22632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1649977179
transform 1 0 23276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1649977179
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_257
timestamp 1649977179
transform 1 0 24748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_261
timestamp 1649977179
transform 1 0 25116 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_270
timestamp 1649977179
transform 1 0 25944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_278
timestamp 1649977179
transform 1 0 26680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_282
timestamp 1649977179
transform 1 0 27048 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_291
timestamp 1649977179
transform 1 0 27876 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_299
timestamp 1649977179
transform 1 0 28612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_303
timestamp 1649977179
transform 1 0 28980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_321
timestamp 1649977179
transform 1 0 30636 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_338
timestamp 1649977179
transform 1 0 32200 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_350
timestamp 1649977179
transform 1 0 33304 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp 1649977179
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_369
timestamp 1649977179
transform 1 0 35052 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_376
timestamp 1649977179
transform 1 0 35696 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_383
timestamp 1649977179
transform 1 0 36340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_390
timestamp 1649977179
transform 1 0 36984 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_399
timestamp 1649977179
transform 1 0 37812 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_407
timestamp 1649977179
transform 1 0 38548 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_411
timestamp 1649977179
transform 1 0 38916 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1649977179
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_426
timestamp 1649977179
transform 1 0 40296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_433
timestamp 1649977179
transform 1 0 40940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_440
timestamp 1649977179
transform 1 0 41584 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_448
timestamp 1649977179
transform 1 0 42320 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_453
timestamp 1649977179
transform 1 0 42780 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_460
timestamp 1649977179
transform 1 0 43424 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_472
timestamp 1649977179
transform 1 0 44528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1649977179
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1649977179
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_494
timestamp 1649977179
transform 1 0 46552 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_501
timestamp 1649977179
transform 1 0 47196 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_510
timestamp 1649977179
transform 1 0 48024 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_517
timestamp 1649977179
transform 1 0 48668 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_529
timestamp 1649977179
transform 1 0 49772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_533
timestamp 1649977179
transform 1 0 50140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_537
timestamp 1649977179
transform 1 0 50508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_544
timestamp 1649977179
transform 1 0 51152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_551
timestamp 1649977179
transform 1 0 51796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_558
timestamp 1649977179
transform 1 0 52440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_565
timestamp 1649977179
transform 1 0 53084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_572
timestamp 1649977179
transform 1 0 53728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_579
timestamp 1649977179
transform 1 0 54372 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1649977179
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_592
timestamp 1649977179
transform 1 0 55568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_599
timestamp 1649977179
transform 1 0 56212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_606
timestamp 1649977179
transform 1 0 56856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_610
timestamp 1649977179
transform 1 0 57224 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_614
timestamp 1649977179
transform 1 0 57592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_621
timestamp 1649977179
transform 1 0 58236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_10
timestamp 1649977179
transform 1 0 2024 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_17
timestamp 1649977179
transform 1 0 2668 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_24
timestamp 1649977179
transform 1 0 3312 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_36
timestamp 1649977179
transform 1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_45
timestamp 1649977179
transform 1 0 5244 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1649977179
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1649977179
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_71
timestamp 1649977179
transform 1 0 7636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_86
timestamp 1649977179
transform 1 0 9016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_94
timestamp 1649977179
transform 1 0 9752 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_100
timestamp 1649977179
transform 1 0 10304 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1649977179
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_124
timestamp 1649977179
transform 1 0 12512 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_133
timestamp 1649977179
transform 1 0 13340 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_140
timestamp 1649977179
transform 1 0 13984 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_147
timestamp 1649977179
transform 1 0 14628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_154
timestamp 1649977179
transform 1 0 15272 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp 1649977179
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1649977179
transform 1 0 16928 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_180
timestamp 1649977179
transform 1 0 17664 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_188
timestamp 1649977179
transform 1 0 18400 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_192
timestamp 1649977179
transform 1 0 18768 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_199
timestamp 1649977179
transform 1 0 19412 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_206
timestamp 1649977179
transform 1 0 20056 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_213
timestamp 1649977179
transform 1 0 20700 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1649977179
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_230
timestamp 1649977179
transform 1 0 22264 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_250
timestamp 1649977179
transform 1 0 24104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_257
timestamp 1649977179
transform 1 0 24748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_263
timestamp 1649977179
transform 1 0 25300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_269
timestamp 1649977179
transform 1 0 25852 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_275
timestamp 1649977179
transform 1 0 26404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1649977179
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1649977179
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_369
timestamp 1649977179
transform 1 0 35052 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_386
timestamp 1649977179
transform 1 0 36616 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1649977179
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1649977179
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1649977179
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1649977179
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1649977179
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1649977179
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1649977179
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1649977179
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1649977179
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1649977179
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1649977179
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_541
timestamp 1649977179
transform 1 0 50876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_547
timestamp 1649977179
transform 1 0 51428 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_554
timestamp 1649977179
transform 1 0 52072 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_564
timestamp 1649977179
transform 1 0 52992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_571
timestamp 1649977179
transform 1 0 53636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_578
timestamp 1649977179
transform 1 0 54280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_585
timestamp 1649977179
transform 1 0 54924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_592
timestamp 1649977179
transform 1 0 55568 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_599
timestamp 1649977179
transform 1 0 56212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_611
timestamp 1649977179
transform 1 0 57316 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1649977179
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_617
timestamp 1649977179
transform 1 0 57868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_621
timestamp 1649977179
transform 1 0 58236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1649977179
transform 1 0 1748 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_10
timestamp 1649977179
transform 1 0 2024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_17
timestamp 1649977179
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1649977179
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_33
timestamp 1649977179
transform 1 0 4140 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_49
timestamp 1649977179
transform 1 0 5612 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_61
timestamp 1649977179
transform 1 0 6716 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_67
timestamp 1649977179
transform 1 0 7268 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1649977179
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_89
timestamp 1649977179
transform 1 0 9292 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_102
timestamp 1649977179
transform 1 0 10488 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_117
timestamp 1649977179
transform 1 0 11868 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_125
timestamp 1649977179
transform 1 0 12604 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_129
timestamp 1649977179
transform 1 0 12972 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1649977179
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_146
timestamp 1649977179
transform 1 0 14536 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_160
timestamp 1649977179
transform 1 0 15824 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_167
timestamp 1649977179
transform 1 0 16468 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_174
timestamp 1649977179
transform 1 0 17112 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_185
timestamp 1649977179
transform 1 0 18124 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1649977179
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_216
timestamp 1649977179
transform 1 0 20976 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_225
timestamp 1649977179
transform 1 0 21804 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_232
timestamp 1649977179
transform 1 0 22448 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_239
timestamp 1649977179
transform 1 0 23092 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_246
timestamp 1649977179
transform 1 0 23736 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_269
timestamp 1649977179
transform 1 0 25852 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_281
timestamp 1649977179
transform 1 0 26956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_299
timestamp 1649977179
transform 1 0 28612 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_343
timestamp 1649977179
transform 1 0 32660 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_355
timestamp 1649977179
transform 1 0 33764 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1649977179
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1649977179
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1649977179
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1649977179
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1649977179
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1649977179
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1649977179
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1649977179
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1649977179
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1649977179
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_545
timestamp 1649977179
transform 1 0 51244 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_553
timestamp 1649977179
transform 1 0 51980 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_558
timestamp 1649977179
transform 1 0 52440 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_565
timestamp 1649977179
transform 1 0 53084 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_572
timestamp 1649977179
transform 1 0 53728 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_579
timestamp 1649977179
transform 1 0 54372 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1649977179
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_592
timestamp 1649977179
transform 1 0 55568 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_599
timestamp 1649977179
transform 1 0 56212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_611
timestamp 1649977179
transform 1 0 57316 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_623
timestamp 1649977179
transform 1 0 58420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_8
timestamp 1649977179
transform 1 0 1840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_28
timestamp 1649977179
transform 1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_32
timestamp 1649977179
transform 1 0 4048 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_36
timestamp 1649977179
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_44
timestamp 1649977179
transform 1 0 5152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1649977179
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_67
timestamp 1649977179
transform 1 0 7268 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_79
timestamp 1649977179
transform 1 0 8372 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_90
timestamp 1649977179
transform 1 0 9384 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_101
timestamp 1649977179
transform 1 0 10396 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_123
timestamp 1649977179
transform 1 0 12420 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_131
timestamp 1649977179
transform 1 0 13156 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_135
timestamp 1649977179
transform 1 0 13524 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_142
timestamp 1649977179
transform 1 0 14168 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_154
timestamp 1649977179
transform 1 0 15272 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_175
timestamp 1649977179
transform 1 0 17204 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_182
timestamp 1649977179
transform 1 0 17848 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_194
timestamp 1649977179
transform 1 0 18952 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_201
timestamp 1649977179
transform 1 0 19596 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_210
timestamp 1649977179
transform 1 0 20424 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_219
timestamp 1649977179
transform 1 0 21252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_227
timestamp 1649977179
transform 1 0 21988 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_234
timestamp 1649977179
transform 1 0 22632 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_240
timestamp 1649977179
transform 1 0 23184 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_246
timestamp 1649977179
transform 1 0 23736 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_252
timestamp 1649977179
transform 1 0 24288 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_258
timestamp 1649977179
transform 1 0 24840 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_270
timestamp 1649977179
transform 1 0 25944 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1649977179
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_292
timestamp 1649977179
transform 1 0 27968 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_304
timestamp 1649977179
transform 1 0 29072 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_312
timestamp 1649977179
transform 1 0 29808 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_324
timestamp 1649977179
transform 1 0 30912 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1649977179
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_410
timestamp 1649977179
transform 1 0 38824 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_422
timestamp 1649977179
transform 1 0 39928 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_434
timestamp 1649977179
transform 1 0 41032 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_446
timestamp 1649977179
transform 1 0 42136 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1649977179
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1649977179
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1649977179
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1649977179
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1649977179
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1649977179
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1649977179
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1649977179
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1649977179
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_561
timestamp 1649977179
transform 1 0 52716 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_569
timestamp 1649977179
transform 1 0 53452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_575
timestamp 1649977179
transform 1 0 54004 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_582
timestamp 1649977179
transform 1 0 54648 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_589
timestamp 1649977179
transform 1 0 55292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_601
timestamp 1649977179
transform 1 0 56396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_613
timestamp 1649977179
transform 1 0 57500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_617
timestamp 1649977179
transform 1 0 57868 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_621
timestamp 1649977179
transform 1 0 58236 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_8
timestamp 1649977179
transform 1 0 1840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_21
timestamp 1649977179
transform 1 0 3036 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1649977179
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_66
timestamp 1649977179
transform 1 0 7176 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_74
timestamp 1649977179
transform 1 0 7912 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1649977179
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1649977179
transform 1 0 9200 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_95
timestamp 1649977179
transform 1 0 9844 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_102
timestamp 1649977179
transform 1 0 10488 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_116
timestamp 1649977179
transform 1 0 11776 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_123
timestamp 1649977179
transform 1 0 12420 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_130
timestamp 1649977179
transform 1 0 13064 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1649977179
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_159
timestamp 1649977179
transform 1 0 15732 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_171
timestamp 1649977179
transform 1 0 16836 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_179
timestamp 1649977179
transform 1 0 17572 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_191
timestamp 1649977179
transform 1 0 18676 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_213
timestamp 1649977179
transform 1 0 20700 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1649977179
transform 1 0 21252 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_222
timestamp 1649977179
transform 1 0 21528 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_228
timestamp 1649977179
transform 1 0 22080 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_232
timestamp 1649977179
transform 1 0 22448 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_240
timestamp 1649977179
transform 1 0 23184 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_246
timestamp 1649977179
transform 1 0 23736 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_255
timestamp 1649977179
transform 1 0 24564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_264
timestamp 1649977179
transform 1 0 25392 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_270
timestamp 1649977179
transform 1 0 25944 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_273
timestamp 1649977179
transform 1 0 26220 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_281
timestamp 1649977179
transform 1 0 26956 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_297
timestamp 1649977179
transform 1 0 28428 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_305
timestamp 1649977179
transform 1 0 29164 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_313
timestamp 1649977179
transform 1 0 29900 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_325
timestamp 1649977179
transform 1 0 31004 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_334
timestamp 1649977179
transform 1 0 31832 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_343
timestamp 1649977179
transform 1 0 32660 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_355
timestamp 1649977179
transform 1 0 33764 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_381
timestamp 1649977179
transform 1 0 36156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_387
timestamp 1649977179
transform 1 0 36708 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_411
timestamp 1649977179
transform 1 0 38916 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1649977179
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1649977179
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1649977179
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1649977179
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1649977179
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1649977179
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1649977179
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1649977179
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1649977179
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1649977179
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1649977179
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1649977179
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1649977179
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1649977179
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1649977179
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1649977179
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1649977179
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_9
timestamp 1649977179
transform 1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_29
timestamp 1649977179
transform 1 0 3772 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_37
timestamp 1649977179
transform 1 0 4508 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_44
timestamp 1649977179
transform 1 0 5152 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_48
timestamp 1649977179
transform 1 0 5520 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1649977179
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_64
timestamp 1649977179
transform 1 0 6992 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_70
timestamp 1649977179
transform 1 0 7544 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_74
timestamp 1649977179
transform 1 0 7912 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_101
timestamp 1649977179
transform 1 0 10396 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1649977179
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_117
timestamp 1649977179
transform 1 0 11868 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_124
timestamp 1649977179
transform 1 0 12512 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_133
timestamp 1649977179
transform 1 0 13340 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_140
timestamp 1649977179
transform 1 0 13984 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1649977179
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_179
timestamp 1649977179
transform 1 0 17572 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_187
timestamp 1649977179
transform 1 0 18308 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_202
timestamp 1649977179
transform 1 0 19688 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_208
timestamp 1649977179
transform 1 0 20240 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_214
timestamp 1649977179
transform 1 0 20792 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1649977179
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_235
timestamp 1649977179
transform 1 0 22724 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_246
timestamp 1649977179
transform 1 0 23736 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_250
timestamp 1649977179
transform 1 0 24104 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_271
timestamp 1649977179
transform 1 0 26036 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_291
timestamp 1649977179
transform 1 0 27876 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_300
timestamp 1649977179
transform 1 0 28704 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_308
timestamp 1649977179
transform 1 0 29440 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_312
timestamp 1649977179
transform 1 0 29808 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_324
timestamp 1649977179
transform 1 0 30912 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_339
timestamp 1649977179
transform 1 0 32292 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_351
timestamp 1649977179
transform 1 0 33396 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_357
timestamp 1649977179
transform 1 0 33948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_363
timestamp 1649977179
transform 1 0 34500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_375
timestamp 1649977179
transform 1 0 35604 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_384
timestamp 1649977179
transform 1 0 36432 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_398
timestamp 1649977179
transform 1 0 37720 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_420
timestamp 1649977179
transform 1 0 39744 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_432
timestamp 1649977179
transform 1 0 40848 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_444
timestamp 1649977179
transform 1 0 41952 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1649977179
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1649977179
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1649977179
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1649977179
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1649977179
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1649977179
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1649977179
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1649977179
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1649977179
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1649977179
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1649977179
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1649977179
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_617
timestamp 1649977179
transform 1 0 57868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_621
timestamp 1649977179
transform 1 0 58236 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_7
timestamp 1649977179
transform 1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_16
timestamp 1649977179
transform 1 0 2576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1649977179
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_31
timestamp 1649977179
transform 1 0 3956 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_37
timestamp 1649977179
transform 1 0 4508 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_43
timestamp 1649977179
transform 1 0 5060 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_49
timestamp 1649977179
transform 1 0 5612 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_56
timestamp 1649977179
transform 1 0 6256 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_63
timestamp 1649977179
transform 1 0 6900 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_70
timestamp 1649977179
transform 1 0 7544 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_88
timestamp 1649977179
transform 1 0 9200 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_98
timestamp 1649977179
transform 1 0 10120 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_118
timestamp 1649977179
transform 1 0 11960 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_122
timestamp 1649977179
transform 1 0 12328 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_126
timestamp 1649977179
transform 1 0 12696 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_145
timestamp 1649977179
transform 1 0 14444 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_151
timestamp 1649977179
transform 1 0 14996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_162
timestamp 1649977179
transform 1 0 16008 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_166
timestamp 1649977179
transform 1 0 16376 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_169
timestamp 1649977179
transform 1 0 16652 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_175
timestamp 1649977179
transform 1 0 17204 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_178
timestamp 1649977179
transform 1 0 17480 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1649977179
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_199
timestamp 1649977179
transform 1 0 19412 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_203
timestamp 1649977179
transform 1 0 19780 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_206
timestamp 1649977179
transform 1 0 20056 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_212
timestamp 1649977179
transform 1 0 20608 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_218
timestamp 1649977179
transform 1 0 21160 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_224
timestamp 1649977179
transform 1 0 21712 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_235
timestamp 1649977179
transform 1 0 22724 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_239
timestamp 1649977179
transform 1 0 23092 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1649977179
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_261
timestamp 1649977179
transform 1 0 25116 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_269
timestamp 1649977179
transform 1 0 25852 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_280
timestamp 1649977179
transform 1 0 26864 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_300
timestamp 1649977179
transform 1 0 28704 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_313
timestamp 1649977179
transform 1 0 29900 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_334
timestamp 1649977179
transform 1 0 31832 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_356
timestamp 1649977179
transform 1 0 33856 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_385
timestamp 1649977179
transform 1 0 36524 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_394
timestamp 1649977179
transform 1 0 37352 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_400
timestamp 1649977179
transform 1 0 37904 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_404
timestamp 1649977179
transform 1 0 38272 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1649977179
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1649977179
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_423
timestamp 1649977179
transform 1 0 40020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_435
timestamp 1649977179
transform 1 0 41124 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_447
timestamp 1649977179
transform 1 0 42228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_459
timestamp 1649977179
transform 1 0 43332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_471
timestamp 1649977179
transform 1 0 44436 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1649977179
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1649977179
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1649977179
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1649977179
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1649977179
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1649977179
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1649977179
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1649977179
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1649977179
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1649977179
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1649977179
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1649977179
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1649977179
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1649977179
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_8
timestamp 1649977179
transform 1 0 1840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_17
timestamp 1649977179
transform 1 0 2668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_30
timestamp 1649977179
transform 1 0 3864 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_36
timestamp 1649977179
transform 1 0 4416 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_45
timestamp 1649977179
transform 1 0 5244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_49
timestamp 1649977179
transform 1 0 5612 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_65
timestamp 1649977179
transform 1 0 7084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_78
timestamp 1649977179
transform 1 0 8280 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_84
timestamp 1649977179
transform 1 0 8832 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_90
timestamp 1649977179
transform 1 0 9384 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_96
timestamp 1649977179
transform 1 0 9936 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_102
timestamp 1649977179
transform 1 0 10488 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_130
timestamp 1649977179
transform 1 0 13064 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_136
timestamp 1649977179
transform 1 0 13616 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_139
timestamp 1649977179
transform 1 0 13892 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_147
timestamp 1649977179
transform 1 0 14628 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_159
timestamp 1649977179
transform 1 0 15732 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_174
timestamp 1649977179
transform 1 0 17112 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_180
timestamp 1649977179
transform 1 0 17664 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_186
timestamp 1649977179
transform 1 0 18216 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_190
timestamp 1649977179
transform 1 0 18584 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_194
timestamp 1649977179
transform 1 0 18952 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_200
timestamp 1649977179
transform 1 0 19504 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_208
timestamp 1649977179
transform 1 0 20240 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_211
timestamp 1649977179
transform 1 0 20516 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1649977179
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_229
timestamp 1649977179
transform 1 0 22172 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_246
timestamp 1649977179
transform 1 0 23736 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_252
timestamp 1649977179
transform 1 0 24288 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_264
timestamp 1649977179
transform 1 0 25392 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_300
timestamp 1649977179
transform 1 0 28704 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_312
timestamp 1649977179
transform 1 0 29808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_332
timestamp 1649977179
transform 1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_357
timestamp 1649977179
transform 1 0 33948 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_365
timestamp 1649977179
transform 1 0 34684 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_376
timestamp 1649977179
transform 1 0 35696 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_384
timestamp 1649977179
transform 1 0 36432 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_403
timestamp 1649977179
transform 1 0 38180 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_412
timestamp 1649977179
transform 1 0 39008 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_424
timestamp 1649977179
transform 1 0 40112 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_436
timestamp 1649977179
transform 1 0 41216 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1649977179
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1649977179
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1649977179
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1649977179
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1649977179
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1649977179
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1649977179
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1649977179
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1649977179
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1649977179
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1649977179
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1649977179
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1649977179
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_617
timestamp 1649977179
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_5
timestamp 1649977179
transform 1 0 1564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_11
timestamp 1649977179
transform 1 0 2116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1649977179
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_32
timestamp 1649977179
transform 1 0 4048 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_38
timestamp 1649977179
transform 1 0 4600 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_48
timestamp 1649977179
transform 1 0 5520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_68
timestamp 1649977179
transform 1 0 7360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_94
timestamp 1649977179
transform 1 0 9752 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_106
timestamp 1649977179
transform 1 0 10856 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_112
timestamp 1649977179
transform 1 0 11408 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_118
timestamp 1649977179
transform 1 0 11960 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_124
timestamp 1649977179
transform 1 0 12512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_130
timestamp 1649977179
transform 1 0 13064 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_145
timestamp 1649977179
transform 1 0 14444 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_159
timestamp 1649977179
transform 1 0 15732 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_167
timestamp 1649977179
transform 1 0 16468 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_170
timestamp 1649977179
transform 1 0 16744 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_176
timestamp 1649977179
transform 1 0 17296 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_188
timestamp 1649977179
transform 1 0 18400 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_201
timestamp 1649977179
transform 1 0 19596 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_214
timestamp 1649977179
transform 1 0 20792 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_225
timestamp 1649977179
transform 1 0 21804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_242
timestamp 1649977179
transform 1 0 23368 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1649977179
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_257
timestamp 1649977179
transform 1 0 24748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_274
timestamp 1649977179
transform 1 0 26312 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_282
timestamp 1649977179
transform 1 0 27048 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_293
timestamp 1649977179
transform 1 0 28060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_305
timestamp 1649977179
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_326
timestamp 1649977179
transform 1 0 31096 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_338
timestamp 1649977179
transform 1 0 32200 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_350
timestamp 1649977179
transform 1 0 33304 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 1649977179
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_376
timestamp 1649977179
transform 1 0 35696 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_388
timestamp 1649977179
transform 1 0 36800 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_400
timestamp 1649977179
transform 1 0 37904 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_412
timestamp 1649977179
transform 1 0 39008 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1649977179
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1649977179
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1649977179
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1649977179
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1649977179
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1649977179
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1649977179
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1649977179
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1649977179
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1649977179
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1649977179
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1649977179
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1649977179
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1649977179
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1649977179
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1649977179
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1649977179
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1649977179
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_613
timestamp 1649977179
transform 1 0 57500 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_617
timestamp 1649977179
transform 1 0 57868 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_621
timestamp 1649977179
transform 1 0 58236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_7
timestamp 1649977179
transform 1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_13
timestamp 1649977179
transform 1 0 2300 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_19
timestamp 1649977179
transform 1 0 2852 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_23
timestamp 1649977179
transform 1 0 3220 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_26
timestamp 1649977179
transform 1 0 3496 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_32
timestamp 1649977179
transform 1 0 4048 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_35
timestamp 1649977179
transform 1 0 4324 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_41
timestamp 1649977179
transform 1 0 4876 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1649977179
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_67
timestamp 1649977179
transform 1 0 7268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_73
timestamp 1649977179
transform 1 0 7820 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_88
timestamp 1649977179
transform 1 0 9200 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_94
timestamp 1649977179
transform 1 0 9752 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_100
timestamp 1649977179
transform 1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_106
timestamp 1649977179
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_122
timestamp 1649977179
transform 1 0 12328 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_128
timestamp 1649977179
transform 1 0 12880 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_136
timestamp 1649977179
transform 1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_144
timestamp 1649977179
transform 1 0 14352 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1649977179
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_174
timestamp 1649977179
transform 1 0 17112 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_180
timestamp 1649977179
transform 1 0 17664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_192
timestamp 1649977179
transform 1 0 18768 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_201
timestamp 1649977179
transform 1 0 19596 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_210
timestamp 1649977179
transform 1 0 20424 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_214
timestamp 1649977179
transform 1 0 20792 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_235
timestamp 1649977179
transform 1 0 22724 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_241
timestamp 1649977179
transform 1 0 23276 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_250
timestamp 1649977179
transform 1 0 24104 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_262
timestamp 1649977179
transform 1 0 25208 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_274
timestamp 1649977179
transform 1 0 26312 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_289
timestamp 1649977179
transform 1 0 27692 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_302
timestamp 1649977179
transform 1 0 28888 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_313
timestamp 1649977179
transform 1 0 29900 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_325
timestamp 1649977179
transform 1 0 31004 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp 1649977179
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_344
timestamp 1649977179
transform 1 0 32752 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_356
timestamp 1649977179
transform 1 0 33856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_364
timestamp 1649977179
transform 1 0 34592 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_376
timestamp 1649977179
transform 1 0 35696 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_384
timestamp 1649977179
transform 1 0 36432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_388
timestamp 1649977179
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_398
timestamp 1649977179
transform 1 0 37720 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_410
timestamp 1649977179
transform 1 0 38824 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_422
timestamp 1649977179
transform 1 0 39928 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_434
timestamp 1649977179
transform 1 0 41032 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_446
timestamp 1649977179
transform 1 0 42136 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1649977179
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1649977179
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1649977179
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1649977179
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1649977179
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1649977179
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1649977179
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1649977179
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1649977179
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1649977179
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1649977179
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1649977179
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1649977179
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1649977179
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1649977179
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1649977179
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_21
timestamp 1649977179
transform 1 0 3036 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1649977179
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_34
timestamp 1649977179
transform 1 0 4232 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_46
timestamp 1649977179
transform 1 0 5336 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_52
timestamp 1649977179
transform 1 0 5888 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_56
timestamp 1649977179
transform 1 0 6256 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_61
timestamp 1649977179
transform 1 0 6716 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_67
timestamp 1649977179
transform 1 0 7268 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_73
timestamp 1649977179
transform 1 0 7820 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1649977179
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1649977179
transform 1 0 9660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_99
timestamp 1649977179
transform 1 0 10212 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_107
timestamp 1649977179
transform 1 0 10948 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_119
timestamp 1649977179
transform 1 0 12052 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_127
timestamp 1649977179
transform 1 0 12788 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_157
timestamp 1649977179
transform 1 0 15548 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_163
timestamp 1649977179
transform 1 0 16100 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_166
timestamp 1649977179
transform 1 0 16376 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_172
timestamp 1649977179
transform 1 0 16928 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1649977179
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_213
timestamp 1649977179
transform 1 0 20700 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_220
timestamp 1649977179
transform 1 0 21344 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_226
timestamp 1649977179
transform 1 0 21896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_237
timestamp 1649977179
transform 1 0 22908 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_243
timestamp 1649977179
transform 1 0 23460 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_293
timestamp 1649977179
transform 1 0 28060 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1649977179
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_328
timestamp 1649977179
transform 1 0 31280 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_339
timestamp 1649977179
transform 1 0 32292 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_350
timestamp 1649977179
transform 1 0 33304 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 1649977179
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_381
timestamp 1649977179
transform 1 0 36156 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_387
timestamp 1649977179
transform 1 0 36708 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_396
timestamp 1649977179
transform 1 0 37536 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_416
timestamp 1649977179
transform 1 0 39376 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1649977179
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1649977179
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1649977179
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1649977179
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1649977179
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1649977179
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1649977179
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1649977179
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1649977179
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1649977179
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1649977179
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1649977179
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1649977179
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1649977179
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1649977179
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1649977179
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_613
timestamp 1649977179
transform 1 0 57500 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_617
timestamp 1649977179
transform 1 0 57868 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_621
timestamp 1649977179
transform 1 0 58236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_9
timestamp 1649977179
transform 1 0 1932 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_26
timestamp 1649977179
transform 1 0 3496 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_38
timestamp 1649977179
transform 1 0 4600 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1649977179
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_59
timestamp 1649977179
transform 1 0 6532 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_71
timestamp 1649977179
transform 1 0 7636 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_83
timestamp 1649977179
transform 1 0 8740 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_95
timestamp 1649977179
transform 1 0 9844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1649977179
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_121
timestamp 1649977179
transform 1 0 12236 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_130
timestamp 1649977179
transform 1 0 13064 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_142
timestamp 1649977179
transform 1 0 14168 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_146
timestamp 1649977179
transform 1 0 14536 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_154
timestamp 1649977179
transform 1 0 15272 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp 1649977179
transform 1 0 15824 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_172
timestamp 1649977179
transform 1 0 16928 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_196
timestamp 1649977179
transform 1 0 19136 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_208
timestamp 1649977179
transform 1 0 20240 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_212
timestamp 1649977179
transform 1 0 20608 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_215
timestamp 1649977179
transform 1 0 20884 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_238
timestamp 1649977179
transform 1 0 23000 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_250
timestamp 1649977179
transform 1 0 24104 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_257
timestamp 1649977179
transform 1 0 24748 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_266
timestamp 1649977179
transform 1 0 25576 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1649977179
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_311
timestamp 1649977179
transform 1 0 29716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_315
timestamp 1649977179
transform 1 0 30084 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1649977179
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_345
timestamp 1649977179
transform 1 0 32844 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_351
timestamp 1649977179
transform 1 0 33396 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_363
timestamp 1649977179
transform 1 0 34500 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_376
timestamp 1649977179
transform 1 0 35696 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_388
timestamp 1649977179
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_400
timestamp 1649977179
transform 1 0 37904 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_420
timestamp 1649977179
transform 1 0 39744 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_432
timestamp 1649977179
transform 1 0 40848 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_444
timestamp 1649977179
transform 1 0 41952 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1649977179
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1649977179
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1649977179
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1649977179
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1649977179
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1649977179
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1649977179
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1649977179
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1649977179
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1649977179
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1649977179
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1649977179
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1649977179
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1649977179
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1649977179
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1649977179
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1649977179
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_11
timestamp 1649977179
transform 1 0 2116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1649977179
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_31
timestamp 1649977179
transform 1 0 3956 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_39
timestamp 1649977179
transform 1 0 4692 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_45
timestamp 1649977179
transform 1 0 5244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_57
timestamp 1649977179
transform 1 0 6348 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_61
timestamp 1649977179
transform 1 0 6716 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_66
timestamp 1649977179
transform 1 0 7176 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_78
timestamp 1649977179
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_94
timestamp 1649977179
transform 1 0 9752 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_100
timestamp 1649977179
transform 1 0 10304 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_134
timestamp 1649977179
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_217
timestamp 1649977179
transform 1 0 21068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_230
timestamp 1649977179
transform 1 0 22264 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_242
timestamp 1649977179
transform 1 0 23368 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1649977179
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_276
timestamp 1649977179
transform 1 0 26496 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_284
timestamp 1649977179
transform 1 0 27232 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_293
timestamp 1649977179
transform 1 0 28060 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1649977179
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_314
timestamp 1649977179
transform 1 0 29992 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_320
timestamp 1649977179
transform 1 0 30544 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_323
timestamp 1649977179
transform 1 0 30820 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_347
timestamp 1649977179
transform 1 0 33028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_359
timestamp 1649977179
transform 1 0 34132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_385
timestamp 1649977179
transform 1 0 36524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_390
timestamp 1649977179
transform 1 0 36984 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_396
timestamp 1649977179
transform 1 0 37536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_408
timestamp 1649977179
transform 1 0 38640 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_414
timestamp 1649977179
transform 1 0 39192 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1649977179
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1649977179
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1649977179
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1649977179
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1649977179
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1649977179
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1649977179
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1649977179
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1649977179
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1649977179
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1649977179
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1649977179
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1649977179
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1649977179
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1649977179
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1649977179
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1649977179
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1649977179
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1649977179
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_11
timestamp 1649977179
transform 1 0 2116 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_33
timestamp 1649977179
transform 1 0 4140 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_38
timestamp 1649977179
transform 1 0 4600 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_50
timestamp 1649977179
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_65
timestamp 1649977179
transform 1 0 7084 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_74
timestamp 1649977179
transform 1 0 7912 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_94
timestamp 1649977179
transform 1 0 9752 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_100
timestamp 1649977179
transform 1 0 10304 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_121
timestamp 1649977179
transform 1 0 12236 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_131
timestamp 1649977179
transform 1 0 13156 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_139
timestamp 1649977179
transform 1 0 13892 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_156
timestamp 1649977179
transform 1 0 15456 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1649977179
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_202
timestamp 1649977179
transform 1 0 19688 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_214
timestamp 1649977179
transform 1 0 20792 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1649977179
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_236
timestamp 1649977179
transform 1 0 22816 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_244
timestamp 1649977179
transform 1 0 23552 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_256
timestamp 1649977179
transform 1 0 24656 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1649977179
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_296
timestamp 1649977179
transform 1 0 28336 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_308
timestamp 1649977179
transform 1 0 29440 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_314
timestamp 1649977179
transform 1 0 29992 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_320
timestamp 1649977179
transform 1 0 30544 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_326
timestamp 1649977179
transform 1 0 31096 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1649977179
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_361
timestamp 1649977179
transform 1 0 34316 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1649977179
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_417
timestamp 1649977179
transform 1 0 39468 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_437
timestamp 1649977179
transform 1 0 41308 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_445
timestamp 1649977179
transform 1 0 42044 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1649977179
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1649977179
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1649977179
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1649977179
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1649977179
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1649977179
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1649977179
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1649977179
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1649977179
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1649977179
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1649977179
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1649977179
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1649977179
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1649977179
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1649977179
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1649977179
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_617
timestamp 1649977179
transform 1 0 57868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_621
timestamp 1649977179
transform 1 0 58236 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_11
timestamp 1649977179
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1649977179
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_32
timestamp 1649977179
transform 1 0 4048 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_44
timestamp 1649977179
transform 1 0 5152 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_66
timestamp 1649977179
transform 1 0 7176 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1649977179
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_88
timestamp 1649977179
transform 1 0 9200 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_100
timestamp 1649977179
transform 1 0 10304 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_112
timestamp 1649977179
transform 1 0 11408 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_117
timestamp 1649977179
transform 1 0 11868 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_125
timestamp 1649977179
transform 1 0 12604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1649977179
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_158
timestamp 1649977179
transform 1 0 15640 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1649977179
transform 1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_174
timestamp 1649977179
transform 1 0 17112 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_180
timestamp 1649977179
transform 1 0 17664 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_183
timestamp 1649977179
transform 1 0 17940 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1649977179
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_203
timestamp 1649977179
transform 1 0 19780 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_211
timestamp 1649977179
transform 1 0 20516 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1649977179
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_239
timestamp 1649977179
transform 1 0 23092 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_246
timestamp 1649977179
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_273
timestamp 1649977179
transform 1 0 26220 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_285
timestamp 1649977179
transform 1 0 27324 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_293
timestamp 1649977179
transform 1 0 28060 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1649977179
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_314
timestamp 1649977179
transform 1 0 29992 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_326
timestamp 1649977179
transform 1 0 31096 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_340
timestamp 1649977179
transform 1 0 32384 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_344
timestamp 1649977179
transform 1 0 32752 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_347
timestamp 1649977179
transform 1 0 33028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_359
timestamp 1649977179
transform 1 0 34132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1649977179
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_367
timestamp 1649977179
transform 1 0 34868 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_379
timestamp 1649977179
transform 1 0 35972 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_388
timestamp 1649977179
transform 1 0 36800 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_396
timestamp 1649977179
transform 1 0 37536 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_404
timestamp 1649977179
transform 1 0 38272 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_416
timestamp 1649977179
transform 1 0 39376 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_423
timestamp 1649977179
transform 1 0 40020 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_435
timestamp 1649977179
transform 1 0 41124 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_447
timestamp 1649977179
transform 1 0 42228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_459
timestamp 1649977179
transform 1 0 43332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_471
timestamp 1649977179
transform 1 0 44436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1649977179
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1649977179
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1649977179
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1649977179
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1649977179
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1649977179
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1649977179
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1649977179
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1649977179
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1649977179
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1649977179
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1649977179
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1649977179
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1649977179
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1649977179
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_35
timestamp 1649977179
transform 1 0 4324 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_44
timestamp 1649977179
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_67
timestamp 1649977179
transform 1 0 7268 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_87
timestamp 1649977179
transform 1 0 9108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_99
timestamp 1649977179
transform 1 0 10212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_123
timestamp 1649977179
transform 1 0 12420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_135
timestamp 1649977179
transform 1 0 13524 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_141
timestamp 1649977179
transform 1 0 14076 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1649977179
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_159
timestamp 1649977179
transform 1 0 15732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_177
timestamp 1649977179
transform 1 0 17388 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_180
timestamp 1649977179
transform 1 0 17664 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_192
timestamp 1649977179
transform 1 0 18768 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_200
timestamp 1649977179
transform 1 0 19504 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1649977179
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_243
timestamp 1649977179
transform 1 0 23460 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_255
timestamp 1649977179
transform 1 0 24564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_259
timestamp 1649977179
transform 1 0 24932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_262
timestamp 1649977179
transform 1 0 25208 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_274
timestamp 1649977179
transform 1 0 26312 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_298
timestamp 1649977179
transform 1 0 28520 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_310
timestamp 1649977179
transform 1 0 29624 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_322
timestamp 1649977179
transform 1 0 30728 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1649977179
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_342
timestamp 1649977179
transform 1 0 32568 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_346
timestamp 1649977179
transform 1 0 32936 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_357
timestamp 1649977179
transform 1 0 33948 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_363
timestamp 1649977179
transform 1 0 34500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_366
timestamp 1649977179
transform 1 0 34776 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_377
timestamp 1649977179
transform 1 0 35788 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_401
timestamp 1649977179
transform 1 0 37996 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_405
timestamp 1649977179
transform 1 0 38364 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_419
timestamp 1649977179
transform 1 0 39652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_431
timestamp 1649977179
transform 1 0 40756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_443
timestamp 1649977179
transform 1 0 41860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1649977179
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1649977179
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1649977179
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1649977179
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1649977179
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1649977179
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1649977179
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1649977179
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1649977179
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1649977179
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1649977179
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1649977179
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1649977179
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1649977179
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1649977179
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_617
timestamp 1649977179
transform 1 0 57868 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_621
timestamp 1649977179
transform 1 0 58236 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_18
timestamp 1649977179
transform 1 0 2760 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1649977179
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_33
timestamp 1649977179
transform 1 0 4140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_36
timestamp 1649977179
transform 1 0 4416 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_49
timestamp 1649977179
transform 1 0 5612 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_57
timestamp 1649977179
transform 1 0 6348 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1649977179
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_87
timestamp 1649977179
transform 1 0 9108 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_99
timestamp 1649977179
transform 1 0 10212 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_129
timestamp 1649977179
transform 1 0 12972 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_152
timestamp 1649977179
transform 1 0 15088 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_158
timestamp 1649977179
transform 1 0 15640 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_170
timestamp 1649977179
transform 1 0 16744 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_202
timestamp 1649977179
transform 1 0 19688 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_218
timestamp 1649977179
transform 1 0 21160 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_230
timestamp 1649977179
transform 1 0 22264 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_236
timestamp 1649977179
transform 1 0 22816 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_246
timestamp 1649977179
transform 1 0 23736 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_255
timestamp 1649977179
transform 1 0 24564 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_261
timestamp 1649977179
transform 1 0 25116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_281
timestamp 1649977179
transform 1 0 26956 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_285
timestamp 1649977179
transform 1 0 27324 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_290
timestamp 1649977179
transform 1 0 27784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_298
timestamp 1649977179
transform 1 0 28520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1649977179
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_324
timestamp 1649977179
transform 1 0 30912 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_336
timestamp 1649977179
transform 1 0 32016 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_356
timestamp 1649977179
transform 1 0 33856 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_375
timestamp 1649977179
transform 1 0 35604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_387
timestamp 1649977179
transform 1 0 36708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_393
timestamp 1649977179
transform 1 0 37260 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_404
timestamp 1649977179
transform 1 0 38272 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_416
timestamp 1649977179
transform 1 0 39376 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1649977179
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1649977179
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1649977179
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1649977179
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1649977179
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1649977179
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1649977179
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1649977179
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1649977179
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1649977179
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1649977179
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1649977179
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1649977179
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1649977179
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1649977179
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1649977179
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1649977179
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1649977179
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1649977179
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_14
timestamp 1649977179
transform 1 0 2392 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_34
timestamp 1649977179
transform 1 0 4232 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1649977179
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_83
timestamp 1649977179
transform 1 0 8740 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_95
timestamp 1649977179
transform 1 0 9844 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_115
timestamp 1649977179
transform 1 0 11684 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_127
timestamp 1649977179
transform 1 0 12788 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_139
timestamp 1649977179
transform 1 0 13892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_150
timestamp 1649977179
transform 1 0 14904 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_156
timestamp 1649977179
transform 1 0 15456 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_189
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_201
timestamp 1649977179
transform 1 0 19596 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_210
timestamp 1649977179
transform 1 0 20424 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_219
timestamp 1649977179
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_229
timestamp 1649977179
transform 1 0 22172 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_251
timestamp 1649977179
transform 1 0 24196 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_259
timestamp 1649977179
transform 1 0 24932 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_265
timestamp 1649977179
transform 1 0 25484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1649977179
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_283
timestamp 1649977179
transform 1 0 27140 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_291
timestamp 1649977179
transform 1 0 27876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_303
timestamp 1649977179
transform 1 0 28980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_309
timestamp 1649977179
transform 1 0 29532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_312
timestamp 1649977179
transform 1 0 29808 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_320
timestamp 1649977179
transform 1 0 30544 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_328
timestamp 1649977179
transform 1 0 31280 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_332
timestamp 1649977179
transform 1 0 31648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_347
timestamp 1649977179
transform 1 0 33028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_359
timestamp 1649977179
transform 1 0 34132 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_369
timestamp 1649977179
transform 1 0 35052 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_383
timestamp 1649977179
transform 1 0 36340 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1649977179
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1649977179
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_423
timestamp 1649977179
transform 1 0 40020 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_435
timestamp 1649977179
transform 1 0 41124 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1649977179
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1649977179
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1649977179
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1649977179
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1649977179
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1649977179
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1649977179
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1649977179
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1649977179
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1649977179
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1649977179
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1649977179
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1649977179
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1649977179
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1649977179
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1649977179
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1649977179
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1649977179
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1649977179
transform 1 0 2116 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_16
timestamp 1649977179
transform 1 0 2576 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_35
timestamp 1649977179
transform 1 0 4324 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_38
timestamp 1649977179
transform 1 0 4600 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_50
timestamp 1649977179
transform 1 0 5704 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_56
timestamp 1649977179
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_71
timestamp 1649977179
transform 1 0 7636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_103
timestamp 1649977179
transform 1 0 10580 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_115
timestamp 1649977179
transform 1 0 11684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_127
timestamp 1649977179
transform 1 0 12788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_146
timestamp 1649977179
transform 1 0 14536 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_158
timestamp 1649977179
transform 1 0 15640 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_170
timestamp 1649977179
transform 1 0 16744 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_178
timestamp 1649977179
transform 1 0 17480 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_185
timestamp 1649977179
transform 1 0 18124 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1649977179
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_201
timestamp 1649977179
transform 1 0 19596 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_206
timestamp 1649977179
transform 1 0 20056 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_212
timestamp 1649977179
transform 1 0 20608 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_222
timestamp 1649977179
transform 1 0 21528 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_234
timestamp 1649977179
transform 1 0 22632 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_244
timestamp 1649977179
transform 1 0 23552 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_260
timestamp 1649977179
transform 1 0 25024 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_268
timestamp 1649977179
transform 1 0 25760 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_271
timestamp 1649977179
transform 1 0 26036 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_295
timestamp 1649977179
transform 1 0 28244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_326
timestamp 1649977179
transform 1 0 31096 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_334
timestamp 1649977179
transform 1 0 31832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_340
timestamp 1649977179
transform 1 0 32384 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1649977179
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_372
timestamp 1649977179
transform 1 0 35328 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_392
timestamp 1649977179
transform 1 0 37168 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_398
timestamp 1649977179
transform 1 0 37720 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_404
timestamp 1649977179
transform 1 0 38272 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1649977179
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1649977179
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_423
timestamp 1649977179
transform 1 0 40020 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_435
timestamp 1649977179
transform 1 0 41124 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_447
timestamp 1649977179
transform 1 0 42228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_459
timestamp 1649977179
transform 1 0 43332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_471
timestamp 1649977179
transform 1 0 44436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1649977179
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1649977179
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1649977179
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1649977179
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1649977179
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1649977179
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1649977179
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1649977179
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1649977179
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1649977179
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1649977179
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1649977179
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1649977179
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_613
timestamp 1649977179
transform 1 0 57500 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_617
timestamp 1649977179
transform 1 0 57868 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_621
timestamp 1649977179
transform 1 0 58236 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_49
timestamp 1649977179
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_89
timestamp 1649977179
transform 1 0 9292 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1649977179
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_121
timestamp 1649977179
transform 1 0 12236 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_129
timestamp 1649977179
transform 1 0 12972 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_147
timestamp 1649977179
transform 1 0 14628 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_159
timestamp 1649977179
transform 1 0 15732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_189
timestamp 1649977179
transform 1 0 18492 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_195
timestamp 1649977179
transform 1 0 19044 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_203
timestamp 1649977179
transform 1 0 19780 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_209
timestamp 1649977179
transform 1 0 20332 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_214
timestamp 1649977179
transform 1 0 20792 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1649977179
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_227
timestamp 1649977179
transform 1 0 21988 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_238
timestamp 1649977179
transform 1 0 23000 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_248
timestamp 1649977179
transform 1 0 23920 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_272
timestamp 1649977179
transform 1 0 26128 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_291
timestamp 1649977179
transform 1 0 27876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_300
timestamp 1649977179
transform 1 0 28704 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_306
timestamp 1649977179
transform 1 0 29256 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_318
timestamp 1649977179
transform 1 0 30360 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_330
timestamp 1649977179
transform 1 0 31464 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_365
timestamp 1649977179
transform 1 0 34684 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_379
timestamp 1649977179
transform 1 0 35972 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_388
timestamp 1649977179
transform 1 0 36800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1649977179
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1649977179
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1649977179
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1649977179
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1649977179
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1649977179
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1649977179
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1649977179
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1649977179
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1649977179
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1649977179
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1649977179
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1649977179
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1649977179
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1649977179
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1649977179
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1649977179
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1649977179
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1649977179
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1649977179
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_37
timestamp 1649977179
transform 1 0 4508 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_47
timestamp 1649977179
transform 1 0 5428 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_59
timestamp 1649977179
transform 1 0 6532 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_67
timestamp 1649977179
transform 1 0 7268 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_78
timestamp 1649977179
transform 1 0 8280 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_87
timestamp 1649977179
transform 1 0 9108 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_95
timestamp 1649977179
transform 1 0 9844 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_107
timestamp 1649977179
transform 1 0 10948 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_119
timestamp 1649977179
transform 1 0 12052 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_131
timestamp 1649977179
transform 1 0 13156 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_145
timestamp 1649977179
transform 1 0 14444 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_157
timestamp 1649977179
transform 1 0 15548 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_167
timestamp 1649977179
transform 1 0 16468 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_187
timestamp 1649977179
transform 1 0 18308 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_199
timestamp 1649977179
transform 1 0 19412 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_206
timestamp 1649977179
transform 1 0 20056 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_220
timestamp 1649977179
transform 1 0 21344 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_227
timestamp 1649977179
transform 1 0 21988 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_242
timestamp 1649977179
transform 1 0 23368 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1649977179
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_255
timestamp 1649977179
transform 1 0 24564 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_259
timestamp 1649977179
transform 1 0 24932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_276
timestamp 1649977179
transform 1 0 26496 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_296
timestamp 1649977179
transform 1 0 28336 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_314
timestamp 1649977179
transform 1 0 29992 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_326
timestamp 1649977179
transform 1 0 31096 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_338
timestamp 1649977179
transform 1 0 32200 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_346
timestamp 1649977179
transform 1 0 32936 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_351
timestamp 1649977179
transform 1 0 33396 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_360
timestamp 1649977179
transform 1 0 34224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_375
timestamp 1649977179
transform 1 0 35604 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_382
timestamp 1649977179
transform 1 0 36248 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_386
timestamp 1649977179
transform 1 0 36616 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_397
timestamp 1649977179
transform 1 0 37628 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_408
timestamp 1649977179
transform 1 0 38640 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_416
timestamp 1649977179
transform 1 0 39376 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_421
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_429
timestamp 1649977179
transform 1 0 40572 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_441
timestamp 1649977179
transform 1 0 41676 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_453
timestamp 1649977179
transform 1 0 42780 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_465
timestamp 1649977179
transform 1 0 43884 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_473
timestamp 1649977179
transform 1 0 44620 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1649977179
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1649977179
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1649977179
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1649977179
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1649977179
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1649977179
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1649977179
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1649977179
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1649977179
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1649977179
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1649977179
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1649977179
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1649977179
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_613
timestamp 1649977179
transform 1 0 57500 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_617
timestamp 1649977179
transform 1 0 57868 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_621
timestamp 1649977179
transform 1 0 58236 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_11
timestamp 1649977179
transform 1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_30
timestamp 1649977179
transform 1 0 3864 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_63
timestamp 1649977179
transform 1 0 6900 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_86
timestamp 1649977179
transform 1 0 9016 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_102
timestamp 1649977179
transform 1 0 10488 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1649977179
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_133
timestamp 1649977179
transform 1 0 13340 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_141
timestamp 1649977179
transform 1 0 14076 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_153
timestamp 1649977179
transform 1 0 15180 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1649977179
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_173
timestamp 1649977179
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_177
timestamp 1649977179
transform 1 0 17388 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_183
timestamp 1649977179
transform 1 0 17940 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_203
timestamp 1649977179
transform 1 0 19780 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_214
timestamp 1649977179
transform 1 0 20792 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1649977179
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_230
timestamp 1649977179
transform 1 0 22264 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_241
timestamp 1649977179
transform 1 0 23276 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_248
timestamp 1649977179
transform 1 0 23920 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_254
timestamp 1649977179
transform 1 0 24472 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_266
timestamp 1649977179
transform 1 0 25576 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1649977179
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_286
timestamp 1649977179
transform 1 0 27416 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_298
timestamp 1649977179
transform 1 0 28520 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_306
timestamp 1649977179
transform 1 0 29256 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_318
timestamp 1649977179
transform 1 0 30360 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_330
timestamp 1649977179
transform 1 0 31464 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_343
timestamp 1649977179
transform 1 0 32660 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_354
timestamp 1649977179
transform 1 0 33672 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_362
timestamp 1649977179
transform 1 0 34408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_373
timestamp 1649977179
transform 1 0 35420 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_382
timestamp 1649977179
transform 1 0 36248 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_388
timestamp 1649977179
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_397
timestamp 1649977179
transform 1 0 37628 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_406
timestamp 1649977179
transform 1 0 38456 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_426
timestamp 1649977179
transform 1 0 40296 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_434
timestamp 1649977179
transform 1 0 41032 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_446
timestamp 1649977179
transform 1 0 42136 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1649977179
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1649977179
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1649977179
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1649977179
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1649977179
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1649977179
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1649977179
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1649977179
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1649977179
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1649977179
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1649977179
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1649977179
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1649977179
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1649977179
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1649977179
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1649977179
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1649977179
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_16
timestamp 1649977179
transform 1 0 2576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_20
timestamp 1649977179
transform 1 0 2944 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1649977179
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_45
timestamp 1649977179
transform 1 0 5244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_57
timestamp 1649977179
transform 1 0 6348 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_61
timestamp 1649977179
transform 1 0 6716 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_71
timestamp 1649977179
transform 1 0 7636 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1649977179
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_101
timestamp 1649977179
transform 1 0 10396 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_105
timestamp 1649977179
transform 1 0 10764 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_108
timestamp 1649977179
transform 1 0 11040 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_144
timestamp 1649977179
transform 1 0 14352 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_168
timestamp 1649977179
transform 1 0 16560 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1649977179
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_200
timestamp 1649977179
transform 1 0 19504 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_206
timestamp 1649977179
transform 1 0 20056 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_213
timestamp 1649977179
transform 1 0 20700 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_223
timestamp 1649977179
transform 1 0 21620 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_229
timestamp 1649977179
transform 1 0 22172 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_236
timestamp 1649977179
transform 1 0 22816 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_240
timestamp 1649977179
transform 1 0 23184 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_243
timestamp 1649977179
transform 1 0 23460 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_255
timestamp 1649977179
transform 1 0 24564 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_267
timestamp 1649977179
transform 1 0 25668 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_279
timestamp 1649977179
transform 1 0 26772 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_288
timestamp 1649977179
transform 1 0 27600 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_294
timestamp 1649977179
transform 1 0 28152 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1649977179
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_325
timestamp 1649977179
transform 1 0 31004 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_334
timestamp 1649977179
transform 1 0 31832 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_338
timestamp 1649977179
transform 1 0 32200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_341
timestamp 1649977179
transform 1 0 32476 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_359
timestamp 1649977179
transform 1 0 34132 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_367
timestamp 1649977179
transform 1 0 34868 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_383
timestamp 1649977179
transform 1 0 36340 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_400
timestamp 1649977179
transform 1 0 37904 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_406
timestamp 1649977179
transform 1 0 38456 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_412
timestamp 1649977179
transform 1 0 39008 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_429
timestamp 1649977179
transform 1 0 40572 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_435
timestamp 1649977179
transform 1 0 41124 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_447
timestamp 1649977179
transform 1 0 42228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_459
timestamp 1649977179
transform 1 0 43332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_471
timestamp 1649977179
transform 1 0 44436 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1649977179
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1649977179
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1649977179
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1649977179
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1649977179
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1649977179
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1649977179
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1649977179
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1649977179
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1649977179
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1649977179
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1649977179
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1649977179
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1649977179
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_8
timestamp 1649977179
transform 1 0 1840 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_32
timestamp 1649977179
transform 1 0 4048 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_38
timestamp 1649977179
transform 1 0 4600 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_50
timestamp 1649977179
transform 1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_73
timestamp 1649977179
transform 1 0 7820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_85
timestamp 1649977179
transform 1 0 8924 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_89
timestamp 1649977179
transform 1 0 9292 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_92
timestamp 1649977179
transform 1 0 9568 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_99
timestamp 1649977179
transform 1 0 10212 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_106
timestamp 1649977179
transform 1 0 10856 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_121
timestamp 1649977179
transform 1 0 12236 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_128
timestamp 1649977179
transform 1 0 12880 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_136
timestamp 1649977179
transform 1 0 13616 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_139
timestamp 1649977179
transform 1 0 13892 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_153
timestamp 1649977179
transform 1 0 15180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1649977179
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_175
timestamp 1649977179
transform 1 0 17204 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_184
timestamp 1649977179
transform 1 0 18032 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_197
timestamp 1649977179
transform 1 0 19228 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_208
timestamp 1649977179
transform 1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_215
timestamp 1649977179
transform 1 0 20884 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_227
timestamp 1649977179
transform 1 0 21988 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_234
timestamp 1649977179
transform 1 0 22632 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_250
timestamp 1649977179
transform 1 0 24104 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_258
timestamp 1649977179
transform 1 0 24840 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_267
timestamp 1649977179
transform 1 0 25668 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1649977179
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_286
timestamp 1649977179
transform 1 0 27416 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_294
timestamp 1649977179
transform 1 0 28152 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_298
timestamp 1649977179
transform 1 0 28520 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_310
timestamp 1649977179
transform 1 0 29624 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_324
timestamp 1649977179
transform 1 0 30912 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_331
timestamp 1649977179
transform 1 0 31556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_369
timestamp 1649977179
transform 1 0 35052 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_381
timestamp 1649977179
transform 1 0 36156 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_389
timestamp 1649977179
transform 1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_405
timestamp 1649977179
transform 1 0 38364 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_409
timestamp 1649977179
transform 1 0 38732 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_426
timestamp 1649977179
transform 1 0 40296 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_440
timestamp 1649977179
transform 1 0 41584 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1649977179
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1649977179
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1649977179
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1649977179
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1649977179
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1649977179
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1649977179
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1649977179
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1649977179
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1649977179
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1649977179
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1649977179
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1649977179
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_617
timestamp 1649977179
transform 1 0 57868 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_621
timestamp 1649977179
transform 1 0 58236 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_7
timestamp 1649977179
transform 1 0 1748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1649977179
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_37
timestamp 1649977179
transform 1 0 4508 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_43
timestamp 1649977179
transform 1 0 5060 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_55
timestamp 1649977179
transform 1 0 6164 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_63
timestamp 1649977179
transform 1 0 6900 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1649977179
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_103
timestamp 1649977179
transform 1 0 10580 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_115
timestamp 1649977179
transform 1 0 11684 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_127
timestamp 1649977179
transform 1 0 12788 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_151
timestamp 1649977179
transform 1 0 14996 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1649977179
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_175
timestamp 1649977179
transform 1 0 17204 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_187
timestamp 1649977179
transform 1 0 18308 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_199
timestamp 1649977179
transform 1 0 19412 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_207
timestamp 1649977179
transform 1 0 20148 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1649977179
transform 1 0 20424 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_216
timestamp 1649977179
transform 1 0 20976 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_228
timestamp 1649977179
transform 1 0 22080 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_240
timestamp 1649977179
transform 1 0 23184 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_257
timestamp 1649977179
transform 1 0 24748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_264
timestamp 1649977179
transform 1 0 25392 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_280
timestamp 1649977179
transform 1 0 26864 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_291
timestamp 1649977179
transform 1 0 27876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_303
timestamp 1649977179
transform 1 0 28980 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_326
timestamp 1649977179
transform 1 0 31096 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_340
timestamp 1649977179
transform 1 0 32384 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_360
timestamp 1649977179
transform 1 0 34224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_373
timestamp 1649977179
transform 1 0 35420 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_376
timestamp 1649977179
transform 1 0 35696 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_384
timestamp 1649977179
transform 1 0 36432 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_395
timestamp 1649977179
transform 1 0 37444 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_407
timestamp 1649977179
transform 1 0 38548 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_411
timestamp 1649977179
transform 1 0 38916 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_416
timestamp 1649977179
transform 1 0 39376 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_426
timestamp 1649977179
transform 1 0 40296 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_438
timestamp 1649977179
transform 1 0 41400 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_450
timestamp 1649977179
transform 1 0 42504 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_462
timestamp 1649977179
transform 1 0 43608 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_474
timestamp 1649977179
transform 1 0 44712 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1649977179
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1649977179
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1649977179
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1649977179
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1649977179
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1649977179
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1649977179
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1649977179
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1649977179
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1649977179
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1649977179
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1649977179
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1649977179
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1649977179
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_37
timestamp 1649977179
transform 1 0 4508 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_43
timestamp 1649977179
transform 1 0 5060 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_46
timestamp 1649977179
transform 1 0 5336 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1649977179
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_67
timestamp 1649977179
transform 1 0 7268 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_79
timestamp 1649977179
transform 1 0 8372 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_91
timestamp 1649977179
transform 1 0 9476 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1649977179
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_118
timestamp 1649977179
transform 1 0 11960 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_124
timestamp 1649977179
transform 1 0 12512 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_130
timestamp 1649977179
transform 1 0 13064 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_138
timestamp 1649977179
transform 1 0 13800 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_144
timestamp 1649977179
transform 1 0 14352 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_160
timestamp 1649977179
transform 1 0 15824 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_171
timestamp 1649977179
transform 1 0 16836 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_179
timestamp 1649977179
transform 1 0 17572 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_191
timestamp 1649977179
transform 1 0 18676 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_203
timestamp 1649977179
transform 1 0 19780 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_215
timestamp 1649977179
transform 1 0 20884 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1649977179
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_233
timestamp 1649977179
transform 1 0 22540 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_239
timestamp 1649977179
transform 1 0 23092 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_255
timestamp 1649977179
transform 1 0 24564 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_263
timestamp 1649977179
transform 1 0 25300 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_275
timestamp 1649977179
transform 1 0 26404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_297
timestamp 1649977179
transform 1 0 28428 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_309
timestamp 1649977179
transform 1 0 29532 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1649977179
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_329
timestamp 1649977179
transform 1 0 31372 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1649977179
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_349
timestamp 1649977179
transform 1 0 33212 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_369
timestamp 1649977179
transform 1 0 35052 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_375
timestamp 1649977179
transform 1 0 35604 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_384
timestamp 1649977179
transform 1 0 36432 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_398
timestamp 1649977179
transform 1 0 37720 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_402
timestamp 1649977179
transform 1 0 38088 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_413
timestamp 1649977179
transform 1 0 39100 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_425
timestamp 1649977179
transform 1 0 40204 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_437
timestamp 1649977179
transform 1 0 41308 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_445
timestamp 1649977179
transform 1 0 42044 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1649977179
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1649977179
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1649977179
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1649977179
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1649977179
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1649977179
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1649977179
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1649977179
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1649977179
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1649977179
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1649977179
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1649977179
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1649977179
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1649977179
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1649977179
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1649977179
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_617
timestamp 1649977179
transform 1 0 57868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_621
timestamp 1649977179
transform 1 0 58236 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_16
timestamp 1649977179
transform 1 0 2576 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1649977179
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_34
timestamp 1649977179
transform 1 0 4232 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_42
timestamp 1649977179
transform 1 0 4968 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_52
timestamp 1649977179
transform 1 0 5888 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_66
timestamp 1649977179
transform 1 0 7176 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_72
timestamp 1649977179
transform 1 0 7728 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_123
timestamp 1649977179
transform 1 0 12420 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_135
timestamp 1649977179
transform 1 0 13524 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_157
timestamp 1649977179
transform 1 0 15548 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_169
timestamp 1649977179
transform 1 0 16652 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_181
timestamp 1649977179
transform 1 0 17756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1649977179
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_205
timestamp 1649977179
transform 1 0 19964 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_214
timestamp 1649977179
transform 1 0 20792 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_234
timestamp 1649977179
transform 1 0 22632 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1649977179
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1649977179
transform 1 0 26036 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_280
timestamp 1649977179
transform 1 0 26864 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_292
timestamp 1649977179
transform 1 0 27968 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1649977179
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_330
timestamp 1649977179
transform 1 0 31464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_334
timestamp 1649977179
transform 1 0 31832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_340
timestamp 1649977179
transform 1 0 32384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_352
timestamp 1649977179
transform 1 0 33488 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_358
timestamp 1649977179
transform 1 0 34040 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_377
timestamp 1649977179
transform 1 0 35788 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_396
timestamp 1649977179
transform 1 0 37536 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_410
timestamp 1649977179
transform 1 0 38824 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_418
timestamp 1649977179
transform 1 0 39560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_421
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_432
timestamp 1649977179
transform 1 0 40848 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_438
timestamp 1649977179
transform 1 0 41400 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_450
timestamp 1649977179
transform 1 0 42504 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_462
timestamp 1649977179
transform 1 0 43608 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_474
timestamp 1649977179
transform 1 0 44712 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1649977179
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1649977179
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1649977179
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1649977179
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1649977179
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1649977179
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1649977179
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1649977179
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1649977179
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1649977179
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1649977179
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1649977179
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1649977179
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1649977179
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_9
timestamp 1649977179
transform 1 0 1932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_18
timestamp 1649977179
transform 1 0 2760 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_33
timestamp 1649977179
transform 1 0 4140 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_45
timestamp 1649977179
transform 1 0 5244 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_49
timestamp 1649977179
transform 1 0 5612 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1649977179
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_77
timestamp 1649977179
transform 1 0 8188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_85
timestamp 1649977179
transform 1 0 8924 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_90
timestamp 1649977179
transform 1 0 9384 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_96
timestamp 1649977179
transform 1 0 9936 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1649977179
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_118
timestamp 1649977179
transform 1 0 11960 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_124
timestamp 1649977179
transform 1 0 12512 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_127
timestamp 1649977179
transform 1 0 12788 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_139
timestamp 1649977179
transform 1 0 13892 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_151
timestamp 1649977179
transform 1 0 14996 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1649977179
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_178
timestamp 1649977179
transform 1 0 17480 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_190
timestamp 1649977179
transform 1 0 18584 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_199
timestamp 1649977179
transform 1 0 19412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_211
timestamp 1649977179
transform 1 0 20516 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_215
timestamp 1649977179
transform 1 0 20884 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1649977179
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_230
timestamp 1649977179
transform 1 0 22264 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_236
timestamp 1649977179
transform 1 0 22816 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_240
timestamp 1649977179
transform 1 0 23184 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_245
timestamp 1649977179
transform 1 0 23644 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_253
timestamp 1649977179
transform 1 0 24380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_301
timestamp 1649977179
transform 1 0 28796 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_305
timestamp 1649977179
transform 1 0 29164 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_313
timestamp 1649977179
transform 1 0 29900 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_325
timestamp 1649977179
transform 1 0 31004 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_333
timestamp 1649977179
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_342
timestamp 1649977179
transform 1 0 32568 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_351
timestamp 1649977179
transform 1 0 33396 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_363
timestamp 1649977179
transform 1 0 34500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_375
timestamp 1649977179
transform 1 0 35604 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_388
timestamp 1649977179
transform 1 0 36800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_399
timestamp 1649977179
transform 1 0 37812 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_404
timestamp 1649977179
transform 1 0 38272 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_410
timestamp 1649977179
transform 1 0 38824 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_427
timestamp 1649977179
transform 1 0 40388 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_439
timestamp 1649977179
transform 1 0 41492 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1649977179
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1649977179
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1649977179
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1649977179
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1649977179
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1649977179
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1649977179
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1649977179
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1649977179
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1649977179
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1649977179
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1649977179
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1649977179
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1649977179
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1649977179
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1649977179
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1649977179
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_617
timestamp 1649977179
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_7
timestamp 1649977179
transform 1 0 1748 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1649977179
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_38
timestamp 1649977179
transform 1 0 4600 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_50
timestamp 1649977179
transform 1 0 5704 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_54
timestamp 1649977179
transform 1 0 6072 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_59
timestamp 1649977179
transform 1 0 6532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_72
timestamp 1649977179
transform 1 0 7728 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_78
timestamp 1649977179
transform 1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1649977179
transform 1 0 9476 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_108
timestamp 1649977179
transform 1 0 11040 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_120
timestamp 1649977179
transform 1 0 12144 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_126
timestamp 1649977179
transform 1 0 12696 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1649977179
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_159
timestamp 1649977179
transform 1 0 15732 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_162
timestamp 1649977179
transform 1 0 16008 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_174
timestamp 1649977179
transform 1 0 17112 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_180
timestamp 1649977179
transform 1 0 17664 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1649977179
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_213
timestamp 1649977179
transform 1 0 20700 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_227
timestamp 1649977179
transform 1 0 21988 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_235
timestamp 1649977179
transform 1 0 22724 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1649977179
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_280
timestamp 1649977179
transform 1 0 26864 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_288
timestamp 1649977179
transform 1 0 27600 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_300
timestamp 1649977179
transform 1 0 28704 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_316
timestamp 1649977179
transform 1 0 30176 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_326
timestamp 1649977179
transform 1 0 31096 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_330
timestamp 1649977179
transform 1 0 31464 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_333
timestamp 1649977179
transform 1 0 31740 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1649977179
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1649977179
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_389
timestamp 1649977179
transform 1 0 36892 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_400
timestamp 1649977179
transform 1 0 37904 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_412
timestamp 1649977179
transform 1 0 39008 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_426
timestamp 1649977179
transform 1 0 40296 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_432
timestamp 1649977179
transform 1 0 40848 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_438
timestamp 1649977179
transform 1 0 41400 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_441
timestamp 1649977179
transform 1 0 41676 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_453
timestamp 1649977179
transform 1 0 42780 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_465
timestamp 1649977179
transform 1 0 43884 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_473
timestamp 1649977179
transform 1 0 44620 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1649977179
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1649977179
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1649977179
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1649977179
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1649977179
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1649977179
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1649977179
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1649977179
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1649977179
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1649977179
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1649977179
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1649977179
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1649977179
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_613
timestamp 1649977179
transform 1 0 57500 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_617
timestamp 1649977179
transform 1 0 57868 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_621
timestamp 1649977179
transform 1 0 58236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_11
timestamp 1649977179
transform 1 0 2116 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_35
timestamp 1649977179
transform 1 0 4324 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_49
timestamp 1649977179
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_61
timestamp 1649977179
transform 1 0 6716 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_74
timestamp 1649977179
transform 1 0 7912 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_83
timestamp 1649977179
transform 1 0 8740 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_89
timestamp 1649977179
transform 1 0 9292 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_101
timestamp 1649977179
transform 1 0 10396 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1649977179
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_115
timestamp 1649977179
transform 1 0 11684 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_127
timestamp 1649977179
transform 1 0 12788 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_139
timestamp 1649977179
transform 1 0 13892 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_143
timestamp 1649977179
transform 1 0 14260 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_185
timestamp 1649977179
transform 1 0 18124 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_197
timestamp 1649977179
transform 1 0 19228 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_209
timestamp 1649977179
transform 1 0 20332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_221
timestamp 1649977179
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_229
timestamp 1649977179
transform 1 0 22172 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_235
timestamp 1649977179
transform 1 0 22724 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_247
timestamp 1649977179
transform 1 0 23828 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_259
timestamp 1649977179
transform 1 0 24932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_263
timestamp 1649977179
transform 1 0 25300 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_271
timestamp 1649977179
transform 1 0 26036 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_287
timestamp 1649977179
transform 1 0 27508 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_299
timestamp 1649977179
transform 1 0 28612 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_307
timestamp 1649977179
transform 1 0 29348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_316
timestamp 1649977179
transform 1 0 30176 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_326
timestamp 1649977179
transform 1 0 31096 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1649977179
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_354
timestamp 1649977179
transform 1 0 33672 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_366
timestamp 1649977179
transform 1 0 34776 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1649977179
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1649977179
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_397
timestamp 1649977179
transform 1 0 37628 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_421
timestamp 1649977179
transform 1 0 39836 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_437
timestamp 1649977179
transform 1 0 41308 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_445
timestamp 1649977179
transform 1 0 42044 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1649977179
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1649977179
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1649977179
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1649977179
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1649977179
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1649977179
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1649977179
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1649977179
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1649977179
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1649977179
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1649977179
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1649977179
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1649977179
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1649977179
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1649977179
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1649977179
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1649977179
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1649977179
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1649977179
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_37
timestamp 1649977179
transform 1 0 4508 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_40
timestamp 1649977179
transform 1 0 4784 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_54
timestamp 1649977179
transform 1 0 6072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_60
timestamp 1649977179
transform 1 0 6624 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1649977179
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_117
timestamp 1649977179
transform 1 0 11868 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_120
timestamp 1649977179
transform 1 0 12144 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_132
timestamp 1649977179
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_145
timestamp 1649977179
transform 1 0 14444 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_151
timestamp 1649977179
transform 1 0 14996 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_163
timestamp 1649977179
transform 1 0 16100 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_175
timestamp 1649977179
transform 1 0 17204 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_187
timestamp 1649977179
transform 1 0 18308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_208
timestamp 1649977179
transform 1 0 20240 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_220
timestamp 1649977179
transform 1 0 21344 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_232
timestamp 1649977179
transform 1 0 22448 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_240
timestamp 1649977179
transform 1 0 23184 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_246
timestamp 1649977179
transform 1 0 23736 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_282
timestamp 1649977179
transform 1 0 27048 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_288
timestamp 1649977179
transform 1 0 27600 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_296
timestamp 1649977179
transform 1 0 28336 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1649977179
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_320
timestamp 1649977179
transform 1 0 30544 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_331
timestamp 1649977179
transform 1 0 31556 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_343
timestamp 1649977179
transform 1 0 32660 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_349
timestamp 1649977179
transform 1 0 33212 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_361
timestamp 1649977179
transform 1 0 34316 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_369
timestamp 1649977179
transform 1 0 35052 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_377
timestamp 1649977179
transform 1 0 35788 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_391
timestamp 1649977179
transform 1 0 37076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_399
timestamp 1649977179
transform 1 0 37812 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_416
timestamp 1649977179
transform 1 0 39376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_421
timestamp 1649977179
transform 1 0 39836 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_430
timestamp 1649977179
transform 1 0 40664 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_442
timestamp 1649977179
transform 1 0 41768 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_454
timestamp 1649977179
transform 1 0 42872 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_466
timestamp 1649977179
transform 1 0 43976 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_474
timestamp 1649977179
transform 1 0 44712 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1649977179
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1649977179
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1649977179
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1649977179
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1649977179
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1649977179
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1649977179
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1649977179
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1649977179
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1649977179
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1649977179
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1649977179
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1649977179
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_613
timestamp 1649977179
transform 1 0 57500 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_617
timestamp 1649977179
transform 1 0 57868 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_621
timestamp 1649977179
transform 1 0 58236 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1649977179
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_75
timestamp 1649977179
transform 1 0 8004 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_87
timestamp 1649977179
transform 1 0 9108 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_99
timestamp 1649977179
transform 1 0 10212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_115
timestamp 1649977179
transform 1 0 11684 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_151
timestamp 1649977179
transform 1 0 14996 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_155
timestamp 1649977179
transform 1 0 15364 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_160
timestamp 1649977179
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_182
timestamp 1649977179
transform 1 0 17848 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_194
timestamp 1649977179
transform 1 0 18952 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_202
timestamp 1649977179
transform 1 0 19688 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_212
timestamp 1649977179
transform 1 0 20608 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_254
timestamp 1649977179
transform 1 0 24472 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_264
timestamp 1649977179
transform 1 0 25392 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1649977179
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_285
timestamp 1649977179
transform 1 0 27324 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_290
timestamp 1649977179
transform 1 0 27784 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_300
timestamp 1649977179
transform 1 0 28704 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_308
timestamp 1649977179
transform 1 0 29440 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_322
timestamp 1649977179
transform 1 0 30728 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1649977179
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_349
timestamp 1649977179
transform 1 0 33212 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_369
timestamp 1649977179
transform 1 0 35052 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_377
timestamp 1649977179
transform 1 0 35788 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_388
timestamp 1649977179
transform 1 0 36800 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1649977179
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_417
timestamp 1649977179
transform 1 0 39468 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_421
timestamp 1649977179
transform 1 0 39836 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_424
timestamp 1649977179
transform 1 0 40112 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_436
timestamp 1649977179
transform 1 0 41216 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1649977179
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1649977179
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1649977179
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1649977179
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1649977179
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1649977179
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1649977179
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1649977179
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1649977179
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1649977179
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1649977179
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1649977179
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1649977179
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1649977179
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1649977179
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1649977179
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1649977179
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1649977179
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_19
timestamp 1649977179
transform 1 0 2852 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_22
timestamp 1649977179
transform 1 0 3128 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_100
timestamp 1649977179
transform 1 0 10304 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_108
timestamp 1649977179
transform 1 0 11040 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_116
timestamp 1649977179
transform 1 0 11776 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_122
timestamp 1649977179
transform 1 0 12328 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_126
timestamp 1649977179
transform 1 0 12696 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_132
timestamp 1649977179
transform 1 0 13248 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_149
timestamp 1649977179
transform 1 0 14812 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_163
timestamp 1649977179
transform 1 0 16100 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_169
timestamp 1649977179
transform 1 0 16652 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_181
timestamp 1649977179
transform 1 0 17756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 1649977179
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_213
timestamp 1649977179
transform 1 0 20700 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_221
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_225
timestamp 1649977179
transform 1 0 21804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_228
timestamp 1649977179
transform 1 0 22080 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_248
timestamp 1649977179
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_269
timestamp 1649977179
transform 1 0 25852 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_275
timestamp 1649977179
transform 1 0 26404 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_283
timestamp 1649977179
transform 1 0 27140 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_286
timestamp 1649977179
transform 1 0 27416 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_298
timestamp 1649977179
transform 1 0 28520 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 1649977179
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_316
timestamp 1649977179
transform 1 0 30176 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_328
timestamp 1649977179
transform 1 0 31280 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_336
timestamp 1649977179
transform 1 0 32016 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_341
timestamp 1649977179
transform 1 0 32476 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_353
timestamp 1649977179
transform 1 0 33580 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_361
timestamp 1649977179
transform 1 0 34316 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_392
timestamp 1649977179
transform 1 0 37168 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_416
timestamp 1649977179
transform 1 0 39376 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_421
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_430
timestamp 1649977179
transform 1 0 40664 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_442
timestamp 1649977179
transform 1 0 41768 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_454
timestamp 1649977179
transform 1 0 42872 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_466
timestamp 1649977179
transform 1 0 43976 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_474
timestamp 1649977179
transform 1 0 44712 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1649977179
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1649977179
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1649977179
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1649977179
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1649977179
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1649977179
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1649977179
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1649977179
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1649977179
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1649977179
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1649977179
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1649977179
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1649977179
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1649977179
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1649977179
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_11
timestamp 1649977179
transform 1 0 2116 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_20
timestamp 1649977179
transform 1 0 2944 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_28
timestamp 1649977179
transform 1 0 3680 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_34
timestamp 1649977179
transform 1 0 4232 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_46
timestamp 1649977179
transform 1 0 5336 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1649977179
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_65
timestamp 1649977179
transform 1 0 7084 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_71
timestamp 1649977179
transform 1 0 7636 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_83
timestamp 1649977179
transform 1 0 8740 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_87
timestamp 1649977179
transform 1 0 9108 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_95
timestamp 1649977179
transform 1 0 9844 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_103
timestamp 1649977179
transform 1 0 10580 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_123
timestamp 1649977179
transform 1 0 12420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_135
timestamp 1649977179
transform 1 0 13524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_143
timestamp 1649977179
transform 1 0 14260 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_150
timestamp 1649977179
transform 1 0 14904 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_159
timestamp 1649977179
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_185
timestamp 1649977179
transform 1 0 18124 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_194
timestamp 1649977179
transform 1 0 18952 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_202
timestamp 1649977179
transform 1 0 19688 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_211
timestamp 1649977179
transform 1 0 20516 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_215
timestamp 1649977179
transform 1 0 20884 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1649977179
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_230
timestamp 1649977179
transform 1 0 22264 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_242
timestamp 1649977179
transform 1 0 23368 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_251
timestamp 1649977179
transform 1 0 24196 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_255
timestamp 1649977179
transform 1 0 24564 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1649977179
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_283
timestamp 1649977179
transform 1 0 27140 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_289
timestamp 1649977179
transform 1 0 27692 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_301
timestamp 1649977179
transform 1 0 28796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_307
timestamp 1649977179
transform 1 0 29348 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_319
timestamp 1649977179
transform 1 0 30452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_331
timestamp 1649977179
transform 1 0 31556 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_343
timestamp 1649977179
transform 1 0 32660 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_353
timestamp 1649977179
transform 1 0 33580 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_365
timestamp 1649977179
transform 1 0 34684 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_377
timestamp 1649977179
transform 1 0 35788 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_389
timestamp 1649977179
transform 1 0 36892 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1649977179
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_423
timestamp 1649977179
transform 1 0 40020 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_435
timestamp 1649977179
transform 1 0 41124 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1649977179
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1649977179
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1649977179
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1649977179
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1649977179
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1649977179
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1649977179
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1649977179
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1649977179
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1649977179
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1649977179
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1649977179
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1649977179
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1649977179
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1649977179
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1649977179
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1649977179
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1649977179
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1649977179
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_617
timestamp 1649977179
transform 1 0 57868 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_621
timestamp 1649977179
transform 1 0 58236 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_7
timestamp 1649977179
transform 1 0 1748 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1649977179
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_45
timestamp 1649977179
transform 1 0 5244 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_69
timestamp 1649977179
transform 1 0 7452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_81
timestamp 1649977179
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_91
timestamp 1649977179
transform 1 0 9476 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_102
timestamp 1649977179
transform 1 0 10488 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_117
timestamp 1649977179
transform 1 0 11868 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_129
timestamp 1649977179
transform 1 0 12972 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_137
timestamp 1649977179
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_151
timestamp 1649977179
transform 1 0 14996 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_160
timestamp 1649977179
transform 1 0 15824 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_174
timestamp 1649977179
transform 1 0 17112 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_190
timestamp 1649977179
transform 1 0 18584 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_206
timestamp 1649977179
transform 1 0 20056 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_210
timestamp 1649977179
transform 1 0 20424 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_231
timestamp 1649977179
transform 1 0 22356 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_243
timestamp 1649977179
transform 1 0 23460 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_257
timestamp 1649977179
transform 1 0 24748 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_269
timestamp 1649977179
transform 1 0 25852 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_281
timestamp 1649977179
transform 1 0 26956 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_293
timestamp 1649977179
transform 1 0 28060 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_300
timestamp 1649977179
transform 1 0 28704 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_343
timestamp 1649977179
transform 1 0 32660 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_353
timestamp 1649977179
transform 1 0 33580 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_361
timestamp 1649977179
transform 1 0 34316 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_391
timestamp 1649977179
transform 1 0 37076 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_397
timestamp 1649977179
transform 1 0 37628 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_409
timestamp 1649977179
transform 1 0 38732 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_417
timestamp 1649977179
transform 1 0 39468 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_421
timestamp 1649977179
transform 1 0 39836 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_427
timestamp 1649977179
transform 1 0 40388 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_439
timestamp 1649977179
transform 1 0 41492 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_451
timestamp 1649977179
transform 1 0 42596 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_463
timestamp 1649977179
transform 1 0 43700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1649977179
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1649977179
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1649977179
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1649977179
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1649977179
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1649977179
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1649977179
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1649977179
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1649977179
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1649977179
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1649977179
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1649977179
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1649977179
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1649977179
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1649977179
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1649977179
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_10
timestamp 1649977179
transform 1 0 2024 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_30
timestamp 1649977179
transform 1 0 3864 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_42
timestamp 1649977179
transform 1 0 4968 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1649977179
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_62
timestamp 1649977179
transform 1 0 6808 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_75
timestamp 1649977179
transform 1 0 8004 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_87
timestamp 1649977179
transform 1 0 9108 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_95
timestamp 1649977179
transform 1 0 9844 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_99
timestamp 1649977179
transform 1 0 10212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_115
timestamp 1649977179
transform 1 0 11684 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_127
timestamp 1649977179
transform 1 0 12788 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_139
timestamp 1649977179
transform 1 0 13892 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_150
timestamp 1649977179
transform 1 0 14904 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_156
timestamp 1649977179
transform 1 0 15456 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_162
timestamp 1649977179
transform 1 0 16008 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_171
timestamp 1649977179
transform 1 0 16836 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_179
timestamp 1649977179
transform 1 0 17572 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_182
timestamp 1649977179
transform 1 0 17848 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_202
timestamp 1649977179
transform 1 0 19688 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_214
timestamp 1649977179
transform 1 0 20792 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1649977179
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_230
timestamp 1649977179
transform 1 0 22264 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_236
timestamp 1649977179
transform 1 0 22816 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_242
timestamp 1649977179
transform 1 0 23368 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_246
timestamp 1649977179
transform 1 0 23736 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_257
timestamp 1649977179
transform 1 0 24748 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_269
timestamp 1649977179
transform 1 0 25852 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1649977179
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1649977179
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1649977179
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1649977179
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_339
timestamp 1649977179
transform 1 0 32292 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_351
timestamp 1649977179
transform 1 0 33396 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_362
timestamp 1649977179
transform 1 0 34408 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_372
timestamp 1649977179
transform 1 0 35328 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_383
timestamp 1649977179
transform 1 0 36340 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1649977179
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_401
timestamp 1649977179
transform 1 0 37996 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_425
timestamp 1649977179
transform 1 0 40204 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_437
timestamp 1649977179
transform 1 0 41308 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_445
timestamp 1649977179
transform 1 0 42044 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1649977179
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1649977179
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1649977179
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1649977179
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1649977179
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1649977179
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1649977179
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1649977179
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1649977179
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1649977179
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1649977179
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1649977179
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1649977179
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1649977179
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1649977179
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1649977179
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1649977179
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_617
timestamp 1649977179
transform 1 0 57868 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_621
timestamp 1649977179
transform 1 0 58236 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_11
timestamp 1649977179
transform 1 0 2116 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1649977179
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_31
timestamp 1649977179
transform 1 0 3956 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_39
timestamp 1649977179
transform 1 0 4692 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_42
timestamp 1649977179
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_54
timestamp 1649977179
transform 1 0 6072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_74
timestamp 1649977179
transform 1 0 7912 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1649977179
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_93
timestamp 1649977179
transform 1 0 9660 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_100
timestamp 1649977179
transform 1 0 10304 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_113
timestamp 1649977179
transform 1 0 11500 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_122
timestamp 1649977179
transform 1 0 12328 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_134
timestamp 1649977179
transform 1 0 13432 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_147
timestamp 1649977179
transform 1 0 14628 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_171
timestamp 1649977179
transform 1 0 16836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_183
timestamp 1649977179
transform 1 0 17940 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1649977179
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1649977179
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_221
timestamp 1649977179
transform 1 0 21436 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_229
timestamp 1649977179
transform 1 0 22172 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_237
timestamp 1649977179
transform 1 0 22908 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_245
timestamp 1649977179
transform 1 0 23644 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1649977179
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_261
timestamp 1649977179
transform 1 0 25116 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_282
timestamp 1649977179
transform 1 0 27048 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_294
timestamp 1649977179
transform 1 0 28152 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_306
timestamp 1649977179
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_311
timestamp 1649977179
transform 1 0 29716 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_323
timestamp 1649977179
transform 1 0 30820 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_331
timestamp 1649977179
transform 1 0 31556 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_340
timestamp 1649977179
transform 1 0 32384 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1649977179
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_369
timestamp 1649977179
transform 1 0 35052 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_377
timestamp 1649977179
transform 1 0 35788 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_397
timestamp 1649977179
transform 1 0 37628 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_409
timestamp 1649977179
transform 1 0 38732 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_413
timestamp 1649977179
transform 1 0 39100 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_416
timestamp 1649977179
transform 1 0 39376 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_421
timestamp 1649977179
transform 1 0 39836 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_425
timestamp 1649977179
transform 1 0 40204 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_434
timestamp 1649977179
transform 1 0 41032 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_446
timestamp 1649977179
transform 1 0 42136 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_458
timestamp 1649977179
transform 1 0 43240 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_470
timestamp 1649977179
transform 1 0 44344 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1649977179
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1649977179
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1649977179
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1649977179
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1649977179
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1649977179
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1649977179
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1649977179
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1649977179
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1649977179
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1649977179
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1649977179
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1649977179
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1649977179
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1649977179
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_16
timestamp 1649977179
transform 1 0 2576 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_28
timestamp 1649977179
transform 1 0 3680 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_40
timestamp 1649977179
transform 1 0 4784 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1649977179
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_59
timestamp 1649977179
transform 1 0 6532 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_63
timestamp 1649977179
transform 1 0 6900 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_74
timestamp 1649977179
transform 1 0 7912 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_78
timestamp 1649977179
transform 1 0 8280 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_95
timestamp 1649977179
transform 1 0 9844 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_107
timestamp 1649977179
transform 1 0 10948 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_129
timestamp 1649977179
transform 1 0 12972 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_138
timestamp 1649977179
transform 1 0 13800 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_146
timestamp 1649977179
transform 1 0 14536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_157
timestamp 1649977179
transform 1 0 15548 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_163
timestamp 1649977179
transform 1 0 16100 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_181
timestamp 1649977179
transform 1 0 17756 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_187
timestamp 1649977179
transform 1 0 18308 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1649977179
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1649977179
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1649977179
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1649977179
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_231
timestamp 1649977179
transform 1 0 22356 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_240
timestamp 1649977179
transform 1 0 23184 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_252
timestamp 1649977179
transform 1 0 24288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_256
timestamp 1649977179
transform 1 0 24656 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1649977179
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_286
timestamp 1649977179
transform 1 0 27416 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_298
timestamp 1649977179
transform 1 0 28520 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_304
timestamp 1649977179
transform 1 0 29072 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_316
timestamp 1649977179
transform 1 0 30176 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_322
timestamp 1649977179
transform 1 0 30728 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1649977179
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1649977179
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1649977179
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_373
timestamp 1649977179
transform 1 0 35420 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_383
timestamp 1649977179
transform 1 0 36340 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1649977179
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_398
timestamp 1649977179
transform 1 0 37720 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_406
timestamp 1649977179
transform 1 0 38456 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_425
timestamp 1649977179
transform 1 0 40204 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_437
timestamp 1649977179
transform 1 0 41308 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_443
timestamp 1649977179
transform 1 0 41860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1649977179
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1649977179
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1649977179
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1649977179
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1649977179
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1649977179
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1649977179
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1649977179
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1649977179
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1649977179
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1649977179
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1649977179
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1649977179
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1649977179
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1649977179
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1649977179
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1649977179
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1649977179
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_617
timestamp 1649977179
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_67
timestamp 1649977179
transform 1 0 7268 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_73
timestamp 1649977179
transform 1 0 7820 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_76
timestamp 1649977179
transform 1 0 8096 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_101
timestamp 1649977179
transform 1 0 10396 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_107
timestamp 1649977179
transform 1 0 10948 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_116
timestamp 1649977179
transform 1 0 11776 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1649977179
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_151
timestamp 1649977179
transform 1 0 14996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_159
timestamp 1649977179
transform 1 0 15732 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_171
timestamp 1649977179
transform 1 0 16836 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_188
timestamp 1649977179
transform 1 0 18400 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_202
timestamp 1649977179
transform 1 0 19688 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_222
timestamp 1649977179
transform 1 0 21528 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_234
timestamp 1649977179
transform 1 0 22632 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_246
timestamp 1649977179
transform 1 0 23736 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_264
timestamp 1649977179
transform 1 0 25392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_276
timestamp 1649977179
transform 1 0 26496 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_286
timestamp 1649977179
transform 1 0 27416 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_292
timestamp 1649977179
transform 1 0 27968 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1649977179
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_311
timestamp 1649977179
transform 1 0 29716 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_323
timestamp 1649977179
transform 1 0 30820 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_329
timestamp 1649977179
transform 1 0 31372 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_341
timestamp 1649977179
transform 1 0 32476 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_353
timestamp 1649977179
transform 1 0 33580 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1649977179
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_383
timestamp 1649977179
transform 1 0 36340 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1649977179
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1649977179
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1649977179
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_421
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_425
timestamp 1649977179
transform 1 0 40204 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_431
timestamp 1649977179
transform 1 0 40756 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_440
timestamp 1649977179
transform 1 0 41584 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_452
timestamp 1649977179
transform 1 0 42688 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_464
timestamp 1649977179
transform 1 0 43792 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1649977179
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1649977179
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1649977179
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1649977179
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1649977179
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1649977179
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1649977179
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1649977179
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1649977179
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1649977179
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1649977179
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1649977179
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1649977179
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1649977179
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_613
timestamp 1649977179
transform 1 0 57500 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_617
timestamp 1649977179
transform 1 0 57868 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_621
timestamp 1649977179
transform 1 0 58236 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_31
timestamp 1649977179
transform 1 0 3956 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_41
timestamp 1649977179
transform 1 0 4876 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_47
timestamp 1649977179
transform 1 0 5428 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_65
timestamp 1649977179
transform 1 0 7084 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_87
timestamp 1649977179
transform 1 0 9108 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_90
timestamp 1649977179
transform 1 0 9384 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_102
timestamp 1649977179
transform 1 0 10488 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1649977179
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_115
timestamp 1649977179
transform 1 0 11684 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_121
timestamp 1649977179
transform 1 0 12236 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_133
timestamp 1649977179
transform 1 0 13340 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_137
timestamp 1649977179
transform 1 0 13708 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_140
timestamp 1649977179
transform 1 0 13984 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_160
timestamp 1649977179
transform 1 0 15824 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_173
timestamp 1649977179
transform 1 0 17020 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_187
timestamp 1649977179
transform 1 0 18308 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_207
timestamp 1649977179
transform 1 0 20148 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_215
timestamp 1649977179
transform 1 0 20884 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1649977179
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_233
timestamp 1649977179
transform 1 0 22540 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_245
timestamp 1649977179
transform 1 0 23644 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_257
timestamp 1649977179
transform 1 0 24748 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_265
timestamp 1649977179
transform 1 0 25484 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_268
timestamp 1649977179
transform 1 0 25760 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_274
timestamp 1649977179
transform 1 0 26312 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_293
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_302
timestamp 1649977179
transform 1 0 28888 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_322
timestamp 1649977179
transform 1 0 30728 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_334
timestamp 1649977179
transform 1 0 31832 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1649977179
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1649977179
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1649977179
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1649977179
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1649977179
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_395
timestamp 1649977179
transform 1 0 37444 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_403
timestamp 1649977179
transform 1 0 38180 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_424
timestamp 1649977179
transform 1 0 40112 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_436
timestamp 1649977179
transform 1 0 41216 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1649977179
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1649977179
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1649977179
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1649977179
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1649977179
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1649977179
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1649977179
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1649977179
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1649977179
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1649977179
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1649977179
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1649977179
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1649977179
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1649977179
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1649977179
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1649977179
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_617
timestamp 1649977179
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_37
timestamp 1649977179
transform 1 0 4508 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_45
timestamp 1649977179
transform 1 0 5244 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_62
timestamp 1649977179
transform 1 0 6808 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_68
timestamp 1649977179
transform 1 0 7360 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_80
timestamp 1649977179
transform 1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_91
timestamp 1649977179
transform 1 0 9476 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_100
timestamp 1649977179
transform 1 0 10304 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_110
timestamp 1649977179
transform 1 0 11224 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_122
timestamp 1649977179
transform 1 0 12328 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_130
timestamp 1649977179
transform 1 0 13064 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_135
timestamp 1649977179
transform 1 0 13524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_146
timestamp 1649977179
transform 1 0 14536 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_155
timestamp 1649977179
transform 1 0 15364 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_175
timestamp 1649977179
transform 1 0 17204 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1649977179
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1649977179
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1649977179
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_221
timestamp 1649977179
transform 1 0 21436 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_238
timestamp 1649977179
transform 1 0 23000 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1649977179
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_271
timestamp 1649977179
transform 1 0 26036 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_283
timestamp 1649977179
transform 1 0 27140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_295
timestamp 1649977179
transform 1 0 28244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1649977179
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_315
timestamp 1649977179
transform 1 0 30084 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_323
timestamp 1649977179
transform 1 0 30820 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_340
timestamp 1649977179
transform 1 0 32384 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_352
timestamp 1649977179
transform 1 0 33488 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_395
timestamp 1649977179
transform 1 0 37444 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_401
timestamp 1649977179
transform 1 0 37996 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_404
timestamp 1649977179
transform 1 0 38272 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_412
timestamp 1649977179
transform 1 0 39008 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_416
timestamp 1649977179
transform 1 0 39376 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_421
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_431
timestamp 1649977179
transform 1 0 40756 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_437
timestamp 1649977179
transform 1 0 41308 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_449
timestamp 1649977179
transform 1 0 42412 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_461
timestamp 1649977179
transform 1 0 43516 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_473
timestamp 1649977179
transform 1 0 44620 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1649977179
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1649977179
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1649977179
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1649977179
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1649977179
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1649977179
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1649977179
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1649977179
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1649977179
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1649977179
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1649977179
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1649977179
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1649977179
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_613
timestamp 1649977179
transform 1 0 57500 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_617
timestamp 1649977179
transform 1 0 57868 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_621
timestamp 1649977179
transform 1 0 58236 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_31
timestamp 1649977179
transform 1 0 3956 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_39
timestamp 1649977179
transform 1 0 4692 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1649977179
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_65
timestamp 1649977179
transform 1 0 7084 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_71
timestamp 1649977179
transform 1 0 7636 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_77
timestamp 1649977179
transform 1 0 8188 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_80
timestamp 1649977179
transform 1 0 8464 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_88
timestamp 1649977179
transform 1 0 9200 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_102
timestamp 1649977179
transform 1 0 10488 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1649977179
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_131
timestamp 1649977179
transform 1 0 13156 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_139
timestamp 1649977179
transform 1 0 13892 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_147
timestamp 1649977179
transform 1 0 14628 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_172
timestamp 1649977179
transform 1 0 16928 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_186
timestamp 1649977179
transform 1 0 18216 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_192
timestamp 1649977179
transform 1 0 18768 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_198
timestamp 1649977179
transform 1 0 19320 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_207
timestamp 1649977179
transform 1 0 20148 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1649977179
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_241
timestamp 1649977179
transform 1 0 23276 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_247
timestamp 1649977179
transform 1 0 23828 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_259
timestamp 1649977179
transform 1 0 24932 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_262
timestamp 1649977179
transform 1 0 25208 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_274
timestamp 1649977179
transform 1 0 26312 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_283
timestamp 1649977179
transform 1 0 27140 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_291
timestamp 1649977179
transform 1 0 27876 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_310
timestamp 1649977179
transform 1 0 29624 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_322
timestamp 1649977179
transform 1 0 30728 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_325
timestamp 1649977179
transform 1 0 31004 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_333
timestamp 1649977179
transform 1 0 31740 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_341
timestamp 1649977179
transform 1 0 32476 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_344
timestamp 1649977179
transform 1 0 32752 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_364
timestamp 1649977179
transform 1 0 34592 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_384
timestamp 1649977179
transform 1 0 36432 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_425
timestamp 1649977179
transform 1 0 40204 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_437
timestamp 1649977179
transform 1 0 41308 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_445
timestamp 1649977179
transform 1 0 42044 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1649977179
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1649977179
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1649977179
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1649977179
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1649977179
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1649977179
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1649977179
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1649977179
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1649977179
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1649977179
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1649977179
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1649977179
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1649977179
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1649977179
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1649977179
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_617
timestamp 1649977179
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1649977179
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_37
timestamp 1649977179
transform 1 0 4508 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_43
timestamp 1649977179
transform 1 0 5060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_55
timestamp 1649977179
transform 1 0 6164 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_63
timestamp 1649977179
transform 1 0 6900 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_68
timestamp 1649977179
transform 1 0 7360 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1649977179
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_115
timestamp 1649977179
transform 1 0 11684 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_120
timestamp 1649977179
transform 1 0 12144 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_128
timestamp 1649977179
transform 1 0 12880 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_161
timestamp 1649977179
transform 1 0 15916 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_166
timestamp 1649977179
transform 1 0 16376 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_175
timestamp 1649977179
transform 1 0 17204 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_183
timestamp 1649977179
transform 1 0 17940 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1649977179
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_199
timestamp 1649977179
transform 1 0 19412 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_211
timestamp 1649977179
transform 1 0 20516 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_215
timestamp 1649977179
transform 1 0 20884 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_236
timestamp 1649977179
transform 1 0 22816 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_242
timestamp 1649977179
transform 1 0 23368 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1649977179
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_262
timestamp 1649977179
transform 1 0 25208 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_282
timestamp 1649977179
transform 1 0 27048 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_291
timestamp 1649977179
transform 1 0 27876 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_299
timestamp 1649977179
transform 1 0 28612 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_304
timestamp 1649977179
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_319
timestamp 1649977179
transform 1 0 30452 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_345
timestamp 1649977179
transform 1 0 32844 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1649977179
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1649977179
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_373
timestamp 1649977179
transform 1 0 35420 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_379
timestamp 1649977179
transform 1 0 35972 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_391
timestamp 1649977179
transform 1 0 37076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_403
timestamp 1649977179
transform 1 0 38180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_415
timestamp 1649977179
transform 1 0 39284 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1649977179
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_421
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_428
timestamp 1649977179
transform 1 0 40480 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_437
timestamp 1649977179
transform 1 0 41308 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_449
timestamp 1649977179
transform 1 0 42412 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_461
timestamp 1649977179
transform 1 0 43516 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_473
timestamp 1649977179
transform 1 0 44620 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1649977179
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1649977179
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1649977179
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1649977179
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1649977179
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1649977179
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1649977179
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1649977179
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1649977179
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1649977179
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1649977179
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1649977179
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1649977179
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1649977179
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1649977179
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_23
timestamp 1649977179
transform 1 0 3220 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_30
timestamp 1649977179
transform 1 0 3864 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_42
timestamp 1649977179
transform 1 0 4968 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1649977179
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_61
timestamp 1649977179
transform 1 0 6716 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_78
timestamp 1649977179
transform 1 0 8280 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_84
timestamp 1649977179
transform 1 0 8832 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_90
timestamp 1649977179
transform 1 0 9384 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_104
timestamp 1649977179
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_124
timestamp 1649977179
transform 1 0 12512 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_138
timestamp 1649977179
transform 1 0 13800 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_150
timestamp 1649977179
transform 1 0 14904 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_162
timestamp 1649977179
transform 1 0 16008 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_188
timestamp 1649977179
transform 1 0 18400 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_212
timestamp 1649977179
transform 1 0 20608 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_247
timestamp 1649977179
transform 1 0 23828 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_253
timestamp 1649977179
transform 1 0 24380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_265
timestamp 1649977179
transform 1 0 25484 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_274
timestamp 1649977179
transform 1 0 26312 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_289
timestamp 1649977179
transform 1 0 27692 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_307
timestamp 1649977179
transform 1 0 29348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_315
timestamp 1649977179
transform 1 0 30084 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_318
timestamp 1649977179
transform 1 0 30360 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1649977179
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_341
timestamp 1649977179
transform 1 0 32476 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_360
timestamp 1649977179
transform 1 0 34224 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_369
timestamp 1649977179
transform 1 0 35052 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_381
timestamp 1649977179
transform 1 0 36156 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_389
timestamp 1649977179
transform 1 0 36892 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_425
timestamp 1649977179
transform 1 0 40204 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_437
timestamp 1649977179
transform 1 0 41308 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_445
timestamp 1649977179
transform 1 0 42044 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1649977179
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1649977179
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1649977179
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1649977179
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1649977179
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1649977179
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1649977179
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1649977179
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1649977179
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1649977179
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1649977179
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1649977179
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1649977179
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1649977179
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1649977179
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1649977179
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_617
timestamp 1649977179
transform 1 0 57868 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_621
timestamp 1649977179
transform 1 0 58236 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1649977179
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_49
timestamp 1649977179
transform 1 0 5612 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_57
timestamp 1649977179
transform 1 0 6348 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_68
timestamp 1649977179
transform 1 0 7360 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1649977179
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1649977179
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_91
timestamp 1649977179
transform 1 0 9476 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_99
timestamp 1649977179
transform 1 0 10212 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_110
timestamp 1649977179
transform 1 0 11224 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_116
timestamp 1649977179
transform 1 0 11776 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1649977179
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_165
timestamp 1649977179
transform 1 0 16284 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_170
timestamp 1649977179
transform 1 0 16744 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_176
timestamp 1649977179
transform 1 0 17296 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_182
timestamp 1649977179
transform 1 0 17848 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1649977179
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_211
timestamp 1649977179
transform 1 0 20516 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_219
timestamp 1649977179
transform 1 0 21252 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_228
timestamp 1649977179
transform 1 0 22080 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_240
timestamp 1649977179
transform 1 0 23184 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_255
timestamp 1649977179
transform 1 0 24564 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_267
timestamp 1649977179
transform 1 0 25668 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_291
timestamp 1649977179
transform 1 0 27876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_303
timestamp 1649977179
transform 1 0 28980 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1649977179
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_314
timestamp 1649977179
transform 1 0 29992 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_328
timestamp 1649977179
transform 1 0 31280 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_340
timestamp 1649977179
transform 1 0 32384 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_351
timestamp 1649977179
transform 1 0 33396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1649977179
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1649977179
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1649977179
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1649977179
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1649977179
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1649977179
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1649977179
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1649977179
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1649977179
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1649977179
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1649977179
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1649977179
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1649977179
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1649977179
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1649977179
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1649977179
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1649977179
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1649977179
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1649977179
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1649977179
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1649977179
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1649977179
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1649977179
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1649977179
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1649977179
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_11
timestamp 1649977179
transform 1 0 2116 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_30
timestamp 1649977179
transform 1 0 3864 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_50
timestamp 1649977179
transform 1 0 5704 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_65
timestamp 1649977179
transform 1 0 7084 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_75
timestamp 1649977179
transform 1 0 8004 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_82
timestamp 1649977179
transform 1 0 8648 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_91
timestamp 1649977179
transform 1 0 9476 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_97
timestamp 1649977179
transform 1 0 10028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1649977179
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_118
timestamp 1649977179
transform 1 0 11960 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_131
timestamp 1649977179
transform 1 0 13156 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_140
timestamp 1649977179
transform 1 0 13984 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_160
timestamp 1649977179
transform 1 0 15824 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_177
timestamp 1649977179
transform 1 0 17388 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_185
timestamp 1649977179
transform 1 0 18124 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_196
timestamp 1649977179
transform 1 0 19136 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_210
timestamp 1649977179
transform 1 0 20424 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1649977179
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_233
timestamp 1649977179
transform 1 0 22540 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_245
timestamp 1649977179
transform 1 0 23644 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_253
timestamp 1649977179
transform 1 0 24380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_265
timestamp 1649977179
transform 1 0 25484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_277
timestamp 1649977179
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_305
timestamp 1649977179
transform 1 0 29164 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_309
timestamp 1649977179
transform 1 0 29532 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_318
timestamp 1649977179
transform 1 0 30360 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1649977179
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_339
timestamp 1649977179
transform 1 0 32292 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_355
timestamp 1649977179
transform 1 0 33764 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_366
timestamp 1649977179
transform 1 0 34776 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_376
timestamp 1649977179
transform 1 0 35696 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 1649977179
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_410
timestamp 1649977179
transform 1 0 38824 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_422
timestamp 1649977179
transform 1 0 39928 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_434
timestamp 1649977179
transform 1 0 41032 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_446
timestamp 1649977179
transform 1 0 42136 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1649977179
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1649977179
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1649977179
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1649977179
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1649977179
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1649977179
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1649977179
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1649977179
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1649977179
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1649977179
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1649977179
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1649977179
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1649977179
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1649977179
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1649977179
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1649977179
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1649977179
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1649977179
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_617
timestamp 1649977179
transform 1 0 57868 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_621
timestamp 1649977179
transform 1 0 58236 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_21
timestamp 1649977179
transform 1 0 3036 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_37
timestamp 1649977179
transform 1 0 4508 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_45
timestamp 1649977179
transform 1 0 5244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_57
timestamp 1649977179
transform 1 0 6348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_69
timestamp 1649977179
transform 1 0 7452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_81
timestamp 1649977179
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_104
timestamp 1649977179
transform 1 0 10672 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_116
timestamp 1649977179
transform 1 0 11776 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_124
timestamp 1649977179
transform 1 0 12512 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1649977179
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_143
timestamp 1649977179
transform 1 0 14260 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_155
timestamp 1649977179
transform 1 0 15364 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_163
timestamp 1649977179
transform 1 0 16100 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_173
timestamp 1649977179
transform 1 0 17020 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_179
timestamp 1649977179
transform 1 0 17572 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_187
timestamp 1649977179
transform 1 0 18308 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1649977179
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1649977179
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1649977179
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_233
timestamp 1649977179
transform 1 0 22540 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_241
timestamp 1649977179
transform 1 0 23276 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_244
timestamp 1649977179
transform 1 0 23552 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_257
timestamp 1649977179
transform 1 0 24748 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_263
timestamp 1649977179
transform 1 0 25300 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_271
timestamp 1649977179
transform 1 0 26036 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_274
timestamp 1649977179
transform 1 0 26312 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_282
timestamp 1649977179
transform 1 0 27048 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_294
timestamp 1649977179
transform 1 0 28152 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1649977179
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_312
timestamp 1649977179
transform 1 0 29808 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_326
timestamp 1649977179
transform 1 0 31096 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_332
timestamp 1649977179
transform 1 0 31648 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_344
timestamp 1649977179
transform 1 0 32752 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_356
timestamp 1649977179
transform 1 0 33856 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_48_372
timestamp 1649977179
transform 1 0 35328 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_378
timestamp 1649977179
transform 1 0 35880 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_387
timestamp 1649977179
transform 1 0 36708 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_396
timestamp 1649977179
transform 1 0 37536 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_408
timestamp 1649977179
transform 1 0 38640 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1649977179
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1649977179
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1649977179
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1649977179
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1649977179
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1649977179
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1649977179
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1649977179
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1649977179
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1649977179
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1649977179
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1649977179
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1649977179
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1649977179
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1649977179
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1649977179
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1649977179
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1649977179
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1649977179
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1649977179
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_613
timestamp 1649977179
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_23
timestamp 1649977179
transform 1 0 3220 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_29
timestamp 1649977179
transform 1 0 3772 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_33
timestamp 1649977179
transform 1 0 4140 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_41
timestamp 1649977179
transform 1 0 4876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1649977179
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_69
timestamp 1649977179
transform 1 0 7452 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_75
timestamp 1649977179
transform 1 0 8004 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_81
timestamp 1649977179
transform 1 0 8556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_87
timestamp 1649977179
transform 1 0 9108 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_99
timestamp 1649977179
transform 1 0 10212 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_108
timestamp 1649977179
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_115
timestamp 1649977179
transform 1 0 11684 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_129
timestamp 1649977179
transform 1 0 12972 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_141
timestamp 1649977179
transform 1 0 14076 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_152
timestamp 1649977179
transform 1 0 15088 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_156
timestamp 1649977179
transform 1 0 15456 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_159
timestamp 1649977179
transform 1 0 15732 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1649977179
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_183
timestamp 1649977179
transform 1 0 17940 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_191
timestamp 1649977179
transform 1 0 18676 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_194
timestamp 1649977179
transform 1 0 18952 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_200
timestamp 1649977179
transform 1 0 19504 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_211
timestamp 1649977179
transform 1 0 20516 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1649977179
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1649977179
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_232
timestamp 1649977179
transform 1 0 22448 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_240
timestamp 1649977179
transform 1 0 23184 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_248
timestamp 1649977179
transform 1 0 23920 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_257
timestamp 1649977179
transform 1 0 24748 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_265
timestamp 1649977179
transform 1 0 25484 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1649977179
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1649977179
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_283
timestamp 1649977179
transform 1 0 27140 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_295
timestamp 1649977179
transform 1 0 28244 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_303
timestamp 1649977179
transform 1 0 28980 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_312
timestamp 1649977179
transform 1 0 29808 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_321
timestamp 1649977179
transform 1 0 30636 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_327
timestamp 1649977179
transform 1 0 31188 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1649977179
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_349
timestamp 1649977179
transform 1 0 33212 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_359
timestamp 1649977179
transform 1 0 34132 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_366
timestamp 1649977179
transform 1 0 34776 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_380
timestamp 1649977179
transform 1 0 36064 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_386
timestamp 1649977179
transform 1 0 36616 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_399
timestamp 1649977179
transform 1 0 37812 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_416
timestamp 1649977179
transform 1 0 39376 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_428
timestamp 1649977179
transform 1 0 40480 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_440
timestamp 1649977179
transform 1 0 41584 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1649977179
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1649977179
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1649977179
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1649977179
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1649977179
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1649977179
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1649977179
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1649977179
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1649977179
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1649977179
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1649977179
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1649977179
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1649977179
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1649977179
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1649977179
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1649977179
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1649977179
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1649977179
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_617
timestamp 1649977179
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_15
timestamp 1649977179
transform 1 0 2484 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_21
timestamp 1649977179
transform 1 0 3036 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_42
timestamp 1649977179
transform 1 0 4968 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_54
timestamp 1649977179
transform 1 0 6072 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_66
timestamp 1649977179
transform 1 0 7176 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_78
timestamp 1649977179
transform 1 0 8280 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_103
timestamp 1649977179
transform 1 0 10580 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_112
timestamp 1649977179
transform 1 0 11408 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_118
timestamp 1649977179
transform 1 0 11960 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_130
timestamp 1649977179
transform 1 0 13064 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1649977179
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_153
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_161
timestamp 1649977179
transform 1 0 15916 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_169
timestamp 1649977179
transform 1 0 16652 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_173
timestamp 1649977179
transform 1 0 17020 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_179
timestamp 1649977179
transform 1 0 17572 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_187
timestamp 1649977179
transform 1 0 18308 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1649977179
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_202
timestamp 1649977179
transform 1 0 19688 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_206
timestamp 1649977179
transform 1 0 20056 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_212
timestamp 1649977179
transform 1 0 20608 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_220
timestamp 1649977179
transform 1 0 21344 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_226
timestamp 1649977179
transform 1 0 21896 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_230
timestamp 1649977179
transform 1 0 22264 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_238
timestamp 1649977179
transform 1 0 23000 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1649977179
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_257
timestamp 1649977179
transform 1 0 24748 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_266
timestamp 1649977179
transform 1 0 25576 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_286
timestamp 1649977179
transform 1 0 27416 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_292
timestamp 1649977179
transform 1 0 27968 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1649977179
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_325
timestamp 1649977179
transform 1 0 31004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_333
timestamp 1649977179
transform 1 0 31740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_336
timestamp 1649977179
transform 1 0 32016 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_348
timestamp 1649977179
transform 1 0 33120 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_359
timestamp 1649977179
transform 1 0 34132 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1649977179
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_382
timestamp 1649977179
transform 1 0 36248 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_394
timestamp 1649977179
transform 1 0 37352 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_416
timestamp 1649977179
transform 1 0 39376 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1649977179
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1649977179
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1649977179
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1649977179
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1649977179
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1649977179
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1649977179
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1649977179
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1649977179
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1649977179
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1649977179
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1649977179
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1649977179
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1649977179
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1649977179
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1649977179
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1649977179
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1649977179
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1649977179
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1649977179
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_613
timestamp 1649977179
transform 1 0 57500 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_617
timestamp 1649977179
transform 1 0 57868 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_621
timestamp 1649977179
transform 1 0 58236 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_19
timestamp 1649977179
transform 1 0 2852 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_28
timestamp 1649977179
transform 1 0 3680 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_40
timestamp 1649977179
transform 1 0 4784 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_52
timestamp 1649977179
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_65
timestamp 1649977179
transform 1 0 7084 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_73
timestamp 1649977179
transform 1 0 7820 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_78
timestamp 1649977179
transform 1 0 8280 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_86
timestamp 1649977179
transform 1 0 9016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_95
timestamp 1649977179
transform 1 0 9844 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_104
timestamp 1649977179
transform 1 0 10672 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_119
timestamp 1649977179
transform 1 0 12052 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1649977179
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1649977179
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_149
timestamp 1649977179
transform 1 0 14812 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_159
timestamp 1649977179
transform 1 0 15732 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1649977179
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_174
timestamp 1649977179
transform 1 0 17112 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_180
timestamp 1649977179
transform 1 0 17664 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_192
timestamp 1649977179
transform 1 0 18768 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_204
timestamp 1649977179
transform 1 0 19872 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1649977179
transform 1 0 21344 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_244
timestamp 1649977179
transform 1 0 23552 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_255
timestamp 1649977179
transform 1 0 24564 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_269
timestamp 1649977179
transform 1 0 25852 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_275
timestamp 1649977179
transform 1 0 26404 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1649977179
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_293
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_301
timestamp 1649977179
transform 1 0 28796 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_307
timestamp 1649977179
transform 1 0 29348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_319
timestamp 1649977179
transform 1 0 30452 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1649977179
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1649977179
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_341
timestamp 1649977179
transform 1 0 32476 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_358
timestamp 1649977179
transform 1 0 34040 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_366
timestamp 1649977179
transform 1 0 34776 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_374
timestamp 1649977179
transform 1 0 35512 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_386
timestamp 1649977179
transform 1 0 36616 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_395
timestamp 1649977179
transform 1 0 37444 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_407
timestamp 1649977179
transform 1 0 38548 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_419
timestamp 1649977179
transform 1 0 39652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_431
timestamp 1649977179
transform 1 0 40756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_443
timestamp 1649977179
transform 1 0 41860 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1649977179
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1649977179
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1649977179
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1649977179
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1649977179
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1649977179
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1649977179
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1649977179
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1649977179
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1649977179
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1649977179
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1649977179
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1649977179
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1649977179
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1649977179
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1649977179
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1649977179
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1649977179
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1649977179
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1649977179
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_7
timestamp 1649977179
transform 1 0 1748 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_24
timestamp 1649977179
transform 1 0 3312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_73
timestamp 1649977179
transform 1 0 7820 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_79
timestamp 1649977179
transform 1 0 8372 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_93
timestamp 1649977179
transform 1 0 9660 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1649977179
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1649977179
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_121
timestamp 1649977179
transform 1 0 12236 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_134
timestamp 1649977179
transform 1 0 13432 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_148
timestamp 1649977179
transform 1 0 14720 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_168
timestamp 1649977179
transform 1 0 16560 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1649977179
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_199
timestamp 1649977179
transform 1 0 19412 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_207
timestamp 1649977179
transform 1 0 20148 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_210
timestamp 1649977179
transform 1 0 20424 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_222
timestamp 1649977179
transform 1 0 21528 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_226
timestamp 1649977179
transform 1 0 21896 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_238
timestamp 1649977179
transform 1 0 23000 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 1649977179
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_259
timestamp 1649977179
transform 1 0 24932 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_263
timestamp 1649977179
transform 1 0 25300 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_280
timestamp 1649977179
transform 1 0 26864 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1649977179
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_311
timestamp 1649977179
transform 1 0 29716 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_325
timestamp 1649977179
transform 1 0 31004 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_329
timestamp 1649977179
transform 1 0 31372 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_332
timestamp 1649977179
transform 1 0 31648 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_344
timestamp 1649977179
transform 1 0 32752 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_348
timestamp 1649977179
transform 1 0 33120 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_356
timestamp 1649977179
transform 1 0 33856 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_369
timestamp 1649977179
transform 1 0 35052 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_375
timestamp 1649977179
transform 1 0 35604 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_387
timestamp 1649977179
transform 1 0 36708 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_393
timestamp 1649977179
transform 1 0 37260 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_399
timestamp 1649977179
transform 1 0 37812 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_416
timestamp 1649977179
transform 1 0 39376 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1649977179
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1649977179
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1649977179
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1649977179
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1649977179
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1649977179
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1649977179
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1649977179
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1649977179
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1649977179
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1649977179
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1649977179
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1649977179
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1649977179
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1649977179
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1649977179
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1649977179
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1649977179
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1649977179
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1649977179
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_613
timestamp 1649977179
transform 1 0 57500 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_617
timestamp 1649977179
transform 1 0 57868 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_621
timestamp 1649977179
transform 1 0 58236 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_11
timestamp 1649977179
transform 1 0 2116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_19
timestamp 1649977179
transform 1 0 2852 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_25
timestamp 1649977179
transform 1 0 3404 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_37
timestamp 1649977179
transform 1 0 4508 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_45
timestamp 1649977179
transform 1 0 5244 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_52
timestamp 1649977179
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_65
timestamp 1649977179
transform 1 0 7084 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_93
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_99
timestamp 1649977179
transform 1 0 10212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1649977179
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_149
timestamp 1649977179
transform 1 0 14812 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_158
timestamp 1649977179
transform 1 0 15640 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1649977179
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_171
timestamp 1649977179
transform 1 0 16836 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_177
timestamp 1649977179
transform 1 0 17388 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_188
timestamp 1649977179
transform 1 0 18400 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_196
timestamp 1649977179
transform 1 0 19136 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_215
timestamp 1649977179
transform 1 0 20884 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1649977179
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_231
timestamp 1649977179
transform 1 0 22356 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_237
timestamp 1649977179
transform 1 0 22908 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_243
timestamp 1649977179
transform 1 0 23460 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_251
timestamp 1649977179
transform 1 0 24196 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_257
timestamp 1649977179
transform 1 0 24748 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_265
timestamp 1649977179
transform 1 0 25484 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1649977179
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1649977179
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_295
timestamp 1649977179
transform 1 0 28244 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_319
timestamp 1649977179
transform 1 0 30452 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_330
timestamp 1649977179
transform 1 0 31464 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_342
timestamp 1649977179
transform 1 0 32568 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_351
timestamp 1649977179
transform 1 0 33396 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_363
timestamp 1649977179
transform 1 0 34500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_375
timestamp 1649977179
transform 1 0 35604 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_382
timestamp 1649977179
transform 1 0 36248 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_390
timestamp 1649977179
transform 1 0 36984 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_393
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1649977179
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1649977179
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1649977179
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1649977179
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1649977179
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1649977179
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1649977179
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1649977179
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1649977179
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1649977179
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1649977179
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1649977179
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1649977179
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1649977179
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1649977179
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1649977179
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1649977179
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1649977179
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1649977179
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1649977179
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1649977179
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1649977179
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_617
timestamp 1649977179
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_19
timestamp 1649977179
transform 1 0 2852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1649977179
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_37
timestamp 1649977179
transform 1 0 4508 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_48
timestamp 1649977179
transform 1 0 5520 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_72
timestamp 1649977179
transform 1 0 7728 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_78
timestamp 1649977179
transform 1 0 8280 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_107
timestamp 1649977179
transform 1 0 10948 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_119
timestamp 1649977179
transform 1 0 12052 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_127
timestamp 1649977179
transform 1 0 12788 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_134
timestamp 1649977179
transform 1 0 13432 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_149
timestamp 1649977179
transform 1 0 14812 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_155
timestamp 1649977179
transform 1 0 15364 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_161
timestamp 1649977179
transform 1 0 15916 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_166
timestamp 1649977179
transform 1 0 16376 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_190
timestamp 1649977179
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1649977179
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_223
timestamp 1649977179
transform 1 0 21620 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_237
timestamp 1649977179
transform 1 0 22908 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_249
timestamp 1649977179
transform 1 0 24012 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_253
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_267
timestamp 1649977179
transform 1 0 25668 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_273
timestamp 1649977179
transform 1 0 26220 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_285
timestamp 1649977179
transform 1 0 27324 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_300
timestamp 1649977179
transform 1 0 28704 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_325
timestamp 1649977179
transform 1 0 31004 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_333
timestamp 1649977179
transform 1 0 31740 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_338
timestamp 1649977179
transform 1 0 32200 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_344
timestamp 1649977179
transform 1 0 32752 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_356
timestamp 1649977179
transform 1 0 33856 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_375
timestamp 1649977179
transform 1 0 35604 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_387
timestamp 1649977179
transform 1 0 36708 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_397
timestamp 1649977179
transform 1 0 37628 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_409
timestamp 1649977179
transform 1 0 38732 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_417
timestamp 1649977179
transform 1 0 39468 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1649977179
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1649977179
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1649977179
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1649977179
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1649977179
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1649977179
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1649977179
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1649977179
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1649977179
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1649977179
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1649977179
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1649977179
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1649977179
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1649977179
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1649977179
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1649977179
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1649977179
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1649977179
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1649977179
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1649977179
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1649977179
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_11
timestamp 1649977179
transform 1 0 2116 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_28
timestamp 1649977179
transform 1 0 3680 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_40
timestamp 1649977179
transform 1 0 4784 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_45
timestamp 1649977179
transform 1 0 5244 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1649977179
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_65
timestamp 1649977179
transform 1 0 7084 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_71
timestamp 1649977179
transform 1 0 7636 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_82
timestamp 1649977179
transform 1 0 8648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_96
timestamp 1649977179
transform 1 0 9936 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_108
timestamp 1649977179
transform 1 0 11040 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_115
timestamp 1649977179
transform 1 0 11684 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_127
timestamp 1649977179
transform 1 0 12788 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_141
timestamp 1649977179
transform 1 0 14076 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_153
timestamp 1649977179
transform 1 0 15180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_165
timestamp 1649977179
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_177
timestamp 1649977179
transform 1 0 17388 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_187
timestamp 1649977179
transform 1 0 18308 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_207
timestamp 1649977179
transform 1 0 20148 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_219
timestamp 1649977179
transform 1 0 21252 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1649977179
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_233
timestamp 1649977179
transform 1 0 22540 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_245
timestamp 1649977179
transform 1 0 23644 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_251
timestamp 1649977179
transform 1 0 24196 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_255
timestamp 1649977179
transform 1 0 24564 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_265
timestamp 1649977179
transform 1 0 25484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_277
timestamp 1649977179
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_293
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_301
timestamp 1649977179
transform 1 0 28796 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_313
timestamp 1649977179
transform 1 0 29900 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_317
timestamp 1649977179
transform 1 0 30268 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_321
timestamp 1649977179
transform 1 0 30636 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_333
timestamp 1649977179
transform 1 0 31740 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_346
timestamp 1649977179
transform 1 0 32936 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_358
timestamp 1649977179
transform 1 0 34040 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_370
timestamp 1649977179
transform 1 0 35144 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_382
timestamp 1649977179
transform 1 0 36248 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_390
timestamp 1649977179
transform 1 0 36984 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_409
timestamp 1649977179
transform 1 0 38732 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_421
timestamp 1649977179
transform 1 0 39836 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_433
timestamp 1649977179
transform 1 0 40940 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_445
timestamp 1649977179
transform 1 0 42044 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1649977179
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1649977179
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1649977179
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1649977179
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1649977179
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1649977179
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1649977179
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1649977179
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1649977179
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1649977179
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1649977179
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1649977179
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1649977179
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1649977179
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1649977179
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1649977179
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1649977179
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1649977179
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_617
timestamp 1649977179
transform 1 0 57868 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_621
timestamp 1649977179
transform 1 0 58236 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_47
timestamp 1649977179
transform 1 0 5428 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_50
timestamp 1649977179
transform 1 0 5704 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_54
timestamp 1649977179
transform 1 0 6072 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_57
timestamp 1649977179
transform 1 0 6348 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_69
timestamp 1649977179
transform 1 0 7452 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_78
timestamp 1649977179
transform 1 0 8280 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_89
timestamp 1649977179
transform 1 0 9292 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_94
timestamp 1649977179
transform 1 0 9752 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_103
timestamp 1649977179
transform 1 0 10580 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_107
timestamp 1649977179
transform 1 0 10948 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_110
timestamp 1649977179
transform 1 0 11224 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_122
timestamp 1649977179
transform 1 0 12328 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_130
timestamp 1649977179
transform 1 0 13064 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_136
timestamp 1649977179
transform 1 0 13616 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_151
timestamp 1649977179
transform 1 0 14996 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_157
timestamp 1649977179
transform 1 0 15548 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_163
timestamp 1649977179
transform 1 0 16100 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_172
timestamp 1649977179
transform 1 0 16928 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_182
timestamp 1649977179
transform 1 0 17848 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_191
timestamp 1649977179
transform 1 0 18676 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1649977179
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1649977179
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_221
timestamp 1649977179
transform 1 0 21436 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_229
timestamp 1649977179
transform 1 0 22172 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_241
timestamp 1649977179
transform 1 0 23276 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1649977179
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_263
timestamp 1649977179
transform 1 0 25300 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_267
timestamp 1649977179
transform 1 0 25668 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_284
timestamp 1649977179
transform 1 0 27232 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_290
timestamp 1649977179
transform 1 0 27784 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_302
timestamp 1649977179
transform 1 0 28888 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_313
timestamp 1649977179
transform 1 0 29900 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_321
timestamp 1649977179
transform 1 0 30636 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_329
timestamp 1649977179
transform 1 0 31372 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_335
timestamp 1649977179
transform 1 0 31924 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_349
timestamp 1649977179
transform 1 0 33212 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_361
timestamp 1649977179
transform 1 0 34316 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_381
timestamp 1649977179
transform 1 0 36156 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_393
timestamp 1649977179
transform 1 0 37260 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_405
timestamp 1649977179
transform 1 0 38364 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_417
timestamp 1649977179
transform 1 0 39468 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1649977179
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1649977179
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1649977179
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1649977179
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1649977179
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1649977179
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1649977179
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1649977179
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1649977179
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1649977179
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1649977179
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1649977179
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1649977179
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1649977179
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1649977179
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1649977179
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1649977179
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1649977179
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1649977179
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1649977179
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1649977179
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_32
timestamp 1649977179
transform 1 0 4048 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_41
timestamp 1649977179
transform 1 0 4876 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_47
timestamp 1649977179
transform 1 0 5428 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_76
timestamp 1649977179
transform 1 0 8096 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_88
timestamp 1649977179
transform 1 0 9200 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_100
timestamp 1649977179
transform 1 0 10304 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_115
timestamp 1649977179
transform 1 0 11684 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_145
timestamp 1649977179
transform 1 0 14444 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_157
timestamp 1649977179
transform 1 0 15548 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_165
timestamp 1649977179
transform 1 0 16284 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_57_174
timestamp 1649977179
transform 1 0 17112 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_180
timestamp 1649977179
transform 1 0 17664 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_183
timestamp 1649977179
transform 1 0 17940 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_191
timestamp 1649977179
transform 1 0 18676 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_195
timestamp 1649977179
transform 1 0 19044 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_200
timestamp 1649977179
transform 1 0 19504 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_206
timestamp 1649977179
transform 1 0 20056 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_218
timestamp 1649977179
transform 1 0 21160 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_57_241
timestamp 1649977179
transform 1 0 23276 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_247
timestamp 1649977179
transform 1 0 23828 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_256
timestamp 1649977179
transform 1 0 24656 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_268
timestamp 1649977179
transform 1 0 25760 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_276
timestamp 1649977179
transform 1 0 26496 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_292
timestamp 1649977179
transform 1 0 27968 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_304
timestamp 1649977179
transform 1 0 29072 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_308
timestamp 1649977179
transform 1 0 29440 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_311
timestamp 1649977179
transform 1 0 29716 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_323
timestamp 1649977179
transform 1 0 30820 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_331
timestamp 1649977179
transform 1 0 31556 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1649977179
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_359
timestamp 1649977179
transform 1 0 34132 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_379
timestamp 1649977179
transform 1 0 35972 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1649977179
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1649977179
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1649977179
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1649977179
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1649977179
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1649977179
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1649977179
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1649977179
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1649977179
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1649977179
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1649977179
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1649977179
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1649977179
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1649977179
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1649977179
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1649977179
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1649977179
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1649977179
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1649977179
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1649977179
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1649977179
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1649977179
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1649977179
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_617
timestamp 1649977179
transform 1 0 57868 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_621
timestamp 1649977179
transform 1 0 58236 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1649977179
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1649977179
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_37
timestamp 1649977179
transform 1 0 4508 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_46
timestamp 1649977179
transform 1 0 5336 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_52
timestamp 1649977179
transform 1 0 5888 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_64
timestamp 1649977179
transform 1 0 6992 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_68
timestamp 1649977179
transform 1 0 7360 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_71
timestamp 1649977179
transform 1 0 7636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_97
timestamp 1649977179
transform 1 0 10028 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_109
timestamp 1649977179
transform 1 0 11132 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_115
timestamp 1649977179
transform 1 0 11684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_127
timestamp 1649977179
transform 1 0 12788 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_131
timestamp 1649977179
transform 1 0 13156 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 1649977179
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_149
timestamp 1649977179
transform 1 0 14812 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_155
timestamp 1649977179
transform 1 0 15364 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_172
timestamp 1649977179
transform 1 0 16928 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_184
timestamp 1649977179
transform 1 0 18032 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_190
timestamp 1649977179
transform 1 0 18584 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_206
timestamp 1649977179
transform 1 0 20056 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_218
timestamp 1649977179
transform 1 0 21160 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_226
timestamp 1649977179
transform 1 0 21896 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_246
timestamp 1649977179
transform 1 0 23736 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_257
timestamp 1649977179
transform 1 0 24748 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_263
timestamp 1649977179
transform 1 0 25300 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_267
timestamp 1649977179
transform 1 0 25668 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_270
timestamp 1649977179
transform 1 0 25944 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_278
timestamp 1649977179
transform 1 0 26680 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_297
timestamp 1649977179
transform 1 0 28428 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_301
timestamp 1649977179
transform 1 0 28796 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_304
timestamp 1649977179
transform 1 0 29072 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_323
timestamp 1649977179
transform 1 0 30820 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_332
timestamp 1649977179
transform 1 0 31648 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_340
timestamp 1649977179
transform 1 0 32384 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_348
timestamp 1649977179
transform 1 0 33120 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 1649977179
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_370
timestamp 1649977179
transform 1 0 35144 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_382
timestamp 1649977179
transform 1 0 36248 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_394
timestamp 1649977179
transform 1 0 37352 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_406
timestamp 1649977179
transform 1 0 38456 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_418
timestamp 1649977179
transform 1 0 39560 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1649977179
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1649977179
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1649977179
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1649977179
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1649977179
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1649977179
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1649977179
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1649977179
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1649977179
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1649977179
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1649977179
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1649977179
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1649977179
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1649977179
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1649977179
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1649977179
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1649977179
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1649977179
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1649977179
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1649977179
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1649977179
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_15
timestamp 1649977179
transform 1 0 2484 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_32
timestamp 1649977179
transform 1 0 4048 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_44
timestamp 1649977179
transform 1 0 5152 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_50
timestamp 1649977179
transform 1 0 5704 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_75
timestamp 1649977179
transform 1 0 8004 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_87
timestamp 1649977179
transform 1 0 9108 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_95
timestamp 1649977179
transform 1 0 9844 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_99
timestamp 1649977179
transform 1 0 10212 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_108
timestamp 1649977179
transform 1 0 11040 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_118
timestamp 1649977179
transform 1 0 11960 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_124
timestamp 1649977179
transform 1 0 12512 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1649977179
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_161
timestamp 1649977179
transform 1 0 15916 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1649977179
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_169
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_173
timestamp 1649977179
transform 1 0 17020 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_182
timestamp 1649977179
transform 1 0 17848 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_190
timestamp 1649977179
transform 1 0 18584 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_197
timestamp 1649977179
transform 1 0 19228 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_209
timestamp 1649977179
transform 1 0 20332 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_215
timestamp 1649977179
transform 1 0 20884 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1649977179
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1649977179
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_249
timestamp 1649977179
transform 1 0 24012 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_255
timestamp 1649977179
transform 1 0 24564 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_258
timestamp 1649977179
transform 1 0 24840 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_270
timestamp 1649977179
transform 1 0 25944 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_278
timestamp 1649977179
transform 1 0 26680 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_294
timestamp 1649977179
transform 1 0 28152 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_300
timestamp 1649977179
transform 1 0 28704 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_312
timestamp 1649977179
transform 1 0 29808 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_332
timestamp 1649977179
transform 1 0 31648 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_351
timestamp 1649977179
transform 1 0 33396 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_363
timestamp 1649977179
transform 1 0 34500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_375
timestamp 1649977179
transform 1 0 35604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_387
timestamp 1649977179
transform 1 0 36708 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1649977179
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1649977179
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1649977179
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1649977179
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1649977179
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1649977179
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1649977179
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1649977179
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1649977179
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1649977179
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1649977179
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1649977179
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1649977179
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1649977179
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1649977179
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1649977179
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1649977179
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1649977179
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1649977179
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1649977179
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1649977179
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1649977179
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1649977179
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1649977179
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_617
timestamp 1649977179
transform 1 0 57868 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_33
timestamp 1649977179
transform 1 0 4140 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_42
timestamp 1649977179
transform 1 0 4968 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_48
timestamp 1649977179
transform 1 0 5520 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_56
timestamp 1649977179
transform 1 0 6256 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_62
timestamp 1649977179
transform 1 0 6808 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_74
timestamp 1649977179
transform 1 0 7912 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_80
timestamp 1649977179
transform 1 0 8464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_99
timestamp 1649977179
transform 1 0 10212 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_119
timestamp 1649977179
transform 1 0 12052 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_127
timestamp 1649977179
transform 1 0 12788 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_136
timestamp 1649977179
transform 1 0 13616 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_173
timestamp 1649977179
transform 1 0 17020 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_190
timestamp 1649977179
transform 1 0 18584 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_201
timestamp 1649977179
transform 1 0 19596 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_207
timestamp 1649977179
transform 1 0 20148 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_224
timestamp 1649977179
transform 1 0 21712 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_230
timestamp 1649977179
transform 1 0 22264 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_242
timestamp 1649977179
transform 1 0 23368 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1649977179
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_261
timestamp 1649977179
transform 1 0 25116 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_267
timestamp 1649977179
transform 1 0 25668 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_279
timestamp 1649977179
transform 1 0 26772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_291
timestamp 1649977179
transform 1 0 27876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_303
timestamp 1649977179
transform 1 0 28980 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_320
timestamp 1649977179
transform 1 0 30544 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_334
timestamp 1649977179
transform 1 0 31832 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_346
timestamp 1649977179
transform 1 0 32936 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_352
timestamp 1649977179
transform 1 0 33488 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_355
timestamp 1649977179
transform 1 0 33764 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1649977179
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1649977179
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1649977179
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1649977179
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1649977179
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1649977179
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1649977179
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1649977179
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1649977179
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1649977179
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1649977179
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1649977179
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1649977179
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1649977179
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1649977179
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1649977179
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1649977179
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1649977179
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1649977179
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1649977179
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1649977179
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1649977179
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1649977179
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1649977179
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1649977179
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_613
timestamp 1649977179
transform 1 0 57500 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_617
timestamp 1649977179
transform 1 0 57868 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_621
timestamp 1649977179
transform 1 0 58236 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_27
timestamp 1649977179
transform 1 0 3588 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_40
timestamp 1649977179
transform 1 0 4784 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_46
timestamp 1649977179
transform 1 0 5336 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1649977179
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_73
timestamp 1649977179
transform 1 0 7820 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_79
timestamp 1649977179
transform 1 0 8372 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_90
timestamp 1649977179
transform 1 0 9384 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_104
timestamp 1649977179
transform 1 0 10672 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_118
timestamp 1649977179
transform 1 0 11960 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_124
timestamp 1649977179
transform 1 0 12512 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_127
timestamp 1649977179
transform 1 0 12788 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_135
timestamp 1649977179
transform 1 0 13524 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_141
timestamp 1649977179
transform 1 0 14076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_153
timestamp 1649977179
transform 1 0 15180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_165
timestamp 1649977179
transform 1 0 16284 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_182
timestamp 1649977179
transform 1 0 17848 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_194
timestamp 1649977179
transform 1 0 18952 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_206
timestamp 1649977179
transform 1 0 20056 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_218
timestamp 1649977179
transform 1 0 21160 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_233
timestamp 1649977179
transform 1 0 22540 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_239
timestamp 1649977179
transform 1 0 23092 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_248
timestamp 1649977179
transform 1 0 23920 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_262
timestamp 1649977179
transform 1 0 25208 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_268
timestamp 1649977179
transform 1 0 25760 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_285
timestamp 1649977179
transform 1 0 27324 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_297
timestamp 1649977179
transform 1 0 28428 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_309
timestamp 1649977179
transform 1 0 29532 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_321
timestamp 1649977179
transform 1 0 30636 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_333
timestamp 1649977179
transform 1 0 31740 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_61_337
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_341
timestamp 1649977179
transform 1 0 32476 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_349
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_355
timestamp 1649977179
transform 1 0 33764 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1649977179
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1649977179
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1649977179
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1649977179
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1649977179
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1649977179
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1649977179
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1649977179
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1649977179
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1649977179
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1649977179
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1649977179
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1649977179
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1649977179
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1649977179
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1649977179
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1649977179
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1649977179
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1649977179
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1649977179
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1649977179
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1649977179
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1649977179
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1649977179
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1649977179
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1649977179
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1649977179
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_617
timestamp 1649977179
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1649977179
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_45
timestamp 1649977179
transform 1 0 5244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_57
timestamp 1649977179
transform 1 0 6348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_60
timestamp 1649977179
transform 1 0 6624 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_72
timestamp 1649977179
transform 1 0 7728 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_94
timestamp 1649977179
transform 1 0 9752 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_114
timestamp 1649977179
transform 1 0 11592 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_122
timestamp 1649977179
transform 1 0 12328 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_127
timestamp 1649977179
transform 1 0 12788 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_131
timestamp 1649977179
transform 1 0 13156 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_136
timestamp 1649977179
transform 1 0 13616 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_149
timestamp 1649977179
transform 1 0 14812 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_155
timestamp 1649977179
transform 1 0 15364 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_163
timestamp 1649977179
transform 1 0 16100 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_166
timestamp 1649977179
transform 1 0 16376 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_178
timestamp 1649977179
transform 1 0 17480 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_190
timestamp 1649977179
transform 1 0 18584 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_221
timestamp 1649977179
transform 1 0 21436 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_227
timestamp 1649977179
transform 1 0 21988 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_235
timestamp 1649977179
transform 1 0 22724 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_248
timestamp 1649977179
transform 1 0 23920 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_255
timestamp 1649977179
transform 1 0 24564 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_277
timestamp 1649977179
transform 1 0 26588 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_283
timestamp 1649977179
transform 1 0 27140 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_295
timestamp 1649977179
transform 1 0 28244 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_304
timestamp 1649977179
transform 1 0 29072 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_314
timestamp 1649977179
transform 1 0 29992 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_320
timestamp 1649977179
transform 1 0 30544 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_328
timestamp 1649977179
transform 1 0 31280 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_331
timestamp 1649977179
transform 1 0 31556 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_345
timestamp 1649977179
transform 1 0 32844 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_351
timestamp 1649977179
transform 1 0 33396 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_360
timestamp 1649977179
transform 1 0 34224 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_370
timestamp 1649977179
transform 1 0 35144 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_374
timestamp 1649977179
transform 1 0 35512 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_391
timestamp 1649977179
transform 1 0 37076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_403
timestamp 1649977179
transform 1 0 38180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_415
timestamp 1649977179
transform 1 0 39284 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1649977179
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1649977179
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1649977179
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1649977179
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1649977179
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1649977179
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1649977179
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1649977179
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1649977179
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1649977179
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1649977179
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1649977179
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1649977179
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1649977179
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1649977179
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1649977179
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1649977179
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1649977179
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1649977179
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1649977179
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1649977179
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_613
timestamp 1649977179
transform 1 0 57500 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_617
timestamp 1649977179
transform 1 0 57868 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_621
timestamp 1649977179
transform 1 0 58236 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_21
timestamp 1649977179
transform 1 0 3036 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_42
timestamp 1649977179
transform 1 0 4968 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_48
timestamp 1649977179
transform 1 0 5520 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_57
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_66
timestamp 1649977179
transform 1 0 7176 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_75
timestamp 1649977179
transform 1 0 8004 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_87
timestamp 1649977179
transform 1 0 9108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_99
timestamp 1649977179
transform 1 0 10212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1649977179
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_117
timestamp 1649977179
transform 1 0 11868 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_122
timestamp 1649977179
transform 1 0 12328 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_130
timestamp 1649977179
transform 1 0 13064 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_147
timestamp 1649977179
transform 1 0 14628 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_155
timestamp 1649977179
transform 1 0 15364 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_164
timestamp 1649977179
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_174
timestamp 1649977179
transform 1 0 17112 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_180
timestamp 1649977179
transform 1 0 17664 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_186
timestamp 1649977179
transform 1 0 18216 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_192
timestamp 1649977179
transform 1 0 18768 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_196
timestamp 1649977179
transform 1 0 19136 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_199
timestamp 1649977179
transform 1 0 19412 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_211
timestamp 1649977179
transform 1 0 20516 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1649977179
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1649977179
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_230
timestamp 1649977179
transform 1 0 22264 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_241
timestamp 1649977179
transform 1 0 23276 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_265
timestamp 1649977179
transform 1 0 25484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_271
timestamp 1649977179
transform 1 0 26036 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1649977179
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_281
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_285
timestamp 1649977179
transform 1 0 27324 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_302
timestamp 1649977179
transform 1 0 28888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_314
timestamp 1649977179
transform 1 0 29992 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_330
timestamp 1649977179
transform 1 0 31464 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_341
timestamp 1649977179
transform 1 0 32476 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_350
timestamp 1649977179
transform 1 0 33304 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_354
timestamp 1649977179
transform 1 0 33672 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_363
timestamp 1649977179
transform 1 0 34500 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_383
timestamp 1649977179
transform 1 0 36340 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1649977179
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1649977179
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1649977179
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1649977179
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1649977179
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1649977179
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1649977179
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1649977179
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1649977179
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1649977179
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1649977179
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1649977179
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1649977179
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1649977179
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1649977179
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1649977179
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1649977179
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1649977179
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1649977179
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1649977179
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1649977179
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1649977179
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1649977179
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1649977179
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1649977179
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_617
timestamp 1649977179
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_7
timestamp 1649977179
transform 1 0 1748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_24
timestamp 1649977179
transform 1 0 3312 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_41
timestamp 1649977179
transform 1 0 4876 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_65
timestamp 1649977179
transform 1 0 7084 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_76
timestamp 1649977179
transform 1 0 8096 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1649977179
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1649977179
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1649977179
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1649977179
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_146
timestamp 1649977179
transform 1 0 14536 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_154
timestamp 1649977179
transform 1 0 15272 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_171
timestamp 1649977179
transform 1 0 16836 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_187
timestamp 1649977179
transform 1 0 18308 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1649977179
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_206
timestamp 1649977179
transform 1 0 20056 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_226
timestamp 1649977179
transform 1 0 21896 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_232
timestamp 1649977179
transform 1 0 22448 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_243
timestamp 1649977179
transform 1 0 23460 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1649977179
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_255
timestamp 1649977179
transform 1 0 24564 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_275
timestamp 1649977179
transform 1 0 26404 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_287
timestamp 1649977179
transform 1 0 27508 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_299
timestamp 1649977179
transform 1 0 28612 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1649977179
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_311
timestamp 1649977179
transform 1 0 29716 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_319
timestamp 1649977179
transform 1 0 30452 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_336
timestamp 1649977179
transform 1 0 32016 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1649977179
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_373
timestamp 1649977179
transform 1 0 35420 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_385
timestamp 1649977179
transform 1 0 36524 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_397
timestamp 1649977179
transform 1 0 37628 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_409
timestamp 1649977179
transform 1 0 38732 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_417
timestamp 1649977179
transform 1 0 39468 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1649977179
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1649977179
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1649977179
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1649977179
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1649977179
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1649977179
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1649977179
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1649977179
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1649977179
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1649977179
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1649977179
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1649977179
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1649977179
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1649977179
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1649977179
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1649977179
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1649977179
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1649977179
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1649977179
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1649977179
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_613
timestamp 1649977179
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1649977179
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_15
timestamp 1649977179
transform 1 0 2484 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_26
timestamp 1649977179
transform 1 0 3496 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_32
timestamp 1649977179
transform 1 0 4048 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_44
timestamp 1649977179
transform 1 0 5152 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1649977179
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_69
timestamp 1649977179
transform 1 0 7452 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_77
timestamp 1649977179
transform 1 0 8188 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_81
timestamp 1649977179
transform 1 0 8556 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_65_89
timestamp 1649977179
transform 1 0 9292 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_97
timestamp 1649977179
transform 1 0 10028 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_104
timestamp 1649977179
transform 1 0 10672 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_120
timestamp 1649977179
transform 1 0 12144 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_132
timestamp 1649977179
transform 1 0 13248 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_144
timestamp 1649977179
transform 1 0 14352 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_156
timestamp 1649977179
transform 1 0 15456 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_169
timestamp 1649977179
transform 1 0 16652 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_175
timestamp 1649977179
transform 1 0 17204 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_184
timestamp 1649977179
transform 1 0 18032 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_204
timestamp 1649977179
transform 1 0 19872 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_213
timestamp 1649977179
transform 1 0 20700 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_221
timestamp 1649977179
transform 1 0 21436 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1649977179
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_237
timestamp 1649977179
transform 1 0 22908 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_243
timestamp 1649977179
transform 1 0 23460 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_249
timestamp 1649977179
transform 1 0 24012 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_261
timestamp 1649977179
transform 1 0 25116 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_270
timestamp 1649977179
transform 1 0 25944 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_278
timestamp 1649977179
transform 1 0 26680 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_281
timestamp 1649977179
transform 1 0 26956 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_289
timestamp 1649977179
transform 1 0 27692 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_310
timestamp 1649977179
transform 1 0 29624 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_316
timestamp 1649977179
transform 1 0 30176 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_325
timestamp 1649977179
transform 1 0 31004 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_331
timestamp 1649977179
transform 1 0 31556 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1649977179
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_337
timestamp 1649977179
transform 1 0 32108 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_355
timestamp 1649977179
transform 1 0 33764 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_365
timestamp 1649977179
transform 1 0 34684 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_377
timestamp 1649977179
transform 1 0 35788 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_389
timestamp 1649977179
transform 1 0 36892 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1649977179
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1649977179
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1649977179
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1649977179
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1649977179
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1649977179
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1649977179
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1649977179
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1649977179
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1649977179
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1649977179
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1649977179
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1649977179
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1649977179
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1649977179
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1649977179
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1649977179
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1649977179
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1649977179
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1649977179
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1649977179
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1649977179
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1649977179
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1649977179
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_617
timestamp 1649977179
transform 1 0 57868 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_621
timestamp 1649977179
transform 1 0 58236 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1649977179
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_15
timestamp 1649977179
transform 1 0 2484 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_24
timestamp 1649977179
transform 1 0 3312 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_34
timestamp 1649977179
transform 1 0 4232 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_46
timestamp 1649977179
transform 1 0 5336 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_62
timestamp 1649977179
transform 1 0 6808 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_68
timestamp 1649977179
transform 1 0 7360 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_80
timestamp 1649977179
transform 1 0 8464 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_85
timestamp 1649977179
transform 1 0 8924 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1649977179
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1649977179
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1649977179
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1649977179
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1649977179
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_153
timestamp 1649977179
transform 1 0 15180 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_166
timestamp 1649977179
transform 1 0 16376 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1649977179
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1649977179
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1649977179
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_197
timestamp 1649977179
transform 1 0 19228 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_206
timestamp 1649977179
transform 1 0 20056 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_218
timestamp 1649977179
transform 1 0 21160 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_230
timestamp 1649977179
transform 1 0 22264 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_242
timestamp 1649977179
transform 1 0 23368 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_250
timestamp 1649977179
transform 1 0 24104 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_253
timestamp 1649977179
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_271
timestamp 1649977179
transform 1 0 26036 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_283
timestamp 1649977179
transform 1 0 27140 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_291
timestamp 1649977179
transform 1 0 27876 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_298
timestamp 1649977179
transform 1 0 28520 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_306
timestamp 1649977179
transform 1 0 29256 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_325
timestamp 1649977179
transform 1 0 31004 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_334
timestamp 1649977179
transform 1 0 31832 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_340
timestamp 1649977179
transform 1 0 32384 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_352
timestamp 1649977179
transform 1 0 33488 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1649977179
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1649977179
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1649977179
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1649977179
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1649977179
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1649977179
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1649977179
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1649977179
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1649977179
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1649977179
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1649977179
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1649977179
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1649977179
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1649977179
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1649977179
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1649977179
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1649977179
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1649977179
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1649977179
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1649977179
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1649977179
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1649977179
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1649977179
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1649977179
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1649977179
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1649977179
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_613
timestamp 1649977179
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_3
timestamp 1649977179
transform 1 0 1380 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_11
timestamp 1649977179
transform 1 0 2116 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_30
timestamp 1649977179
transform 1 0 3864 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_42
timestamp 1649977179
transform 1 0 4968 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_48
timestamp 1649977179
transform 1 0 5520 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_62
timestamp 1649977179
transform 1 0 6808 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_66
timestamp 1649977179
transform 1 0 7176 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_77
timestamp 1649977179
transform 1 0 8188 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_83
timestamp 1649977179
transform 1 0 8740 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_95
timestamp 1649977179
transform 1 0 9844 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_104
timestamp 1649977179
transform 1 0 10672 0 -1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_67_115
timestamp 1649977179
transform 1 0 11684 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_127
timestamp 1649977179
transform 1 0 12788 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_131
timestamp 1649977179
transform 1 0 13156 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_143
timestamp 1649977179
transform 1 0 14260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_155
timestamp 1649977179
transform 1 0 15364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1649977179
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_169
timestamp 1649977179
transform 1 0 16652 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1649977179
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1649977179
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1649977179
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1649977179
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_225
timestamp 1649977179
transform 1 0 21804 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_233
timestamp 1649977179
transform 1 0 22540 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_241
timestamp 1649977179
transform 1 0 23276 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_245
timestamp 1649977179
transform 1 0 23644 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_248
timestamp 1649977179
transform 1 0 23920 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_260
timestamp 1649977179
transform 1 0 25024 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_272
timestamp 1649977179
transform 1 0 26128 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_283
timestamp 1649977179
transform 1 0 27140 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_295
timestamp 1649977179
transform 1 0 28244 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_307
timestamp 1649977179
transform 1 0 29348 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_312
timestamp 1649977179
transform 1 0 29808 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_324
timestamp 1649977179
transform 1 0 30912 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1649977179
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1649977179
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1649977179
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1649977179
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1649977179
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1649977179
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1649977179
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1649977179
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1649977179
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1649977179
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1649977179
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1649977179
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1649977179
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1649977179
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1649977179
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1649977179
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1649977179
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1649977179
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1649977179
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1649977179
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1649977179
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1649977179
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1649977179
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1649977179
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1649977179
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1649977179
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1649977179
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1649977179
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1649977179
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1649977179
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_617
timestamp 1649977179
transform 1 0 57868 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_621
timestamp 1649977179
transform 1 0 58236 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1649977179
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1649977179
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1649977179
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_37
timestamp 1649977179
transform 1 0 4508 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_43
timestamp 1649977179
transform 1 0 5060 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_47
timestamp 1649977179
transform 1 0 5428 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_64
timestamp 1649977179
transform 1 0 6992 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_78
timestamp 1649977179
transform 1 0 8280 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_68_85
timestamp 1649977179
transform 1 0 8924 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_104
timestamp 1649977179
transform 1 0 10672 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_113
timestamp 1649977179
transform 1 0 11500 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_119
timestamp 1649977179
transform 1 0 12052 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_136
timestamp 1649977179
transform 1 0 13616 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_151
timestamp 1649977179
transform 1 0 14996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_163
timestamp 1649977179
transform 1 0 16100 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_68_173
timestamp 1649977179
transform 1 0 17020 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_185
timestamp 1649977179
transform 1 0 18124 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_193
timestamp 1649977179
transform 1 0 18860 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1649977179
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_209
timestamp 1649977179
transform 1 0 20332 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_215
timestamp 1649977179
transform 1 0 20884 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_232
timestamp 1649977179
transform 1 0 22448 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_68_246
timestamp 1649977179
transform 1 0 23736 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_269
timestamp 1649977179
transform 1 0 25852 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_281
timestamp 1649977179
transform 1 0 26956 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_300
timestamp 1649977179
transform 1 0 28704 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_68_309
timestamp 1649977179
transform 1 0 29532 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_319
timestamp 1649977179
transform 1 0 30452 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_331
timestamp 1649977179
transform 1 0 31556 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_340
timestamp 1649977179
transform 1 0 32384 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_352
timestamp 1649977179
transform 1 0 33488 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1649977179
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1649977179
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1649977179
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1649977179
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1649977179
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1649977179
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1649977179
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1649977179
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1649977179
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1649977179
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1649977179
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1649977179
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1649977179
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1649977179
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1649977179
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1649977179
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1649977179
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1649977179
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1649977179
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1649977179
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1649977179
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1649977179
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1649977179
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1649977179
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1649977179
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_601
timestamp 1649977179
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_613
timestamp 1649977179
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1649977179
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_15
timestamp 1649977179
transform 1 0 2484 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_32
timestamp 1649977179
transform 1 0 4048 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_44
timestamp 1649977179
transform 1 0 5152 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_57
timestamp 1649977179
transform 1 0 6348 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_64
timestamp 1649977179
transform 1 0 6992 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_84
timestamp 1649977179
transform 1 0 8832 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_104
timestamp 1649977179
transform 1 0 10672 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_69_121
timestamp 1649977179
transform 1 0 12236 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_143
timestamp 1649977179
transform 1 0 14260 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1649977179
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1649977179
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1649977179
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_185
timestamp 1649977179
transform 1 0 18124 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_205
timestamp 1649977179
transform 1 0 19964 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_213
timestamp 1649977179
transform 1 0 20700 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_220
timestamp 1649977179
transform 1 0 21344 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_225
timestamp 1649977179
transform 1 0 21804 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_231
timestamp 1649977179
transform 1 0 22356 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_240
timestamp 1649977179
transform 1 0 23184 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_260
timestamp 1649977179
transform 1 0 25024 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_272
timestamp 1649977179
transform 1 0 26128 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_281
timestamp 1649977179
transform 1 0 26956 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_284
timestamp 1649977179
transform 1 0 27232 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_296
timestamp 1649977179
transform 1 0 28336 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1649977179
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1649977179
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1649977179
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1649977179
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1649977179
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1649977179
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1649977179
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1649977179
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1649977179
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1649977179
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1649977179
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1649977179
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1649977179
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1649977179
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1649977179
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1649977179
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1649977179
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1649977179
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1649977179
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1649977179
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1649977179
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1649977179
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1649977179
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1649977179
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1649977179
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1649977179
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1649977179
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1649977179
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1649977179
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1649977179
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1649977179
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1649977179
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1649977179
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1649977179
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_617
timestamp 1649977179
transform 1 0 57868 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1649977179
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1649977179
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1649977179
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_34
timestamp 1649977179
transform 1 0 4232 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_46
timestamp 1649977179
transform 1 0 5336 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_70_70
timestamp 1649977179
transform 1 0 7544 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_82
timestamp 1649977179
transform 1 0 8648 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_85
timestamp 1649977179
transform 1 0 8924 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_91
timestamp 1649977179
transform 1 0 9476 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_100
timestamp 1649977179
transform 1 0 10304 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_120
timestamp 1649977179
transform 1 0 12144 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_126
timestamp 1649977179
transform 1 0 12696 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_130
timestamp 1649977179
transform 1 0 13064 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_136
timestamp 1649977179
transform 1 0 13616 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_151
timestamp 1649977179
transform 1 0 14996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_179
timestamp 1649977179
transform 1 0 17572 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_187
timestamp 1649977179
transform 1 0 18308 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_192
timestamp 1649977179
transform 1 0 18768 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_213
timestamp 1649977179
transform 1 0 20700 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_233
timestamp 1649977179
transform 1 0 22540 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_237
timestamp 1649977179
transform 1 0 22908 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_243
timestamp 1649977179
transform 1 0 23460 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1649977179
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1649977179
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1649977179
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_277
timestamp 1649977179
transform 1 0 26588 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1649977179
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1649977179
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1649977179
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_321
timestamp 1649977179
transform 1 0 30636 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_343
timestamp 1649977179
transform 1 0 32660 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_355
timestamp 1649977179
transform 1 0 33764 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1649977179
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1649977179
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1649977179
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1649977179
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1649977179
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1649977179
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1649977179
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1649977179
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1649977179
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1649977179
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1649977179
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1649977179
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1649977179
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1649977179
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1649977179
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1649977179
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1649977179
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1649977179
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1649977179
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1649977179
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1649977179
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1649977179
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1649977179
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1649977179
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1649977179
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1649977179
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1649977179
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_613
timestamp 1649977179
transform 1 0 57500 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_617
timestamp 1649977179
transform 1 0 57868 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_621
timestamp 1649977179
transform 1 0 58236 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1649977179
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1649977179
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1649977179
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1649977179
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1649977179
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1649977179
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_65
timestamp 1649977179
transform 1 0 7084 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_71
timestamp 1649977179
transform 1 0 7636 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_83
timestamp 1649977179
transform 1 0 8740 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_95
timestamp 1649977179
transform 1 0 9844 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_104
timestamp 1649977179
transform 1 0 10672 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1649977179
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_133
timestamp 1649977179
transform 1 0 13340 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_145
timestamp 1649977179
transform 1 0 14444 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_154
timestamp 1649977179
transform 1 0 15272 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_160
timestamp 1649977179
transform 1 0 15824 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_71_174
timestamp 1649977179
transform 1 0 17112 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_180
timestamp 1649977179
transform 1 0 17664 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_189
timestamp 1649977179
transform 1 0 18492 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_201
timestamp 1649977179
transform 1 0 19596 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_210
timestamp 1649977179
transform 1 0 20424 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_216
timestamp 1649977179
transform 1 0 20976 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_71_225
timestamp 1649977179
transform 1 0 21804 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_235
timestamp 1649977179
transform 1 0 22724 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_239
timestamp 1649977179
transform 1 0 23092 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_242
timestamp 1649977179
transform 1 0 23368 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_254
timestamp 1649977179
transform 1 0 24472 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_266
timestamp 1649977179
transform 1 0 25576 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_278
timestamp 1649977179
transform 1 0 26680 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1649977179
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1649977179
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1649977179
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1649977179
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1649977179
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1649977179
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1649977179
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1649977179
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1649977179
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1649977179
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1649977179
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1649977179
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1649977179
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1649977179
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1649977179
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1649977179
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1649977179
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1649977179
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1649977179
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1649977179
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1649977179
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1649977179
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1649977179
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1649977179
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1649977179
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1649977179
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1649977179
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1649977179
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1649977179
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1649977179
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1649977179
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1649977179
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1649977179
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1649977179
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1649977179
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1649977179
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_617
timestamp 1649977179
transform 1 0 57868 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1649977179
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1649977179
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1649977179
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1649977179
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1649977179
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1649977179
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1649977179
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1649977179
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1649977179
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1649977179
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_97
timestamp 1649977179
transform 1 0 10028 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_102
timestamp 1649977179
transform 1 0 10488 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_114
timestamp 1649977179
transform 1 0 11592 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_122
timestamp 1649977179
transform 1 0 12328 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_130
timestamp 1649977179
transform 1 0 13064 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_136
timestamp 1649977179
transform 1 0 13616 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_149
timestamp 1649977179
transform 1 0 14812 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_155
timestamp 1649977179
transform 1 0 15364 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_159
timestamp 1649977179
transform 1 0 15732 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_168
timestamp 1649977179
transform 1 0 16560 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_180
timestamp 1649977179
transform 1 0 17664 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_188
timestamp 1649977179
transform 1 0 18400 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_191
timestamp 1649977179
transform 1 0 18676 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1649977179
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_202
timestamp 1649977179
transform 1 0 19688 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_208
timestamp 1649977179
transform 1 0 20240 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_220
timestamp 1649977179
transform 1 0 21344 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_232
timestamp 1649977179
transform 1 0 22448 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_244
timestamp 1649977179
transform 1 0 23552 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1649977179
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1649977179
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1649977179
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1649977179
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1649977179
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1649977179
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1649977179
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1649977179
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1649977179
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1649977179
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1649977179
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1649977179
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1649977179
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1649977179
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1649977179
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1649977179
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1649977179
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1649977179
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1649977179
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1649977179
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1649977179
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1649977179
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1649977179
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1649977179
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1649977179
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1649977179
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1649977179
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1649977179
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1649977179
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1649977179
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1649977179
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1649977179
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1649977179
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1649977179
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1649977179
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1649977179
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1649977179
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1649977179
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_613
timestamp 1649977179
transform 1 0 57500 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_617
timestamp 1649977179
transform 1 0 57868 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_621
timestamp 1649977179
transform 1 0 58236 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1649977179
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1649977179
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1649977179
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1649977179
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1649977179
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1649977179
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1649977179
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1649977179
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1649977179
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1649977179
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1649977179
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1649977179
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1649977179
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1649977179
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1649977179
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1649977179
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1649977179
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1649977179
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_174
timestamp 1649977179
transform 1 0 17112 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_182
timestamp 1649977179
transform 1 0 17848 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_194
timestamp 1649977179
transform 1 0 18952 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_206
timestamp 1649977179
transform 1 0 20056 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_218
timestamp 1649977179
transform 1 0 21160 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1649977179
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1649977179
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1649977179
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1649977179
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1649977179
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1649977179
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1649977179
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1649977179
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1649977179
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1649977179
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1649977179
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1649977179
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1649977179
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1649977179
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1649977179
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1649977179
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1649977179
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1649977179
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1649977179
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1649977179
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1649977179
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1649977179
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1649977179
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1649977179
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1649977179
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1649977179
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1649977179
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1649977179
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1649977179
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1649977179
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1649977179
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1649977179
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1649977179
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1649977179
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1649977179
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1649977179
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1649977179
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1649977179
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1649977179
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1649977179
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1649977179
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1649977179
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_617
timestamp 1649977179
transform 1 0 57868 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1649977179
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1649977179
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1649977179
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1649977179
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1649977179
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1649977179
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1649977179
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1649977179
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1649977179
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1649977179
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1649977179
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1649977179
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1649977179
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1649977179
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1649977179
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1649977179
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1649977179
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_165
timestamp 1649977179
transform 1 0 16284 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_170
timestamp 1649977179
transform 1 0 16744 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_182
timestamp 1649977179
transform 1 0 17848 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_194
timestamp 1649977179
transform 1 0 18952 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1649977179
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1649977179
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1649977179
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1649977179
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1649977179
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1649977179
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1649977179
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1649977179
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1649977179
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1649977179
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1649977179
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1649977179
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1649977179
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1649977179
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1649977179
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1649977179
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1649977179
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1649977179
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1649977179
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1649977179
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1649977179
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1649977179
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1649977179
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1649977179
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1649977179
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1649977179
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1649977179
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1649977179
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1649977179
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1649977179
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1649977179
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1649977179
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1649977179
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1649977179
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1649977179
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1649977179
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1649977179
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1649977179
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1649977179
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1649977179
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1649977179
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1649977179
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1649977179
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1649977179
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_613
timestamp 1649977179
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1649977179
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1649977179
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1649977179
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1649977179
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1649977179
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1649977179
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1649977179
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1649977179
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1649977179
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1649977179
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1649977179
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1649977179
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1649977179
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1649977179
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1649977179
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1649977179
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1649977179
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1649977179
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1649977179
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1649977179
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1649977179
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1649977179
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1649977179
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1649977179
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1649977179
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1649977179
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1649977179
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1649977179
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1649977179
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1649977179
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1649977179
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1649977179
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1649977179
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1649977179
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1649977179
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1649977179
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1649977179
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1649977179
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1649977179
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1649977179
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1649977179
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1649977179
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1649977179
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1649977179
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1649977179
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1649977179
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1649977179
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1649977179
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1649977179
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1649977179
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1649977179
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1649977179
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1649977179
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1649977179
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1649977179
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1649977179
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1649977179
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1649977179
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1649977179
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1649977179
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1649977179
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1649977179
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1649977179
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1649977179
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1649977179
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1649977179
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_617
timestamp 1649977179
transform 1 0 57868 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_621
timestamp 1649977179
transform 1 0 58236 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1649977179
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1649977179
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1649977179
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1649977179
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1649977179
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1649977179
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1649977179
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1649977179
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1649977179
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1649977179
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1649977179
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1649977179
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1649977179
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1649977179
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1649977179
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1649977179
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1649977179
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1649977179
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1649977179
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1649977179
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1649977179
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1649977179
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1649977179
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1649977179
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1649977179
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1649977179
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1649977179
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1649977179
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1649977179
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1649977179
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1649977179
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1649977179
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1649977179
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1649977179
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1649977179
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1649977179
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1649977179
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1649977179
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1649977179
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1649977179
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1649977179
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1649977179
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1649977179
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1649977179
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1649977179
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1649977179
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1649977179
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1649977179
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1649977179
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1649977179
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1649977179
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1649977179
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1649977179
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1649977179
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1649977179
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1649977179
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1649977179
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1649977179
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1649977179
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1649977179
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1649977179
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1649977179
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1649977179
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1649977179
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1649977179
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_613
timestamp 1649977179
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1649977179
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1649977179
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1649977179
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1649977179
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1649977179
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1649977179
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1649977179
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1649977179
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1649977179
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1649977179
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1649977179
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1649977179
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1649977179
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1649977179
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1649977179
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1649977179
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1649977179
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1649977179
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1649977179
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1649977179
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1649977179
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1649977179
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1649977179
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1649977179
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1649977179
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1649977179
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1649977179
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1649977179
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1649977179
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1649977179
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1649977179
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1649977179
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1649977179
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1649977179
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1649977179
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1649977179
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1649977179
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1649977179
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1649977179
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1649977179
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1649977179
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1649977179
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1649977179
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1649977179
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1649977179
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1649977179
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1649977179
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1649977179
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1649977179
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1649977179
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1649977179
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1649977179
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1649977179
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1649977179
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1649977179
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1649977179
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1649977179
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1649977179
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1649977179
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1649977179
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1649977179
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1649977179
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1649977179
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1649977179
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1649977179
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1649977179
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_617
timestamp 1649977179
transform 1 0 57868 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_621
timestamp 1649977179
transform 1 0 58236 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1649977179
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1649977179
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1649977179
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1649977179
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1649977179
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1649977179
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1649977179
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1649977179
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1649977179
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1649977179
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1649977179
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1649977179
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1649977179
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1649977179
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1649977179
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1649977179
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1649977179
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1649977179
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1649977179
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1649977179
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1649977179
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1649977179
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1649977179
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1649977179
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1649977179
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1649977179
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1649977179
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1649977179
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1649977179
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1649977179
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1649977179
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1649977179
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1649977179
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1649977179
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1649977179
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1649977179
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1649977179
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1649977179
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1649977179
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1649977179
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1649977179
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1649977179
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1649977179
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1649977179
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1649977179
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1649977179
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1649977179
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1649977179
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1649977179
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1649977179
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1649977179
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1649977179
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1649977179
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1649977179
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1649977179
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1649977179
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1649977179
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1649977179
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1649977179
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1649977179
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1649977179
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1649977179
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1649977179
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1649977179
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1649977179
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_613
timestamp 1649977179
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1649977179
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1649977179
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1649977179
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1649977179
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1649977179
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1649977179
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1649977179
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1649977179
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1649977179
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1649977179
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1649977179
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1649977179
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1649977179
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1649977179
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1649977179
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1649977179
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1649977179
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1649977179
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1649977179
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1649977179
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1649977179
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1649977179
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1649977179
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1649977179
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1649977179
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1649977179
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1649977179
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1649977179
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1649977179
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1649977179
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1649977179
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1649977179
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1649977179
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1649977179
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1649977179
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1649977179
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1649977179
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1649977179
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1649977179
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1649977179
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1649977179
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1649977179
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1649977179
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1649977179
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1649977179
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1649977179
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1649977179
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1649977179
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1649977179
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1649977179
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1649977179
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1649977179
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1649977179
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1649977179
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1649977179
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1649977179
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1649977179
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1649977179
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1649977179
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1649977179
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1649977179
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1649977179
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1649977179
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1649977179
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1649977179
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1649977179
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_617
timestamp 1649977179
transform 1 0 57868 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1649977179
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1649977179
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1649977179
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1649977179
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1649977179
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1649977179
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1649977179
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1649977179
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1649977179
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1649977179
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1649977179
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1649977179
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1649977179
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1649977179
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1649977179
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1649977179
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1649977179
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1649977179
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1649977179
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1649977179
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1649977179
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1649977179
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1649977179
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1649977179
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1649977179
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1649977179
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1649977179
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1649977179
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1649977179
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1649977179
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1649977179
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1649977179
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1649977179
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1649977179
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1649977179
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1649977179
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1649977179
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1649977179
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1649977179
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1649977179
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1649977179
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1649977179
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1649977179
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1649977179
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1649977179
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1649977179
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1649977179
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1649977179
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1649977179
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1649977179
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1649977179
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1649977179
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1649977179
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1649977179
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1649977179
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1649977179
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1649977179
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1649977179
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1649977179
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1649977179
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1649977179
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1649977179
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1649977179
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1649977179
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1649977179
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_613
timestamp 1649977179
transform 1 0 57500 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_617
timestamp 1649977179
transform 1 0 57868 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_621
timestamp 1649977179
transform 1 0 58236 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1649977179
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1649977179
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1649977179
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1649977179
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1649977179
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1649977179
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1649977179
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1649977179
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1649977179
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1649977179
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1649977179
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1649977179
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1649977179
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1649977179
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1649977179
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1649977179
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1649977179
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1649977179
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1649977179
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1649977179
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1649977179
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1649977179
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1649977179
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1649977179
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1649977179
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1649977179
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1649977179
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1649977179
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1649977179
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1649977179
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1649977179
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1649977179
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1649977179
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1649977179
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1649977179
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1649977179
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1649977179
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1649977179
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1649977179
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1649977179
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1649977179
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1649977179
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1649977179
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1649977179
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1649977179
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1649977179
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1649977179
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1649977179
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1649977179
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1649977179
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1649977179
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1649977179
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1649977179
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1649977179
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1649977179
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1649977179
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1649977179
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1649977179
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1649977179
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1649977179
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1649977179
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1649977179
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1649977179
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1649977179
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1649977179
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1649977179
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_617
timestamp 1649977179
transform 1 0 57868 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1649977179
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1649977179
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1649977179
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1649977179
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1649977179
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1649977179
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1649977179
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1649977179
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1649977179
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1649977179
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1649977179
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1649977179
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1649977179
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1649977179
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1649977179
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1649977179
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1649977179
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1649977179
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1649977179
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1649977179
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1649977179
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1649977179
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1649977179
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1649977179
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1649977179
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1649977179
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1649977179
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1649977179
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1649977179
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1649977179
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1649977179
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1649977179
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1649977179
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1649977179
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1649977179
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1649977179
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1649977179
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1649977179
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1649977179
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1649977179
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1649977179
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1649977179
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1649977179
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1649977179
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1649977179
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1649977179
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1649977179
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1649977179
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1649977179
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1649977179
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1649977179
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1649977179
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1649977179
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1649977179
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1649977179
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1649977179
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1649977179
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1649977179
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1649977179
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1649977179
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1649977179
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1649977179
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1649977179
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1649977179
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1649977179
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_613
timestamp 1649977179
transform 1 0 57500 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_617
timestamp 1649977179
transform 1 0 57868 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_621
timestamp 1649977179
transform 1 0 58236 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1649977179
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1649977179
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1649977179
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1649977179
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1649977179
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1649977179
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1649977179
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1649977179
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1649977179
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1649977179
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1649977179
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1649977179
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1649977179
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1649977179
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1649977179
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1649977179
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1649977179
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1649977179
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1649977179
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1649977179
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1649977179
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1649977179
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1649977179
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1649977179
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1649977179
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1649977179
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1649977179
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1649977179
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1649977179
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1649977179
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1649977179
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1649977179
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1649977179
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1649977179
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1649977179
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1649977179
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1649977179
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1649977179
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1649977179
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1649977179
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1649977179
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1649977179
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1649977179
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1649977179
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1649977179
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1649977179
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1649977179
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1649977179
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1649977179
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1649977179
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1649977179
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1649977179
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1649977179
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1649977179
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1649977179
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1649977179
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1649977179
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1649977179
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1649977179
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1649977179
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1649977179
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1649977179
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1649977179
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1649977179
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1649977179
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1649977179
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_617
timestamp 1649977179
transform 1 0 57868 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_84_6
timestamp 1649977179
transform 1 0 1656 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_18
timestamp 1649977179
transform 1 0 2760 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_26
timestamp 1649977179
transform 1 0 3496 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1649977179
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1649977179
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1649977179
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1649977179
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1649977179
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1649977179
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1649977179
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1649977179
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1649977179
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1649977179
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1649977179
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1649977179
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1649977179
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1649977179
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1649977179
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1649977179
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1649977179
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1649977179
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1649977179
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1649977179
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1649977179
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1649977179
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1649977179
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1649977179
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1649977179
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1649977179
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1649977179
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1649977179
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1649977179
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1649977179
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1649977179
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1649977179
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1649977179
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1649977179
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1649977179
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1649977179
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1649977179
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1649977179
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1649977179
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1649977179
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1649977179
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1649977179
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1649977179
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1649977179
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1649977179
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1649977179
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1649977179
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1649977179
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1649977179
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1649977179
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1649977179
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1649977179
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1649977179
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1649977179
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1649977179
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1649977179
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1649977179
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1649977179
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1649977179
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1649977179
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1649977179
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1649977179
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_613
timestamp 1649977179
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1649977179
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1649977179
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1649977179
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1649977179
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1649977179
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1649977179
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1649977179
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1649977179
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1649977179
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1649977179
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1649977179
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1649977179
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1649977179
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1649977179
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1649977179
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1649977179
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1649977179
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1649977179
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1649977179
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1649977179
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1649977179
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1649977179
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1649977179
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1649977179
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1649977179
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1649977179
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1649977179
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1649977179
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1649977179
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1649977179
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1649977179
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1649977179
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1649977179
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1649977179
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1649977179
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1649977179
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1649977179
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1649977179
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1649977179
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1649977179
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1649977179
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1649977179
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1649977179
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1649977179
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1649977179
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1649977179
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1649977179
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1649977179
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1649977179
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1649977179
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1649977179
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1649977179
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1649977179
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1649977179
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1649977179
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1649977179
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1649977179
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1649977179
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1649977179
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1649977179
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1649977179
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1649977179
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1649977179
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1649977179
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1649977179
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1649977179
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_617
timestamp 1649977179
transform 1 0 57868 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_621
timestamp 1649977179
transform 1 0 58236 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_6
timestamp 1649977179
transform 1 0 1656 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_18
timestamp 1649977179
transform 1 0 2760 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_26
timestamp 1649977179
transform 1 0 3496 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1649977179
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1649977179
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1649977179
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1649977179
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1649977179
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1649977179
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1649977179
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1649977179
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1649977179
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1649977179
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1649977179
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1649977179
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1649977179
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1649977179
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1649977179
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1649977179
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1649977179
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1649977179
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1649977179
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1649977179
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1649977179
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1649977179
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1649977179
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1649977179
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1649977179
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1649977179
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1649977179
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1649977179
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1649977179
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1649977179
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1649977179
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1649977179
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1649977179
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1649977179
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1649977179
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1649977179
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1649977179
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1649977179
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1649977179
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1649977179
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1649977179
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1649977179
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1649977179
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1649977179
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1649977179
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1649977179
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1649977179
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1649977179
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1649977179
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1649977179
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1649977179
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1649977179
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1649977179
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1649977179
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1649977179
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1649977179
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1649977179
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1649977179
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1649977179
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1649977179
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1649977179
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1649977179
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_613
timestamp 1649977179
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1649977179
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1649977179
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1649977179
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1649977179
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1649977179
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1649977179
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1649977179
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1649977179
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1649977179
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1649977179
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1649977179
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1649977179
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1649977179
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1649977179
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1649977179
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1649977179
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1649977179
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1649977179
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1649977179
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1649977179
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1649977179
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1649977179
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1649977179
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1649977179
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1649977179
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1649977179
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1649977179
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1649977179
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1649977179
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1649977179
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1649977179
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1649977179
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1649977179
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1649977179
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1649977179
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1649977179
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1649977179
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1649977179
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1649977179
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1649977179
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1649977179
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1649977179
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1649977179
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1649977179
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1649977179
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1649977179
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1649977179
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1649977179
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1649977179
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1649977179
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1649977179
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1649977179
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1649977179
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1649977179
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1649977179
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1649977179
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1649977179
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1649977179
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1649977179
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1649977179
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1649977179
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1649977179
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1649977179
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1649977179
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1649977179
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1649977179
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_87_617
timestamp 1649977179
transform 1 0 57868 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_621
timestamp 1649977179
transform 1 0 58236 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_6
timestamp 1649977179
transform 1 0 1656 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_18
timestamp 1649977179
transform 1 0 2760 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_26
timestamp 1649977179
transform 1 0 3496 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1649977179
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1649977179
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1649977179
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1649977179
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1649977179
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1649977179
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1649977179
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1649977179
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1649977179
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1649977179
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1649977179
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1649977179
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1649977179
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1649977179
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1649977179
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1649977179
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1649977179
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1649977179
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1649977179
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1649977179
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1649977179
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1649977179
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1649977179
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1649977179
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1649977179
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1649977179
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1649977179
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1649977179
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1649977179
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1649977179
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1649977179
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1649977179
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1649977179
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1649977179
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1649977179
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1649977179
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1649977179
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1649977179
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1649977179
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1649977179
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1649977179
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1649977179
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1649977179
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1649977179
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1649977179
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1649977179
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1649977179
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1649977179
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1649977179
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1649977179
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1649977179
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1649977179
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1649977179
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1649977179
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1649977179
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1649977179
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1649977179
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1649977179
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1649977179
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1649977179
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1649977179
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1649977179
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_613
timestamp 1649977179
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1649977179
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1649977179
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1649977179
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1649977179
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1649977179
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1649977179
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1649977179
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1649977179
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1649977179
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1649977179
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1649977179
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1649977179
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1649977179
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1649977179
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1649977179
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1649977179
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1649977179
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1649977179
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1649977179
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1649977179
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1649977179
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1649977179
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1649977179
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1649977179
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1649977179
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1649977179
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1649977179
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1649977179
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1649977179
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1649977179
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1649977179
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1649977179
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1649977179
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1649977179
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1649977179
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1649977179
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1649977179
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1649977179
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1649977179
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1649977179
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1649977179
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1649977179
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1649977179
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1649977179
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1649977179
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1649977179
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1649977179
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1649977179
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1649977179
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1649977179
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1649977179
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1649977179
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1649977179
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1649977179
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1649977179
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1649977179
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1649977179
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1649977179
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1649977179
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1649977179
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1649977179
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1649977179
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1649977179
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1649977179
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1649977179
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1649977179
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_617
timestamp 1649977179
transform 1 0 57868 0 -1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_90_6
timestamp 1649977179
transform 1 0 1656 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_18
timestamp 1649977179
transform 1 0 2760 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_26
timestamp 1649977179
transform 1 0 3496 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1649977179
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1649977179
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1649977179
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1649977179
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1649977179
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1649977179
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1649977179
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1649977179
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1649977179
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1649977179
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1649977179
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1649977179
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1649977179
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1649977179
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1649977179
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1649977179
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1649977179
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1649977179
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1649977179
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1649977179
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1649977179
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1649977179
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1649977179
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1649977179
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1649977179
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1649977179
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1649977179
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1649977179
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1649977179
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1649977179
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1649977179
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1649977179
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1649977179
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1649977179
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1649977179
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1649977179
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1649977179
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1649977179
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1649977179
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1649977179
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1649977179
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1649977179
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1649977179
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1649977179
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1649977179
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1649977179
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1649977179
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1649977179
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1649977179
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1649977179
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1649977179
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1649977179
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1649977179
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1649977179
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1649977179
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1649977179
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1649977179
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1649977179
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1649977179
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1649977179
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1649977179
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1649977179
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_613
timestamp 1649977179
transform 1 0 57500 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_617
timestamp 1649977179
transform 1 0 57868 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_621
timestamp 1649977179
transform 1 0 58236 0 1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1649977179
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1649977179
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1649977179
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1649977179
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1649977179
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1649977179
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1649977179
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1649977179
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1649977179
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1649977179
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1649977179
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1649977179
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1649977179
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1649977179
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1649977179
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1649977179
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1649977179
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1649977179
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1649977179
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1649977179
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1649977179
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1649977179
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1649977179
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1649977179
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1649977179
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1649977179
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1649977179
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1649977179
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1649977179
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1649977179
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1649977179
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1649977179
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1649977179
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1649977179
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1649977179
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1649977179
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1649977179
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1649977179
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1649977179
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1649977179
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1649977179
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1649977179
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1649977179
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1649977179
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1649977179
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1649977179
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1649977179
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1649977179
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1649977179
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1649977179
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1649977179
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1649977179
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1649977179
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1649977179
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1649977179
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1649977179
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1649977179
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1649977179
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1649977179
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1649977179
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1649977179
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1649977179
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1649977179
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1649977179
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1649977179
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1649977179
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_617
timestamp 1649977179
transform 1 0 57868 0 -1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_92_6
timestamp 1649977179
transform 1 0 1656 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_18
timestamp 1649977179
transform 1 0 2760 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_26
timestamp 1649977179
transform 1 0 3496 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1649977179
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1649977179
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1649977179
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1649977179
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1649977179
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1649977179
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1649977179
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1649977179
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1649977179
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1649977179
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1649977179
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1649977179
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1649977179
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1649977179
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1649977179
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1649977179
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1649977179
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1649977179
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1649977179
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1649977179
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1649977179
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1649977179
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1649977179
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1649977179
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1649977179
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1649977179
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1649977179
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1649977179
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1649977179
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1649977179
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1649977179
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1649977179
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1649977179
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1649977179
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1649977179
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1649977179
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1649977179
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1649977179
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1649977179
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1649977179
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1649977179
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1649977179
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1649977179
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1649977179
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1649977179
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1649977179
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1649977179
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1649977179
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1649977179
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1649977179
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1649977179
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1649977179
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1649977179
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1649977179
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1649977179
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1649977179
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1649977179
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1649977179
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1649977179
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1649977179
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1649977179
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1649977179
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_613
timestamp 1649977179
transform 1 0 57500 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_617
timestamp 1649977179
transform 1 0 57868 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_621
timestamp 1649977179
transform 1 0 58236 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1649977179
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1649977179
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1649977179
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1649977179
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1649977179
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1649977179
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1649977179
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1649977179
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1649977179
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1649977179
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1649977179
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1649977179
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1649977179
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1649977179
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1649977179
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1649977179
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1649977179
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1649977179
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1649977179
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1649977179
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1649977179
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1649977179
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1649977179
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1649977179
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1649977179
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1649977179
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1649977179
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1649977179
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1649977179
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1649977179
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1649977179
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1649977179
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1649977179
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1649977179
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1649977179
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1649977179
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1649977179
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1649977179
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1649977179
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1649977179
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1649977179
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1649977179
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1649977179
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1649977179
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1649977179
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1649977179
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1649977179
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1649977179
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1649977179
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1649977179
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1649977179
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1649977179
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1649977179
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1649977179
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1649977179
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1649977179
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1649977179
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1649977179
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1649977179
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1649977179
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1649977179
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1649977179
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1649977179
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1649977179
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1649977179
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1649977179
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_617
timestamp 1649977179
transform 1 0 57868 0 -1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_6
timestamp 1649977179
transform 1 0 1656 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_18
timestamp 1649977179
transform 1 0 2760 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_26
timestamp 1649977179
transform 1 0 3496 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1649977179
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1649977179
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1649977179
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1649977179
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1649977179
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1649977179
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1649977179
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1649977179
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1649977179
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1649977179
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1649977179
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1649977179
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1649977179
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1649977179
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1649977179
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1649977179
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1649977179
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1649977179
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1649977179
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1649977179
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1649977179
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1649977179
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1649977179
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1649977179
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1649977179
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1649977179
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1649977179
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1649977179
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1649977179
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1649977179
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1649977179
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1649977179
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1649977179
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1649977179
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1649977179
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1649977179
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1649977179
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1649977179
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1649977179
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1649977179
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1649977179
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1649977179
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1649977179
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1649977179
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1649977179
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1649977179
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1649977179
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1649977179
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1649977179
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1649977179
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1649977179
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1649977179
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1649977179
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1649977179
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1649977179
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1649977179
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1649977179
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1649977179
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1649977179
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1649977179
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1649977179
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1649977179
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1649977179
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1649977179
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1649977179
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1649977179
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1649977179
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1649977179
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1649977179
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1649977179
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1649977179
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1649977179
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1649977179
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1649977179
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1649977179
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1649977179
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1649977179
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1649977179
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1649977179
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1649977179
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1649977179
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1649977179
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1649977179
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1649977179
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1649977179
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1649977179
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1649977179
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1649977179
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1649977179
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1649977179
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1649977179
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1649977179
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1649977179
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1649977179
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1649977179
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1649977179
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1649977179
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1649977179
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1649977179
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1649977179
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1649977179
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1649977179
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1649977179
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1649977179
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1649977179
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1649977179
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1649977179
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1649977179
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1649977179
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1649977179
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1649977179
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1649977179
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1649977179
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1649977179
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1649977179
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1649977179
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1649977179
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1649977179
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1649977179
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1649977179
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1649977179
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1649977179
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1649977179
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1649977179
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1649977179
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1649977179
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1649977179
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1649977179
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1649977179
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_95_617
timestamp 1649977179
transform 1 0 57868 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_621
timestamp 1649977179
transform 1 0 58236 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_6
timestamp 1649977179
transform 1 0 1656 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_18
timestamp 1649977179
transform 1 0 2760 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_26
timestamp 1649977179
transform 1 0 3496 0 1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1649977179
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1649977179
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1649977179
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1649977179
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1649977179
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1649977179
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1649977179
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1649977179
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1649977179
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1649977179
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1649977179
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1649977179
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1649977179
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1649977179
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1649977179
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1649977179
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1649977179
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1649977179
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1649977179
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1649977179
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1649977179
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1649977179
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1649977179
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1649977179
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1649977179
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1649977179
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1649977179
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1649977179
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1649977179
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1649977179
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1649977179
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1649977179
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1649977179
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1649977179
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1649977179
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1649977179
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1649977179
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1649977179
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1649977179
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1649977179
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1649977179
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1649977179
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1649977179
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1649977179
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1649977179
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1649977179
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1649977179
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1649977179
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1649977179
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1649977179
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1649977179
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1649977179
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1649977179
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1649977179
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1649977179
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1649977179
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1649977179
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1649977179
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1649977179
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1649977179
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1649977179
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1649977179
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_613
timestamp 1649977179
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1649977179
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1649977179
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1649977179
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1649977179
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1649977179
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1649977179
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1649977179
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1649977179
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1649977179
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1649977179
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1649977179
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1649977179
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1649977179
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1649977179
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1649977179
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1649977179
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1649977179
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1649977179
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1649977179
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_183
timestamp 1649977179
transform 1 0 17940 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_97_191
timestamp 1649977179
transform 1 0 18676 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_194
timestamp 1649977179
transform 1 0 18952 0 -1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_97_204
timestamp 1649977179
transform 1 0 19872 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_216
timestamp 1649977179
transform 1 0 20976 0 -1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1649977179
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1649977179
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1649977179
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1649977179
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1649977179
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1649977179
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1649977179
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1649977179
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1649977179
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1649977179
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1649977179
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1649977179
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1649977179
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1649977179
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1649977179
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1649977179
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1649977179
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1649977179
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1649977179
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1649977179
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1649977179
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_429
timestamp 1649977179
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1649977179
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1649977179
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1649977179
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1649977179
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1649977179
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1649977179
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1649977179
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1649977179
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1649977179
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1649977179
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1649977179
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1649977179
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1649977179
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1649977179
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1649977179
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1649977179
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1649977179
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1649977179
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1649977179
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1649977179
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_97_617
timestamp 1649977179
transform 1 0 57868 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_621
timestamp 1649977179
transform 1 0 58236 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_6
timestamp 1649977179
transform 1 0 1656 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_18
timestamp 1649977179
transform 1 0 2760 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_26
timestamp 1649977179
transform 1 0 3496 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1649977179
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1649977179
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1649977179
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1649977179
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1649977179
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1649977179
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1649977179
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1649977179
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1649977179
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1649977179
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1649977179
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1649977179
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1649977179
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_153
timestamp 1649977179
transform 1 0 15180 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_161
timestamp 1649977179
transform 1 0 15916 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_164
timestamp 1649977179
transform 1 0 16192 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_98_174
timestamp 1649977179
transform 1 0 17112 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_181
timestamp 1649977179
transform 1 0 17756 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_98_192
timestamp 1649977179
transform 1 0 18768 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_197
timestamp 1649977179
transform 1 0 19228 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_204
timestamp 1649977179
transform 1 0 19872 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_210
timestamp 1649977179
transform 1 0 20424 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_214
timestamp 1649977179
transform 1 0 20792 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_217
timestamp 1649977179
transform 1 0 21068 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_223
timestamp 1649977179
transform 1 0 21620 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_226
timestamp 1649977179
transform 1 0 21896 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_230
timestamp 1649977179
transform 1 0 22264 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_233
timestamp 1649977179
transform 1 0 22540 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_237
timestamp 1649977179
transform 1 0 22908 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_240
timestamp 1649977179
transform 1 0 23184 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_244
timestamp 1649977179
transform 1 0 23552 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_247
timestamp 1649977179
transform 1 0 23828 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1649977179
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_255
timestamp 1649977179
transform 1 0 24564 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_261
timestamp 1649977179
transform 1 0 25116 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_269
timestamp 1649977179
transform 1 0 25852 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_98_273
timestamp 1649977179
transform 1 0 26220 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_98_281
timestamp 1649977179
transform 1 0 26956 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_293
timestamp 1649977179
transform 1 0 28060 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_98_305
timestamp 1649977179
transform 1 0 29164 0 1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_98_311
timestamp 1649977179
transform 1 0 29716 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_323
timestamp 1649977179
transform 1 0 30820 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_326
timestamp 1649977179
transform 1 0 31096 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_338
timestamp 1649977179
transform 1 0 32200 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_350
timestamp 1649977179
transform 1 0 33304 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_98_362
timestamp 1649977179
transform 1 0 34408 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1649977179
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1649977179
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1649977179
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1649977179
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1649977179
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1649977179
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1649977179
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1649977179
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1649977179
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1649977179
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1649977179
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1649977179
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1649977179
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1649977179
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1649977179
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1649977179
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1649977179
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1649977179
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1649977179
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1649977179
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1649977179
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1649977179
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1649977179
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1649977179
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1649977179
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1649977179
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_613
timestamp 1649977179
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1649977179
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1649977179
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1649977179
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1649977179
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1649977179
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1649977179
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1649977179
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1649977179
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1649977179
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1649977179
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1649977179
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1649977179
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1649977179
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_125
timestamp 1649977179
transform 1 0 12604 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_133
timestamp 1649977179
transform 1 0 13340 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_138
timestamp 1649977179
transform 1 0 13800 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_99_144
timestamp 1649977179
transform 1 0 14352 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_156
timestamp 1649977179
transform 1 0 15456 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_99_162
timestamp 1649977179
transform 1 0 16008 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_99_169
timestamp 1649977179
transform 1 0 16652 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_174
timestamp 1649977179
transform 1 0 17112 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_181
timestamp 1649977179
transform 1 0 17756 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_188
timestamp 1649977179
transform 1 0 18400 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_195
timestamp 1649977179
transform 1 0 19044 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_202
timestamp 1649977179
transform 1 0 19688 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_209
timestamp 1649977179
transform 1 0 20332 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_99_220
timestamp 1649977179
transform 1 0 21344 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_225
timestamp 1649977179
transform 1 0 21804 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_229
timestamp 1649977179
transform 1 0 22172 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_236
timestamp 1649977179
transform 1 0 22816 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_243
timestamp 1649977179
transform 1 0 23460 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_250
timestamp 1649977179
transform 1 0 24104 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_257
timestamp 1649977179
transform 1 0 24748 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_264
timestamp 1649977179
transform 1 0 25392 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_272
timestamp 1649977179
transform 1 0 26128 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_276
timestamp 1649977179
transform 1 0 26496 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_284
timestamp 1649977179
transform 1 0 27232 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_99_294
timestamp 1649977179
transform 1 0 28152 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_301
timestamp 1649977179
transform 1 0 28796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_308
timestamp 1649977179
transform 1 0 29440 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_312
timestamp 1649977179
transform 1 0 29808 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_315
timestamp 1649977179
transform 1 0 30084 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_322
timestamp 1649977179
transform 1 0 30728 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1649977179
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1649977179
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_340
timestamp 1649977179
transform 1 0 32384 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_99_346
timestamp 1649977179
transform 1 0 32936 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_358
timestamp 1649977179
transform 1 0 34040 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_370
timestamp 1649977179
transform 1 0 35144 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_377
timestamp 1649977179
transform 1 0 35788 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_383
timestamp 1649977179
transform 1 0 36340 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1649977179
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1649977179
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1649977179
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1649977179
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1649977179
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1649977179
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1649977179
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1649977179
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_461
timestamp 1649977179
transform 1 0 43516 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_467
timestamp 1649977179
transform 1 0 44068 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1649977179
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_485
timestamp 1649977179
transform 1 0 45724 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_492
timestamp 1649977179
transform 1 0 46368 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_498
timestamp 1649977179
transform 1 0 46920 0 -1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1649977179
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1649977179
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1649977179
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1649977179
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1649977179
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1649977179
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1649977179
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1649977179
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1649977179
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1649977179
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1649977179
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1649977179
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_99_617
timestamp 1649977179
transform 1 0 57868 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_621
timestamp 1649977179
transform 1 0 58236 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_6
timestamp 1649977179
transform 1 0 1656 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_18
timestamp 1649977179
transform 1 0 2760 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_26
timestamp 1649977179
transform 1 0 3496 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1649977179
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1649977179
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1649977179
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1649977179
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1649977179
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1649977179
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1649977179
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1649977179
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1649977179
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1649977179
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1649977179
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1649977179
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1649977179
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1649977179
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1649977179
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_179
timestamp 1649977179
transform 1 0 17572 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_185
timestamp 1649977179
transform 1 0 18124 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_192
timestamp 1649977179
transform 1 0 18768 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_197
timestamp 1649977179
transform 1 0 19228 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_201
timestamp 1649977179
transform 1 0 19596 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_208
timestamp 1649977179
transform 1 0 20240 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_214
timestamp 1649977179
transform 1 0 20792 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_226
timestamp 1649977179
transform 1 0 21896 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_238
timestamp 1649977179
transform 1 0 23000 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_250
timestamp 1649977179
transform 1 0 24104 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1649977179
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1649977179
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1649977179
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_289
timestamp 1649977179
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1649977179
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1649977179
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1649977179
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1649977179
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1649977179
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_345
timestamp 1649977179
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1649977179
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1649977179
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1649977179
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1649977179
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1649977179
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1649977179
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1649977179
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1649977179
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_421
timestamp 1649977179
transform 1 0 39836 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_429
timestamp 1649977179
transform 1 0 40572 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1649977179
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_445
timestamp 1649977179
transform 1 0 42044 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_100_450
timestamp 1649977179
transform 1 0 42504 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_462
timestamp 1649977179
transform 1 0 43608 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_474
timestamp 1649977179
transform 1 0 44712 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1649977179
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1649977179
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1649977179
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1649977179
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1649977179
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1649977179
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1649977179
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1649977179
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1649977179
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1649977179
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1649977179
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1649977179
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1649977179
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_601
timestamp 1649977179
transform 1 0 56396 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_609
timestamp 1649977179
transform 1 0 57132 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_614
timestamp 1649977179
transform 1 0 57592 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_621
timestamp 1649977179
transform 1 0 58236 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_3
timestamp 1649977179
transform 1 0 1380 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_7
timestamp 1649977179
transform 1 0 1748 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_12
timestamp 1649977179
transform 1 0 2208 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_18
timestamp 1649977179
transform 1 0 2760 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_26
timestamp 1649977179
transform 1 0 3496 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_33
timestamp 1649977179
transform 1 0 4140 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_41
timestamp 1649977179
transform 1 0 4876 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_46
timestamp 1649977179
transform 1 0 5336 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_54
timestamp 1649977179
transform 1 0 6072 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_57
timestamp 1649977179
transform 1 0 6348 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_63
timestamp 1649977179
transform 1 0 6900 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_75
timestamp 1649977179
transform 1 0 8004 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_80
timestamp 1649977179
transform 1 0 8464 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_85
timestamp 1649977179
transform 1 0 8924 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_97
timestamp 1649977179
transform 1 0 10028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_109
timestamp 1649977179
transform 1 0 11132 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_117
timestamp 1649977179
transform 1 0 11868 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_125
timestamp 1649977179
transform 1 0 12604 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_131
timestamp 1649977179
transform 1 0 13156 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_139
timestamp 1649977179
transform 1 0 13892 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_141
timestamp 1649977179
transform 1 0 14076 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_148
timestamp 1649977179
transform 1 0 14720 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_160
timestamp 1649977179
transform 1 0 15824 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_173
timestamp 1649977179
transform 1 0 17020 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_177
timestamp 1649977179
transform 1 0 17388 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_182
timestamp 1649977179
transform 1 0 17848 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_192
timestamp 1649977179
transform 1 0 18768 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_201
timestamp 1649977179
transform 1 0 19596 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_207
timestamp 1649977179
transform 1 0 20148 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_211
timestamp 1649977179
transform 1 0 20516 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_216
timestamp 1649977179
transform 1 0 20976 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_225
timestamp 1649977179
transform 1 0 21804 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_233
timestamp 1649977179
transform 1 0 22540 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_245
timestamp 1649977179
transform 1 0 23644 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_251
timestamp 1649977179
transform 1 0 24196 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_257
timestamp 1649977179
transform 1 0 24748 0 -1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_101_267
timestamp 1649977179
transform 1 0 25668 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_279
timestamp 1649977179
transform 1 0 26772 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_285
timestamp 1649977179
transform 1 0 27324 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_301
timestamp 1649977179
transform 1 0 28796 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_307
timestamp 1649977179
transform 1 0 29348 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_309
timestamp 1649977179
transform 1 0 29532 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_313
timestamp 1649977179
transform 1 0 29900 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_318
timestamp 1649977179
transform 1 0 30360 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_330
timestamp 1649977179
transform 1 0 31464 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_101_341
timestamp 1649977179
transform 1 0 32476 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_347
timestamp 1649977179
transform 1 0 33028 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_352
timestamp 1649977179
transform 1 0 33488 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_369
timestamp 1649977179
transform 1 0 35052 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_381
timestamp 1649977179
transform 1 0 36156 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_386
timestamp 1649977179
transform 1 0 36616 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_101_393
timestamp 1649977179
transform 1 0 37260 0 -1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_101_403
timestamp 1649977179
transform 1 0 38180 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_415
timestamp 1649977179
transform 1 0 39284 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_419
timestamp 1649977179
transform 1 0 39652 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_425
timestamp 1649977179
transform 1 0 40204 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_101_437
timestamp 1649977179
transform 1 0 41308 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_445
timestamp 1649977179
transform 1 0 42044 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_101_449
timestamp 1649977179
transform 1 0 42412 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_454
timestamp 1649977179
transform 1 0 42872 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_466
timestamp 1649977179
transform 1 0 43976 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_471
timestamp 1649977179
transform 1 0 44436 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_475
timestamp 1649977179
transform 1 0 44804 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_477
timestamp 1649977179
transform 1 0 44988 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_483
timestamp 1649977179
transform 1 0 45540 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_488
timestamp 1649977179
transform 1 0 46000 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_500
timestamp 1649977179
transform 1 0 47104 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_509
timestamp 1649977179
transform 1 0 47932 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_517
timestamp 1649977179
transform 1 0 48668 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_521
timestamp 1649977179
transform 1 0 49036 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_529
timestamp 1649977179
transform 1 0 49772 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_533
timestamp 1649977179
transform 1 0 50140 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_538
timestamp 1649977179
transform 1 0 50600 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_550
timestamp 1649977179
transform 1 0 51704 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_555
timestamp 1649977179
transform 1 0 52164 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_559
timestamp 1649977179
transform 1 0 52532 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_561
timestamp 1649977179
transform 1 0 52716 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_572
timestamp 1649977179
transform 1 0 53728 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_584
timestamp 1649977179
transform 1 0 54832 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_592
timestamp 1649977179
transform 1 0 55568 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_600
timestamp 1649977179
transform 1 0 56304 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_606
timestamp 1649977179
transform 1 0 56856 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_614
timestamp 1649977179
transform 1 0 57592 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_101_617
timestamp 1649977179
transform 1 0 57868 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_621
timestamp 1649977179
transform 1 0 58236 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1649977179
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1649977179
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1649977179
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1649977179
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1649977179
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1649977179
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1649977179
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1649977179
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1649977179
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1649977179
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1649977179
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1649977179
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1649977179
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1649977179
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1649977179
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1649977179
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1649977179
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1649977179
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1649977179
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1649977179
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1649977179
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1649977179
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1649977179
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1649977179
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1649977179
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1649977179
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1649977179
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1649977179
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1649977179
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1649977179
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1649977179
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1649977179
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1649977179
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1649977179
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1649977179
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1649977179
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1649977179
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1649977179
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1649977179
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1649977179
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1649977179
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1649977179
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1649977179
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1649977179
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1649977179
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1649977179
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1649977179
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1649977179
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1649977179
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1649977179
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1649977179
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1649977179
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1649977179
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1649977179
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1649977179
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1649977179
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1649977179
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1649977179
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1649977179
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1649977179
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1649977179
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1649977179
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1649977179
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1649977179
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1649977179
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1649977179
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1649977179
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1649977179
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1649977179
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1649977179
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1649977179
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1649977179
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1649977179
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1649977179
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1649977179
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1649977179
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1649977179
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1649977179
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1649977179
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1649977179
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1649977179
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1649977179
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1649977179
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1649977179
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1649977179
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1649977179
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1649977179
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1649977179
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1649977179
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1649977179
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1649977179
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1649977179
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1649977179
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1649977179
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1649977179
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1649977179
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1649977179
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1649977179
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1649977179
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1649977179
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1649977179
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1649977179
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1649977179
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1649977179
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1649977179
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1649977179
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1649977179
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1649977179
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1649977179
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1649977179
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1649977179
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1649977179
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1649977179
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1649977179
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1649977179
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1649977179
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1649977179
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1649977179
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1649977179
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1649977179
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1649977179
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1649977179
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1649977179
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1649977179
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1649977179
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1649977179
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1649977179
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1649977179
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1649977179
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1649977179
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1649977179
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1649977179
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1649977179
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1649977179
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1649977179
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1649977179
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1649977179
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1649977179
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1649977179
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1649977179
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1649977179
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1649977179
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1649977179
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1649977179
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1649977179
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1649977179
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1649977179
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1649977179
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1649977179
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1649977179
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1649977179
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1649977179
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1649977179
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1649977179
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1649977179
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1649977179
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1649977179
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1649977179
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1649977179
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1649977179
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1649977179
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1649977179
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1649977179
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1649977179
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1649977179
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1649977179
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1649977179
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1649977179
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1649977179
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1649977179
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1649977179
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1649977179
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1649977179
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1649977179
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1649977179
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1649977179
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1649977179
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1649977179
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1649977179
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1649977179
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1649977179
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1649977179
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1649977179
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1649977179
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1649977179
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1649977179
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1649977179
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1649977179
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1649977179
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1649977179
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1649977179
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1649977179
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1649977179
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1649977179
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1649977179
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1649977179
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1649977179
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1649977179
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1649977179
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1649977179
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1649977179
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1649977179
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1649977179
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1649977179
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1649977179
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1649977179
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1649977179
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1649977179
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1649977179
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1649977179
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1649977179
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1649977179
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1649977179
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1649977179
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1649977179
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1649977179
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1649977179
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1649977179
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1649977179
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1649977179
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1649977179
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1649977179
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1649977179
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1649977179
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1649977179
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1649977179
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1649977179
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1649977179
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1649977179
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1649977179
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1649977179
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1649977179
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1649977179
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1649977179
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1649977179
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1649977179
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1649977179
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1649977179
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1649977179
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1649977179
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1649977179
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1649977179
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1649977179
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1649977179
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1649977179
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1649977179
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1649977179
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1649977179
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1649977179
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1649977179
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1649977179
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1649977179
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1649977179
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1649977179
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1649977179
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1649977179
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1649977179
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1649977179
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1649977179
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1649977179
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1649977179
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1649977179
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1649977179
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1649977179
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1649977179
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1649977179
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1649977179
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1649977179
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1649977179
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1649977179
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1649977179
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1649977179
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1649977179
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1649977179
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1649977179
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1649977179
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1649977179
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1649977179
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1649977179
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1649977179
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1649977179
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1649977179
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1649977179
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1649977179
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1649977179
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1649977179
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1649977179
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1649977179
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1649977179
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1649977179
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1649977179
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1649977179
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1649977179
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1649977179
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1649977179
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1649977179
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1649977179
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1649977179
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1649977179
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1649977179
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1649977179
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1649977179
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1649977179
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1649977179
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1649977179
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1649977179
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1649977179
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1649977179
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1649977179
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1649977179
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1649977179
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1649977179
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1649977179
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1649977179
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1649977179
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1649977179
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1649977179
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1649977179
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1649977179
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1649977179
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1649977179
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1649977179
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1649977179
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1649977179
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1649977179
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1649977179
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1649977179
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1649977179
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1649977179
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1649977179
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1649977179
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1649977179
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1649977179
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1649977179
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1649977179
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1649977179
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1649977179
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1649977179
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1649977179
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1649977179
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1649977179
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1649977179
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1649977179
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1649977179
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1649977179
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1649977179
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1649977179
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1649977179
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1649977179
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1649977179
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1649977179
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1649977179
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1649977179
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1649977179
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1649977179
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1649977179
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1649977179
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1649977179
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1649977179
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1649977179
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1649977179
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1649977179
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1649977179
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1649977179
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1649977179
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1649977179
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1649977179
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1649977179
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1649977179
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1649977179
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1649977179
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1649977179
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1649977179
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1649977179
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1649977179
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1649977179
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1649977179
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1649977179
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1649977179
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1649977179
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1649977179
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1649977179
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1649977179
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1649977179
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1649977179
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1649977179
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1649977179
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1649977179
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1649977179
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1649977179
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1649977179
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1649977179
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1649977179
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1649977179
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1649977179
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1649977179
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1649977179
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1649977179
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1649977179
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1649977179
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1649977179
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1649977179
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1649977179
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1649977179
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1649977179
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1649977179
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1649977179
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1649977179
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1649977179
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1649977179
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1649977179
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1649977179
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1649977179
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1649977179
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1649977179
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1649977179
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1649977179
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1649977179
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1649977179
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1649977179
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1649977179
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1649977179
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1649977179
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1649977179
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1649977179
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1649977179
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1649977179
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1649977179
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1649977179
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1649977179
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1649977179
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1649977179
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1649977179
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1649977179
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1649977179
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1649977179
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1649977179
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1649977179
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1649977179
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1649977179
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1649977179
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1649977179
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1649977179
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1649977179
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1649977179
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1649977179
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1649977179
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1649977179
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1649977179
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1649977179
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1649977179
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1649977179
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1649977179
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1649977179
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1649977179
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1649977179
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1649977179
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1649977179
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1649977179
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1649977179
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1649977179
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1649977179
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1649977179
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1649977179
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1649977179
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1649977179
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1649977179
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1649977179
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1649977179
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1649977179
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1649977179
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1649977179
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1649977179
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1649977179
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1649977179
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1649977179
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1649977179
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1649977179
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1649977179
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1649977179
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1649977179
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1649977179
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1649977179
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1649977179
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1649977179
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1649977179
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1649977179
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1649977179
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1649977179
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1649977179
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1649977179
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1649977179
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1649977179
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1649977179
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1649977179
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1649977179
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1649977179
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1649977179
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1649977179
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1649977179
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1649977179
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1649977179
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1649977179
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1649977179
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0855_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0856_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6808 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0857_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9660 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0858_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6900 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0859_
timestamp 1649977179
transform -1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0860_
timestamp 1649977179
transform -1 0 5888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0861_
timestamp 1649977179
transform -1 0 7912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0862_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8740 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0863_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14996 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0864_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5428 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0865_
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _0866_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0867_
timestamp 1649977179
transform -1 0 4600 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0868_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4784 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0869_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5152 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0870_
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0871_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0872_
timestamp 1649977179
transform 1 0 2300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0873_
timestamp 1649977179
transform 1 0 4600 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0874_
timestamp 1649977179
transform 1 0 1932 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0875_
timestamp 1649977179
transform -1 0 2760 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0876_
timestamp 1649977179
transform 1 0 3220 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0877_
timestamp 1649977179
transform -1 0 2576 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0878_
timestamp 1649977179
transform -1 0 2484 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0879_
timestamp 1649977179
transform 1 0 3312 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0880_
timestamp 1649977179
transform -1 0 2576 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0881_
timestamp 1649977179
transform -1 0 1932 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0882_
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0883_
timestamp 1649977179
transform -1 0 2760 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0884_
timestamp 1649977179
transform 1 0 2208 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0885_
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0886_
timestamp 1649977179
transform 1 0 4600 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0887_
timestamp 1649977179
transform -1 0 4692 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0888_
timestamp 1649977179
transform -1 0 3312 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0889_
timestamp 1649977179
transform -1 0 3312 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0890_
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0891_
timestamp 1649977179
transform 1 0 1656 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0892_
timestamp 1649977179
transform -1 0 2484 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0893_
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0894_
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0895_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0896_
timestamp 1649977179
transform 1 0 3036 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0897_
timestamp 1649977179
transform 1 0 2208 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0898_
timestamp 1649977179
transform 1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0899_
timestamp 1649977179
transform 1 0 12604 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0900_
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0901_
timestamp 1649977179
transform -1 0 13340 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0902_
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0903_
timestamp 1649977179
transform 1 0 2116 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0904_
timestamp 1649977179
transform -1 0 2484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0905_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0906_
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0907_
timestamp 1649977179
transform -1 0 7084 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0908_
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0909_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7176 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0910_
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0911_
timestamp 1649977179
transform 1 0 17940 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_4  _0912_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0913_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0914_
timestamp 1649977179
transform -1 0 12144 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0915_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7544 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0916_
timestamp 1649977179
transform -1 0 8188 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0917_
timestamp 1649977179
transform -1 0 11960 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0918_
timestamp 1649977179
transform 1 0 8280 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0919_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0920_
timestamp 1649977179
transform 1 0 7360 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0921_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0922_
timestamp 1649977179
transform -1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0923_
timestamp 1649977179
transform 1 0 3772 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0924_
timestamp 1649977179
transform 1 0 4232 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0925_
timestamp 1649977179
transform -1 0 7268 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0926_
timestamp 1649977179
transform -1 0 3496 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0927_
timestamp 1649977179
transform 1 0 2576 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0928_
timestamp 1649977179
transform -1 0 8004 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0929_
timestamp 1649977179
transform 1 0 6348 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0930_
timestamp 1649977179
transform 1 0 6072 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0931_
timestamp 1649977179
transform -1 0 12420 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0932_
timestamp 1649977179
transform 1 0 6532 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0933_
timestamp 1649977179
transform 1 0 6348 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0934_
timestamp 1649977179
transform -1 0 25484 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0935_
timestamp 1649977179
transform 1 0 14076 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0936_
timestamp 1649977179
transform -1 0 13156 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0937_
timestamp 1649977179
transform -1 0 13064 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0938_
timestamp 1649977179
transform 1 0 14076 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0939_
timestamp 1649977179
transform 1 0 12604 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0940_
timestamp 1649977179
transform 1 0 25852 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0941_
timestamp 1649977179
transform 1 0 16652 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0942_
timestamp 1649977179
transform -1 0 17664 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0943_
timestamp 1649977179
transform -1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0944_
timestamp 1649977179
transform 1 0 16652 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0945_
timestamp 1649977179
transform -1 0 16560 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0946_
timestamp 1649977179
transform -1 0 26220 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0947_
timestamp 1649977179
transform -1 0 15272 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0948_
timestamp 1649977179
transform 1 0 13708 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0949_
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0950_
timestamp 1649977179
transform 1 0 13156 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0951_
timestamp 1649977179
transform 1 0 14076 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0952_
timestamp 1649977179
transform -1 0 17020 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0953_
timestamp 1649977179
transform 1 0 12972 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0954_
timestamp 1649977179
transform 1 0 13248 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0955_
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0956_
timestamp 1649977179
transform -1 0 14628 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0957_
timestamp 1649977179
transform 1 0 12052 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0958_
timestamp 1649977179
transform 1 0 12880 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _0959_
timestamp 1649977179
transform -1 0 11868 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0960_
timestamp 1649977179
transform -1 0 20884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0961_
timestamp 1649977179
transform 1 0 30360 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0962_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0963_
timestamp 1649977179
transform 1 0 30084 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0964_
timestamp 1649977179
transform 1 0 16744 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0965_
timestamp 1649977179
transform 1 0 29900 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0966_
timestamp 1649977179
transform -1 0 30636 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0967_
timestamp 1649977179
transform -1 0 29992 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0968_
timestamp 1649977179
transform -1 0 29992 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0969_
timestamp 1649977179
transform -1 0 29072 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0970_
timestamp 1649977179
transform 1 0 27508 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0971_
timestamp 1649977179
transform -1 0 28152 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0972_
timestamp 1649977179
transform 1 0 27232 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0973_
timestamp 1649977179
transform -1 0 30544 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0974_
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0975_
timestamp 1649977179
transform 1 0 29900 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0976_
timestamp 1649977179
transform 1 0 29072 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0977_
timestamp 1649977179
transform 1 0 31188 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0978_
timestamp 1649977179
transform 1 0 30084 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0979_
timestamp 1649977179
transform 1 0 35144 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0980_
timestamp 1649977179
transform -1 0 34776 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0981_
timestamp 1649977179
transform 1 0 35788 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0982_
timestamp 1649977179
transform -1 0 36708 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0983_
timestamp 1649977179
transform 1 0 35144 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0984_
timestamp 1649977179
transform -1 0 36708 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0985_
timestamp 1649977179
transform 1 0 35052 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0986_
timestamp 1649977179
transform -1 0 36616 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0987_
timestamp 1649977179
transform 1 0 35788 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0988_
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0989_
timestamp 1649977179
transform -1 0 36708 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0990_
timestamp 1649977179
transform 1 0 37076 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0991_
timestamp 1649977179
transform -1 0 36800 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0992_
timestamp 1649977179
transform 1 0 34592 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0993_
timestamp 1649977179
transform -1 0 35420 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0994_
timestamp 1649977179
transform 1 0 32936 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0995_
timestamp 1649977179
transform 1 0 33212 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_2  _0996_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0997_
timestamp 1649977179
transform -1 0 20700 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0998_
timestamp 1649977179
transform -1 0 31096 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0999_
timestamp 1649977179
transform 1 0 30360 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1000_
timestamp 1649977179
transform -1 0 31556 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1001_
timestamp 1649977179
transform -1 0 32568 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1002_
timestamp 1649977179
transform -1 0 31832 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1003_
timestamp 1649977179
transform -1 0 29348 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1004_
timestamp 1649977179
transform 1 0 28336 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1005_
timestamp 1649977179
transform -1 0 29164 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1006_
timestamp 1649977179
transform -1 0 31464 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1007_
timestamp 1649977179
transform 1 0 27600 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1008_
timestamp 1649977179
transform -1 0 28520 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1009_
timestamp 1649977179
transform 1 0 27508 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1010_
timestamp 1649977179
transform -1 0 31832 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1011_
timestamp 1649977179
transform -1 0 31004 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1012_
timestamp 1649977179
transform 1 0 31924 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1013_
timestamp 1649977179
transform -1 0 31556 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1014_
timestamp 1649977179
transform 1 0 32292 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1649977179
transform -1 0 32476 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1016_
timestamp 1649977179
transform -1 0 33764 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1017_
timestamp 1649977179
transform 1 0 32568 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1018_
timestamp 1649977179
transform 1 0 32660 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1019_
timestamp 1649977179
transform 1 0 31924 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1020_
timestamp 1649977179
transform -1 0 34224 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1021_
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1022_
timestamp 1649977179
transform -1 0 34500 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1023_
timestamp 1649977179
transform 1 0 34684 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1024_
timestamp 1649977179
transform -1 0 34500 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1025_
timestamp 1649977179
transform 1 0 33764 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1026_
timestamp 1649977179
transform -1 0 35420 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1027_
timestamp 1649977179
transform 1 0 31464 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1028_
timestamp 1649977179
transform -1 0 32936 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1029_
timestamp 1649977179
transform 1 0 32936 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1030_
timestamp 1649977179
transform 1 0 30268 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1031_
timestamp 1649977179
transform -1 0 32752 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _1032_
timestamp 1649977179
transform 1 0 8004 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1033_
timestamp 1649977179
transform -1 0 9660 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1034_
timestamp 1649977179
transform 1 0 9568 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1035_
timestamp 1649977179
transform 1 0 8372 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1036_
timestamp 1649977179
transform -1 0 8648 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1037_
timestamp 1649977179
transform 1 0 12512 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1038_
timestamp 1649977179
transform -1 0 17112 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1649977179
transform 1 0 5612 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1040_
timestamp 1649977179
transform -1 0 5888 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1041_
timestamp 1649977179
transform 1 0 4784 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1042_
timestamp 1649977179
transform -1 0 5336 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1043_
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1044_
timestamp 1649977179
transform -1 0 4876 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1045_
timestamp 1649977179
transform 1 0 4416 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1046_
timestamp 1649977179
transform 1 0 6624 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1047_
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1048_
timestamp 1649977179
transform 1 0 6348 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1049_
timestamp 1649977179
transform 1 0 11500 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1050_
timestamp 1649977179
transform 1 0 24564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1051_
timestamp 1649977179
transform -1 0 19504 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1052_
timestamp 1649977179
transform 1 0 7176 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1053_
timestamp 1649977179
transform 1 0 16008 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1054_
timestamp 1649977179
transform 1 0 17480 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1055_
timestamp 1649977179
transform 1 0 20240 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1056_
timestamp 1649977179
transform -1 0 20516 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1057_
timestamp 1649977179
transform -1 0 19688 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1058_
timestamp 1649977179
transform -1 0 18492 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1059_
timestamp 1649977179
transform -1 0 20424 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1060_
timestamp 1649977179
transform -1 0 19596 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1061_
timestamp 1649977179
transform 1 0 18768 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1062_
timestamp 1649977179
transform -1 0 20332 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1063_
timestamp 1649977179
transform -1 0 18676 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1064_
timestamp 1649977179
transform -1 0 18676 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1065_
timestamp 1649977179
transform -1 0 18308 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1066_
timestamp 1649977179
transform 1 0 14260 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1067_
timestamp 1649977179
transform -1 0 15732 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1068_
timestamp 1649977179
transform 1 0 14628 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1069_
timestamp 1649977179
transform -1 0 15364 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1070_
timestamp 1649977179
transform -1 0 19504 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1071_
timestamp 1649977179
transform -1 0 18492 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1072_
timestamp 1649977179
transform -1 0 16744 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1073_
timestamp 1649977179
transform -1 0 15916 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1074_
timestamp 1649977179
transform 1 0 16744 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1075_
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1076_
timestamp 1649977179
transform 1 0 9844 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1077_
timestamp 1649977179
transform 1 0 10212 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1078_
timestamp 1649977179
transform 1 0 9844 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1079_
timestamp 1649977179
transform 1 0 9752 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1080_
timestamp 1649977179
transform -1 0 12328 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1081_
timestamp 1649977179
transform 1 0 23828 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1082_
timestamp 1649977179
transform 1 0 11040 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1083_
timestamp 1649977179
transform -1 0 13800 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1084_
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1085_
timestamp 1649977179
transform -1 0 15364 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1086_
timestamp 1649977179
transform 1 0 14260 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1087_
timestamp 1649977179
transform 1 0 24748 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1088_
timestamp 1649977179
transform -1 0 24564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1089_
timestamp 1649977179
transform 1 0 23460 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1090_
timestamp 1649977179
transform -1 0 25208 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1091_
timestamp 1649977179
transform 1 0 23460 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1092_
timestamp 1649977179
transform -1 0 25116 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1093_
timestamp 1649977179
transform 1 0 25484 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1094_
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1095_
timestamp 1649977179
transform 1 0 24380 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1096_
timestamp 1649977179
transform 1 0 24840 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1097_
timestamp 1649977179
transform -1 0 25760 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1098_
timestamp 1649977179
transform 1 0 23460 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1099_
timestamp 1649977179
transform 1 0 23920 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1100_
timestamp 1649977179
transform 1 0 24472 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1101_
timestamp 1649977179
transform -1 0 25852 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1102_
timestamp 1649977179
transform 1 0 24288 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1103_
timestamp 1649977179
transform -1 0 25576 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1104_
timestamp 1649977179
transform 1 0 14904 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1105_
timestamp 1649977179
transform 1 0 20884 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1106_
timestamp 1649977179
transform 1 0 21068 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1107_
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1108_
timestamp 1649977179
transform 1 0 23460 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1109_
timestamp 1649977179
transform -1 0 24656 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1110_
timestamp 1649977179
transform 1 0 21804 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1111_
timestamp 1649977179
transform -1 0 24748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1112_
timestamp 1649977179
transform -1 0 23736 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1113_
timestamp 1649977179
transform -1 0 24196 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1114_
timestamp 1649977179
transform 1 0 23368 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1115_
timestamp 1649977179
transform 1 0 14812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1116_
timestamp 1649977179
transform 1 0 24380 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1117_
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1118_
timestamp 1649977179
transform 1 0 13984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1119_
timestamp 1649977179
transform -1 0 25392 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1120_
timestamp 1649977179
transform 1 0 23184 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1121_
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1122_
timestamp 1649977179
transform 1 0 25760 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1123_
timestamp 1649977179
transform -1 0 25392 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1124_
timestamp 1649977179
transform 1 0 18308 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1125_
timestamp 1649977179
transform -1 0 25576 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1126_
timestamp 1649977179
transform -1 0 25484 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1127_
timestamp 1649977179
transform 1 0 29072 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1128_
timestamp 1649977179
transform 1 0 28152 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1129_
timestamp 1649977179
transform -1 0 28336 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1130_
timestamp 1649977179
transform 1 0 30636 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1131_
timestamp 1649977179
transform 1 0 33028 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1132_
timestamp 1649977179
transform -1 0 32384 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1133_
timestamp 1649977179
transform 1 0 30360 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1134_
timestamp 1649977179
transform 1 0 30176 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1135_
timestamp 1649977179
transform 1 0 31924 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1136_
timestamp 1649977179
transform -1 0 33028 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1137_
timestamp 1649977179
transform 1 0 29532 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1138_
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1139_
timestamp 1649977179
transform -1 0 32016 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1140_
timestamp 1649977179
transform 1 0 27416 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1141_
timestamp 1649977179
transform 1 0 30820 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1142_
timestamp 1649977179
transform -1 0 32844 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1143_
timestamp 1649977179
transform 1 0 27232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1144_
timestamp 1649977179
transform -1 0 29992 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1145_
timestamp 1649977179
transform 1 0 28704 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1146_
timestamp 1649977179
transform 1 0 19688 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1147_
timestamp 1649977179
transform 1 0 22356 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1148_
timestamp 1649977179
transform -1 0 27784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1149_
timestamp 1649977179
transform 1 0 22172 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1150_
timestamp 1649977179
transform 1 0 19136 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1151_
timestamp 1649977179
transform 1 0 25760 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1152_
timestamp 1649977179
transform 1 0 25576 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1153_
timestamp 1649977179
transform -1 0 20056 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1154_
timestamp 1649977179
transform 1 0 20424 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1155_
timestamp 1649977179
transform 1 0 21712 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1156_
timestamp 1649977179
transform -1 0 21160 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1157_
timestamp 1649977179
transform -1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1158_
timestamp 1649977179
transform 1 0 20424 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1159_
timestamp 1649977179
transform 1 0 20332 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1160_
timestamp 1649977179
transform 1 0 20148 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1161_
timestamp 1649977179
transform -1 0 13616 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1162_
timestamp 1649977179
transform 1 0 14444 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1163_
timestamp 1649977179
transform 1 0 13616 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1164_
timestamp 1649977179
transform 1 0 14352 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1165_
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1166_
timestamp 1649977179
transform 1 0 14168 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1167_
timestamp 1649977179
transform -1 0 19688 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1168_
timestamp 1649977179
transform -1 0 28520 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1169_
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1170_
timestamp 1649977179
transform 1 0 17664 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1171_
timestamp 1649977179
transform 1 0 18032 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1172_
timestamp 1649977179
transform 1 0 23276 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1173_
timestamp 1649977179
transform 1 0 23000 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1174_
timestamp 1649977179
transform 1 0 28428 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1175_
timestamp 1649977179
transform 1 0 28336 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1176_
timestamp 1649977179
transform 1 0 29624 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1177_
timestamp 1649977179
transform -1 0 30820 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1178_
timestamp 1649977179
transform 1 0 28612 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1179_
timestamp 1649977179
transform 1 0 29440 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1180_
timestamp 1649977179
transform 1 0 28244 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1181_
timestamp 1649977179
transform 1 0 28152 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1182_
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1183_
timestamp 1649977179
transform 1 0 25944 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1184_
timestamp 1649977179
transform 1 0 25760 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1185_
timestamp 1649977179
transform 1 0 20792 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1186_
timestamp 1649977179
transform 1 0 21528 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1187_
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1188_
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _1189_
timestamp 1649977179
transform 1 0 8004 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1190_
timestamp 1649977179
transform -1 0 23920 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1191_
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1192_
timestamp 1649977179
transform 1 0 35052 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1193_
timestamp 1649977179
transform 1 0 38732 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1194_
timestamp 1649977179
transform 1 0 33764 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1195_
timestamp 1649977179
transform -1 0 38272 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1196_
timestamp 1649977179
transform -1 0 36800 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1197_
timestamp 1649977179
transform 1 0 35236 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1198_
timestamp 1649977179
transform 1 0 38548 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1199_
timestamp 1649977179
transform 1 0 36156 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1200_
timestamp 1649977179
transform 1 0 38364 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1201_
timestamp 1649977179
transform -1 0 37720 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1202_
timestamp 1649977179
transform -1 0 37352 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1203_
timestamp 1649977179
transform 1 0 37444 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1204_
timestamp 1649977179
transform -1 0 38640 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1205_
timestamp 1649977179
transform 1 0 37812 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1206_
timestamp 1649977179
transform -1 0 39376 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1207_
timestamp 1649977179
transform -1 0 39376 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1208_
timestamp 1649977179
transform -1 0 39100 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1209_
timestamp 1649977179
transform -1 0 37720 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1210_
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1211_
timestamp 1649977179
transform 1 0 41124 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1212_
timestamp 1649977179
transform 1 0 33212 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1213_
timestamp 1649977179
transform 1 0 40664 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1214_
timestamp 1649977179
transform 1 0 40296 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1215_
timestamp 1649977179
transform 1 0 40296 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1216_
timestamp 1649977179
transform 1 0 40572 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1217_
timestamp 1649977179
transform 1 0 40204 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1218_
timestamp 1649977179
transform 1 0 40480 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1219_
timestamp 1649977179
transform 1 0 39836 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1220_
timestamp 1649977179
transform 1 0 40572 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1221_
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1222_
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1223_
timestamp 1649977179
transform -1 0 36800 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1224_
timestamp 1649977179
transform -1 0 35972 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1225_
timestamp 1649977179
transform 1 0 35604 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1226_
timestamp 1649977179
transform -1 0 22264 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1227_
timestamp 1649977179
transform -1 0 35420 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1228_
timestamp 1649977179
transform 1 0 35972 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1229_
timestamp 1649977179
transform -1 0 39376 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1230_
timestamp 1649977179
transform 1 0 35788 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1231_
timestamp 1649977179
transform -1 0 37628 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1232_
timestamp 1649977179
transform 1 0 35236 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1233_
timestamp 1649977179
transform 1 0 34960 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1234_
timestamp 1649977179
transform -1 0 36432 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1235_
timestamp 1649977179
transform 1 0 35052 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1236_
timestamp 1649977179
transform -1 0 34684 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1237_
timestamp 1649977179
transform 1 0 34868 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1238_
timestamp 1649977179
transform -1 0 37720 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1239_
timestamp 1649977179
transform -1 0 37536 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1240_
timestamp 1649977179
transform 1 0 38180 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1241_
timestamp 1649977179
transform 1 0 40204 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1242_
timestamp 1649977179
transform -1 0 39100 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1243_
timestamp 1649977179
transform -1 0 38272 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1244_
timestamp 1649977179
transform 1 0 37904 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1245_
timestamp 1649977179
transform -1 0 36892 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1246_
timestamp 1649977179
transform 1 0 37260 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1247_
timestamp 1649977179
transform 1 0 40848 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1248_
timestamp 1649977179
transform 1 0 40020 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1249_
timestamp 1649977179
transform 1 0 40020 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1250_
timestamp 1649977179
transform 1 0 40572 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1251_
timestamp 1649977179
transform 1 0 40204 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1252_
timestamp 1649977179
transform 1 0 40388 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1253_
timestamp 1649977179
transform 1 0 40388 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1254_
timestamp 1649977179
transform 1 0 40664 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1255_
timestamp 1649977179
transform 1 0 40756 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1256_
timestamp 1649977179
transform 1 0 37444 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1257_
timestamp 1649977179
transform -1 0 38456 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1258_
timestamp 1649977179
transform -1 0 37720 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1259_
timestamp 1649977179
transform -1 0 36432 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1260_
timestamp 1649977179
transform -1 0 22816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1261_
timestamp 1649977179
transform 1 0 23184 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1262_
timestamp 1649977179
transform -1 0 27600 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1263_
timestamp 1649977179
transform 1 0 29992 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1264_
timestamp 1649977179
transform -1 0 27876 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1265_
timestamp 1649977179
transform -1 0 31556 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1266_
timestamp 1649977179
transform -1 0 28704 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1267_
timestamp 1649977179
transform 1 0 27140 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1268_
timestamp 1649977179
transform -1 0 27416 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1269_
timestamp 1649977179
transform 1 0 26956 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1270_
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1271_
timestamp 1649977179
transform -1 0 33672 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1272_
timestamp 1649977179
transform -1 0 30360 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1273_
timestamp 1649977179
transform -1 0 30268 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1274_
timestamp 1649977179
transform 1 0 28888 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1275_
timestamp 1649977179
transform 1 0 31372 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1276_
timestamp 1649977179
transform 1 0 29624 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1277_
timestamp 1649977179
transform 1 0 31464 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1278_
timestamp 1649977179
transform -1 0 31464 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1279_
timestamp 1649977179
transform 1 0 31924 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1280_
timestamp 1649977179
transform -1 0 33488 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1281_
timestamp 1649977179
transform 1 0 32936 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1282_
timestamp 1649977179
transform -1 0 33212 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1283_
timestamp 1649977179
transform 1 0 32200 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1284_
timestamp 1649977179
transform 1 0 15916 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1285_
timestamp 1649977179
transform 1 0 24748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1286_
timestamp 1649977179
transform -1 0 33396 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1287_
timestamp 1649977179
transform 1 0 32752 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1288_
timestamp 1649977179
transform -1 0 33212 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1289_
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1290_
timestamp 1649977179
transform -1 0 32844 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1291_
timestamp 1649977179
transform -1 0 26496 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1292_
timestamp 1649977179
transform -1 0 26864 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1293_
timestamp 1649977179
transform -1 0 26864 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1294_
timestamp 1649977179
transform 1 0 25668 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1295_
timestamp 1649977179
transform 1 0 5520 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1296_
timestamp 1649977179
transform 1 0 20884 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1297_
timestamp 1649977179
transform -1 0 17388 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1298_
timestamp 1649977179
transform -1 0 17112 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_2  _1299_
timestamp 1649977179
transform -1 0 11500 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1300_
timestamp 1649977179
transform -1 0 7912 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1301_
timestamp 1649977179
transform -1 0 15824 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1302_
timestamp 1649977179
transform 1 0 7176 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1303_
timestamp 1649977179
transform 1 0 3772 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1304_
timestamp 1649977179
transform -1 0 7268 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1305_
timestamp 1649977179
transform 1 0 4232 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1306_
timestamp 1649977179
transform 1 0 4600 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1307_
timestamp 1649977179
transform -1 0 2024 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1308_
timestamp 1649977179
transform 1 0 2300 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1309_
timestamp 1649977179
transform 1 0 4140 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1310_
timestamp 1649977179
transform 1 0 2116 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1311_
timestamp 1649977179
transform 1 0 2208 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1312_
timestamp 1649977179
transform 1 0 6164 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1313_
timestamp 1649977179
transform 1 0 5428 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1314_
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1315_
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1316_
timestamp 1649977179
transform -1 0 6808 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1317_
timestamp 1649977179
transform -1 0 6072 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1318_
timestamp 1649977179
transform 1 0 22172 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1319_
timestamp 1649977179
transform 1 0 20976 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1320_
timestamp 1649977179
transform -1 0 21344 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1321_
timestamp 1649977179
transform 1 0 20884 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1322_
timestamp 1649977179
transform -1 0 22908 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1323_
timestamp 1649977179
transform 1 0 21804 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1324_
timestamp 1649977179
transform -1 0 25484 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1325_
timestamp 1649977179
transform -1 0 23276 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1326_
timestamp 1649977179
transform -1 0 23184 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1327_
timestamp 1649977179
transform 1 0 26680 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1328_
timestamp 1649977179
transform 1 0 23000 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1329_
timestamp 1649977179
transform -1 0 23736 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1330_
timestamp 1649977179
transform 1 0 15732 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1331_
timestamp 1649977179
transform 1 0 22448 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1332_
timestamp 1649977179
transform 1 0 22264 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1333_
timestamp 1649977179
transform 1 0 17020 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1334_
timestamp 1649977179
transform 1 0 21436 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1335_
timestamp 1649977179
transform -1 0 22908 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1336_
timestamp 1649977179
transform 1 0 11408 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1337_
timestamp 1649977179
transform -1 0 19688 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1338_
timestamp 1649977179
transform 1 0 17940 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1339_
timestamp 1649977179
transform 1 0 18032 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1340_
timestamp 1649977179
transform 1 0 9108 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1341_
timestamp 1649977179
transform -1 0 20608 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1342_
timestamp 1649977179
transform -1 0 19872 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_4  _1343_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7360 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1344_
timestamp 1649977179
transform 1 0 22356 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1345_
timestamp 1649977179
transform -1 0 23184 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1346_
timestamp 1649977179
transform -1 0 22172 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1347_
timestamp 1649977179
transform -1 0 21988 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1348_
timestamp 1649977179
transform 1 0 14260 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1349_
timestamp 1649977179
transform -1 0 22264 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1350_
timestamp 1649977179
transform 1 0 20976 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1351_
timestamp 1649977179
transform -1 0 18032 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1352_
timestamp 1649977179
transform -1 0 17204 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1353_
timestamp 1649977179
transform -1 0 19228 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1354_
timestamp 1649977179
transform -1 0 18308 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1355_
timestamp 1649977179
transform -1 0 17204 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1356_
timestamp 1649977179
transform 1 0 15364 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1357_
timestamp 1649977179
transform -1 0 17480 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1358_
timestamp 1649977179
transform 1 0 16836 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1359_
timestamp 1649977179
transform 1 0 16376 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1360_
timestamp 1649977179
transform -1 0 19412 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1361_
timestamp 1649977179
transform -1 0 18768 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1362_
timestamp 1649977179
transform 1 0 23828 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1363_
timestamp 1649977179
transform -1 0 24748 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1364_
timestamp 1649977179
transform -1 0 27416 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1365_
timestamp 1649977179
transform -1 0 25392 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1366_
timestamp 1649977179
transform -1 0 26036 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1367_
timestamp 1649977179
transform -1 0 25208 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1368_
timestamp 1649977179
transform -1 0 26312 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1369_
timestamp 1649977179
transform -1 0 26312 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1370_
timestamp 1649977179
transform 1 0 27416 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1371_
timestamp 1649977179
transform 1 0 11684 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1372_
timestamp 1649977179
transform -1 0 9476 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1373_
timestamp 1649977179
transform -1 0 25484 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1374_
timestamp 1649977179
transform 1 0 25944 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1375_
timestamp 1649977179
transform 1 0 25760 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1376_
timestamp 1649977179
transform -1 0 24196 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1377_
timestamp 1649977179
transform 1 0 22724 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1378_
timestamp 1649977179
transform -1 0 23736 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1379_
timestamp 1649977179
transform -1 0 23368 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1380_
timestamp 1649977179
transform 1 0 9936 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1381_
timestamp 1649977179
transform 1 0 9752 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1382_
timestamp 1649977179
transform 1 0 9200 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1383_
timestamp 1649977179
transform -1 0 8280 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1384_
timestamp 1649977179
transform 1 0 10856 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1385_
timestamp 1649977179
transform -1 0 12052 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1386_
timestamp 1649977179
transform -1 0 9936 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1387_
timestamp 1649977179
transform 1 0 7728 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1388_
timestamp 1649977179
transform 1 0 7728 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1389_
timestamp 1649977179
transform -1 0 3312 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1390_
timestamp 1649977179
transform -1 0 9200 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1391_
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1392_
timestamp 1649977179
transform 1 0 3404 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1393_
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1394_
timestamp 1649977179
transform 1 0 5428 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1395_
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1396_
timestamp 1649977179
transform -1 0 8280 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1397_
timestamp 1649977179
transform 1 0 6716 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1398_
timestamp 1649977179
transform 1 0 13248 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1399_
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1400_
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1401_
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1402_
timestamp 1649977179
transform -1 0 17112 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1403_
timestamp 1649977179
transform 1 0 11960 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1404_
timestamp 1649977179
transform 1 0 15456 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1405_
timestamp 1649977179
transform 1 0 17756 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1406_
timestamp 1649977179
transform -1 0 18308 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1407_
timestamp 1649977179
transform 1 0 17388 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1408_
timestamp 1649977179
transform 1 0 17112 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1409_
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1410_
timestamp 1649977179
transform 1 0 17296 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1411_
timestamp 1649977179
transform 1 0 13156 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1412_
timestamp 1649977179
transform 1 0 14812 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1413_
timestamp 1649977179
transform -1 0 10672 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1414_
timestamp 1649977179
transform 1 0 9384 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1415_
timestamp 1649977179
transform 1 0 9108 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1416_
timestamp 1649977179
transform 1 0 10580 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1417_
timestamp 1649977179
transform -1 0 11224 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1418_
timestamp 1649977179
transform 1 0 9200 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1419_
timestamp 1649977179
transform -1 0 9844 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1420_
timestamp 1649977179
transform -1 0 11408 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1421_
timestamp 1649977179
transform -1 0 9384 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1422_
timestamp 1649977179
transform 1 0 2576 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1423_
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1424_
timestamp 1649977179
transform -1 0 3680 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1425_
timestamp 1649977179
transform 1 0 2116 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1426_
timestamp 1649977179
transform -1 0 2852 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1427_
timestamp 1649977179
transform 1 0 2116 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1428_
timestamp 1649977179
transform 1 0 4324 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1429_
timestamp 1649977179
transform 1 0 4232 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1430_
timestamp 1649977179
transform -1 0 8004 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1431_
timestamp 1649977179
transform 1 0 9752 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1432_
timestamp 1649977179
transform 1 0 6992 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1433_
timestamp 1649977179
transform -1 0 10212 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1434_
timestamp 1649977179
transform -1 0 9752 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1435_
timestamp 1649977179
transform 1 0 11040 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1436_
timestamp 1649977179
transform -1 0 12236 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1437_
timestamp 1649977179
transform -1 0 10672 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1438_
timestamp 1649977179
transform 1 0 9568 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1439_
timestamp 1649977179
transform 1 0 10212 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1440_
timestamp 1649977179
transform 1 0 9936 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1441_
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1442_
timestamp 1649977179
transform -1 0 11132 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1443_
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1444_
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1445_
timestamp 1649977179
transform 1 0 10672 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1446_
timestamp 1649977179
transform 1 0 10304 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1447_
timestamp 1649977179
transform 1 0 10120 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1448_
timestamp 1649977179
transform 1 0 10304 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1449_
timestamp 1649977179
transform -1 0 11040 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1450_
timestamp 1649977179
transform 1 0 9476 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1451_
timestamp 1649977179
transform -1 0 14352 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1452_
timestamp 1649977179
transform 1 0 14260 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1453_
timestamp 1649977179
transform 1 0 13984 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1454_
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1455_
timestamp 1649977179
transform 1 0 14904 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1456_
timestamp 1649977179
transform -1 0 15732 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1457_
timestamp 1649977179
transform 1 0 14628 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1458_
timestamp 1649977179
transform -1 0 11960 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1459_
timestamp 1649977179
transform 1 0 10304 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1460_
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1461_
timestamp 1649977179
transform 1 0 11408 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1462_
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1463_
timestamp 1649977179
transform 1 0 14444 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1464_
timestamp 1649977179
transform 1 0 12788 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1465_
timestamp 1649977179
transform -1 0 14352 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1466_
timestamp 1649977179
transform -1 0 13892 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1467_
timestamp 1649977179
transform 1 0 12788 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1468_
timestamp 1649977179
transform 1 0 12512 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1469_
timestamp 1649977179
transform 1 0 17480 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1470_
timestamp 1649977179
transform -1 0 18308 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1471_
timestamp 1649977179
transform -1 0 19688 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1472_
timestamp 1649977179
transform -1 0 18308 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1473_
timestamp 1649977179
transform -1 0 19320 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1474_
timestamp 1649977179
transform -1 0 18768 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1475_
timestamp 1649977179
transform 1 0 20884 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1476_
timestamp 1649977179
transform -1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1477_
timestamp 1649977179
transform -1 0 23276 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1478_
timestamp 1649977179
transform 1 0 21620 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1479_
timestamp 1649977179
transform -1 0 22540 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1480_
timestamp 1649977179
transform -1 0 20148 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1481_
timestamp 1649977179
transform 1 0 17480 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1482_
timestamp 1649977179
transform 1 0 18492 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1483_
timestamp 1649977179
transform 1 0 17020 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1484_
timestamp 1649977179
transform -1 0 18768 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1485_
timestamp 1649977179
transform -1 0 18584 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1486_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7636 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1487_
timestamp 1649977179
transform 1 0 12696 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1488_
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1489_
timestamp 1649977179
transform -1 0 21436 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1490_
timestamp 1649977179
transform -1 0 18768 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1491_
timestamp 1649977179
transform 1 0 20884 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1492_
timestamp 1649977179
transform 1 0 18676 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1493_
timestamp 1649977179
transform -1 0 17112 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1494_
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1495_
timestamp 1649977179
transform 1 0 14996 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1496_
timestamp 1649977179
transform -1 0 17204 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1497_
timestamp 1649977179
transform 1 0 16100 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1498_
timestamp 1649977179
transform -1 0 16008 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1499_
timestamp 1649977179
transform 1 0 14536 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1500_
timestamp 1649977179
transform 1 0 19228 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1501_
timestamp 1649977179
transform -1 0 18952 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1502_
timestamp 1649977179
transform -1 0 18860 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1503_
timestamp 1649977179
transform -1 0 18676 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1504_
timestamp 1649977179
transform 1 0 25944 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1505_
timestamp 1649977179
transform -1 0 28704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1506_
timestamp 1649977179
transform -1 0 31096 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1507_
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1508_
timestamp 1649977179
transform 1 0 30176 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1509_
timestamp 1649977179
transform -1 0 31832 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1510_
timestamp 1649977179
transform -1 0 30912 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1511_
timestamp 1649977179
transform 1 0 32200 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1512_
timestamp 1649977179
transform -1 0 31004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1513_
timestamp 1649977179
transform -1 0 28704 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1514_
timestamp 1649977179
transform 1 0 27324 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1515_
timestamp 1649977179
transform -1 0 28428 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1516_
timestamp 1649977179
transform 1 0 27232 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1517_
timestamp 1649977179
transform -1 0 20424 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1518_
timestamp 1649977179
transform 1 0 11868 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1519_
timestamp 1649977179
transform 1 0 17664 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1520_
timestamp 1649977179
transform -1 0 19596 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1521_
timestamp 1649977179
transform -1 0 18768 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1522_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7636 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1523_
timestamp 1649977179
transform -1 0 7176 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1524_
timestamp 1649977179
transform -1 0 5152 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _1525_
timestamp 1649977179
transform -1 0 7268 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1526_
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1527_
timestamp 1649977179
transform 1 0 7544 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__nor3_1  _1528_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6624 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_2  _1529_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1530_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5244 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1531_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 35788 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1532_
timestamp 1649977179
transform 1 0 22724 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1533_
timestamp 1649977179
transform 1 0 22264 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1534_
timestamp 1649977179
transform -1 0 29808 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1535_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 25024 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1536_
timestamp 1649977179
transform 1 0 4600 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1537_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1538_
timestamp 1649977179
transform 1 0 9936 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1539_
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1540_
timestamp 1649977179
transform -1 0 10488 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1541_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7176 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1542_
timestamp 1649977179
transform -1 0 35696 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1543_
timestamp 1649977179
transform 1 0 22632 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1544_
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1545_
timestamp 1649977179
transform -1 0 28796 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1546_
timestamp 1649977179
transform -1 0 23920 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1547_
timestamp 1649977179
transform 1 0 4232 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1548_
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1549_
timestamp 1649977179
transform 1 0 9844 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1550_
timestamp 1649977179
transform 1 0 10948 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1551_
timestamp 1649977179
transform -1 0 8464 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1552_
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a21bo_1  _1553_
timestamp 1649977179
transform 1 0 6348 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1554_
timestamp 1649977179
transform 1 0 6624 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1555_
timestamp 1649977179
transform -1 0 35696 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1556_
timestamp 1649977179
transform 1 0 22356 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1557_
timestamp 1649977179
transform 1 0 23092 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1558_
timestamp 1649977179
transform -1 0 28704 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1559_
timestamp 1649977179
transform -1 0 23552 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1560_
timestamp 1649977179
transform 1 0 4324 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1561_
timestamp 1649977179
transform 1 0 4968 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1562_
timestamp 1649977179
transform 1 0 11224 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1563_
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1564_
timestamp 1649977179
transform -1 0 7452 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1565_
timestamp 1649977179
transform -1 0 5888 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a21bo_1  _1566_
timestamp 1649977179
transform 1 0 5612 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1567_
timestamp 1649977179
transform 1 0 6808 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1568_
timestamp 1649977179
transform 1 0 35420 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1569_
timestamp 1649977179
transform 1 0 36156 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1570_
timestamp 1649977179
transform 1 0 35236 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1571_
timestamp 1649977179
transform 1 0 35880 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1572_
timestamp 1649977179
transform -1 0 35788 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1573_
timestamp 1649977179
transform 1 0 23644 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1574_
timestamp 1649977179
transform 1 0 29808 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1575_
timestamp 1649977179
transform 1 0 23000 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1576_
timestamp 1649977179
transform 1 0 29624 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1577_
timestamp 1649977179
transform 1 0 29532 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1578_
timestamp 1649977179
transform 1 0 21988 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1579_
timestamp 1649977179
transform 1 0 28152 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1580_
timestamp 1649977179
transform 1 0 21804 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1581_
timestamp 1649977179
transform 1 0 27968 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1582_
timestamp 1649977179
transform 1 0 27416 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1583_
timestamp 1649977179
transform 1 0 30728 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1584_
timestamp 1649977179
transform -1 0 33856 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1585_
timestamp 1649977179
transform -1 0 31648 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1586_
timestamp 1649977179
transform -1 0 33764 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1587_
timestamp 1649977179
transform -1 0 31464 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1588_
timestamp 1649977179
transform -1 0 31096 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1589_
timestamp 1649977179
transform 1 0 12880 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1590_
timestamp 1649977179
transform -1 0 13524 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1591_
timestamp 1649977179
transform 1 0 11592 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1592_
timestamp 1649977179
transform -1 0 12788 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1593_
timestamp 1649977179
transform 1 0 6532 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1594_
timestamp 1649977179
transform 1 0 6624 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1595_
timestamp 1649977179
transform 1 0 19504 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1596_
timestamp 1649977179
transform 1 0 22172 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1597_
timestamp 1649977179
transform 1 0 18216 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1598_
timestamp 1649977179
transform 1 0 22816 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1599_
timestamp 1649977179
transform -1 0 14904 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1600_
timestamp 1649977179
transform 1 0 14260 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1601_
timestamp 1649977179
transform -1 0 8740 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1602_
timestamp 1649977179
transform 1 0 4508 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1603_
timestamp 1649977179
transform -1 0 8740 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1604_
timestamp 1649977179
transform 1 0 6900 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1605_
timestamp 1649977179
transform -1 0 36524 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1606_
timestamp 1649977179
transform -1 0 31556 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1607_
timestamp 1649977179
transform 1 0 27416 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1608_
timestamp 1649977179
transform -1 0 31372 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1609_
timestamp 1649977179
transform -1 0 30176 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1610_
timestamp 1649977179
transform -1 0 14812 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1611_
timestamp 1649977179
transform -1 0 12604 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1612_
timestamp 1649977179
transform 1 0 7452 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1613_
timestamp 1649977179
transform 1 0 8372 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1614_
timestamp 1649977179
transform 1 0 21068 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1615_
timestamp 1649977179
transform 1 0 15456 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1616_
timestamp 1649977179
transform 1 0 14904 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1617_
timestamp 1649977179
transform 1 0 15364 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1618_
timestamp 1649977179
transform -1 0 9660 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1619_
timestamp 1649977179
transform 1 0 4968 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1620_
timestamp 1649977179
transform 1 0 7084 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1621_
timestamp 1649977179
transform 1 0 9292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1622_
timestamp 1649977179
transform -1 0 35788 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1623_
timestamp 1649977179
transform -1 0 34408 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1624_
timestamp 1649977179
transform 1 0 31648 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1625_
timestamp 1649977179
transform -1 0 33856 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1626_
timestamp 1649977179
transform -1 0 33580 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1627_
timestamp 1649977179
transform 1 0 11500 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1628_
timestamp 1649977179
transform 1 0 19320 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1629_
timestamp 1649977179
transform -1 0 22724 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1630_
timestamp 1649977179
transform 1 0 20792 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1631_
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1632_
timestamp 1649977179
transform 1 0 5796 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1633_
timestamp 1649977179
transform -1 0 8280 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1634_
timestamp 1649977179
transform -1 0 36340 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1635_
timestamp 1649977179
transform 1 0 31740 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1636_
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1637_
timestamp 1649977179
transform -1 0 34132 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1638_
timestamp 1649977179
transform -1 0 33580 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1639_
timestamp 1649977179
transform 1 0 16744 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1640_
timestamp 1649977179
transform 1 0 17296 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1641_
timestamp 1649977179
transform -1 0 23276 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1642_
timestamp 1649977179
transform -1 0 22632 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1643_
timestamp 1649977179
transform -1 0 20056 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1644_
timestamp 1649977179
transform 1 0 6348 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1645_
timestamp 1649977179
transform 1 0 4600 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1646_
timestamp 1649977179
transform 1 0 9200 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1647_
timestamp 1649977179
transform -1 0 36340 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1648_
timestamp 1649977179
transform 1 0 32016 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1649_
timestamp 1649977179
transform 1 0 32660 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1650_
timestamp 1649977179
transform -1 0 34132 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1651_
timestamp 1649977179
transform 1 0 34776 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1652_
timestamp 1649977179
transform 1 0 15732 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1653_
timestamp 1649977179
transform 1 0 19320 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1654_
timestamp 1649977179
transform -1 0 23460 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1655_
timestamp 1649977179
transform 1 0 22908 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1656_
timestamp 1649977179
transform -1 0 21344 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1657_
timestamp 1649977179
transform -1 0 5888 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a21bo_1  _1658_
timestamp 1649977179
transform -1 0 10948 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1659_
timestamp 1649977179
transform 1 0 10212 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1660_
timestamp 1649977179
transform -1 0 37168 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1661_
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1662_
timestamp 1649977179
transform 1 0 29256 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1663_
timestamp 1649977179
transform -1 0 35328 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1664_
timestamp 1649977179
transform -1 0 30452 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1665_
timestamp 1649977179
transform 1 0 12972 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1666_
timestamp 1649977179
transform 1 0 19320 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1667_
timestamp 1649977179
transform -1 0 23000 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1668_
timestamp 1649977179
transform 1 0 22448 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1669_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 22908 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1670_
timestamp 1649977179
transform 1 0 10120 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1671_
timestamp 1649977179
transform -1 0 12328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1672_
timestamp 1649977179
transform -1 0 37904 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1673_
timestamp 1649977179
transform 1 0 28428 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1674_
timestamp 1649977179
transform 1 0 28428 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1675_
timestamp 1649977179
transform -1 0 34776 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1676_
timestamp 1649977179
transform -1 0 31096 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1677_
timestamp 1649977179
transform 1 0 13064 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1678_
timestamp 1649977179
transform 1 0 16192 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1679_
timestamp 1649977179
transform -1 0 24564 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1680_
timestamp 1649977179
transform -1 0 20240 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1681_
timestamp 1649977179
transform -1 0 17848 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1682_
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1683_
timestamp 1649977179
transform -1 0 12052 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1684_
timestamp 1649977179
transform -1 0 37444 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1685_
timestamp 1649977179
transform 1 0 24472 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1686_
timestamp 1649977179
transform 1 0 22356 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1687_
timestamp 1649977179
transform -1 0 34224 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1688_
timestamp 1649977179
transform -1 0 25392 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1689_
timestamp 1649977179
transform 1 0 12788 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1690_
timestamp 1649977179
transform 1 0 14904 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1691_
timestamp 1649977179
transform 1 0 19872 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1692_
timestamp 1649977179
transform -1 0 20608 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1693_
timestamp 1649977179
transform -1 0 19964 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1694_
timestamp 1649977179
transform 1 0 4508 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1695_
timestamp 1649977179
transform -1 0 5520 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1696_
timestamp 1649977179
transform -1 0 36800 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1697_
timestamp 1649977179
transform 1 0 25392 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1698_
timestamp 1649977179
transform 1 0 25852 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1699_
timestamp 1649977179
transform -1 0 33212 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1700_
timestamp 1649977179
transform -1 0 27508 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1701_
timestamp 1649977179
transform 1 0 12512 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1702_
timestamp 1649977179
transform 1 0 13340 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1703_
timestamp 1649977179
transform -1 0 22448 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1704_
timestamp 1649977179
transform -1 0 20700 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1705_
timestamp 1649977179
transform -1 0 14996 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1706_
timestamp 1649977179
transform 1 0 7728 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1707_
timestamp 1649977179
transform -1 0 9752 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1708_
timestamp 1649977179
transform -1 0 5244 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1709_
timestamp 1649977179
transform -1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1710_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2760 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1711_
timestamp 1649977179
transform 1 0 2852 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1712_
timestamp 1649977179
transform 1 0 2392 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1713_
timestamp 1649977179
transform 1 0 1840 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 1649977179
transform 1 0 1840 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1716_
timestamp 1649977179
transform 1 0 2024 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1717_
timestamp 1649977179
transform 1 0 8280 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1718_
timestamp 1649977179
transform 1 0 2300 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1719_
timestamp 1649977179
transform -1 0 15548 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 1649977179
transform 1 0 2208 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1721_
timestamp 1649977179
transform 1 0 5888 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1722_
timestamp 1649977179
transform 1 0 2576 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1723_
timestamp 1649977179
transform 1 0 2392 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1724_
timestamp 1649977179
transform 1 0 1840 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1725_
timestamp 1649977179
transform 1 0 5520 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1726_
timestamp 1649977179
transform 1 0 6072 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1727_
timestamp 1649977179
transform 1 0 10672 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1728_
timestamp 1649977179
transform -1 0 18124 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1729_
timestamp 1649977179
transform 1 0 16100 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1730_
timestamp 1649977179
transform -1 0 13616 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1731_
timestamp 1649977179
transform -1 0 14260 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1732_
timestamp 1649977179
transform -1 0 13708 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1733_
timestamp 1649977179
transform 1 0 12144 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1734_
timestamp 1649977179
transform -1 0 31004 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1735_
timestamp 1649977179
transform 1 0 27416 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1736_
timestamp 1649977179
transform 1 0 26956 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1737_
timestamp 1649977179
transform 1 0 30176 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1738_
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1739_
timestamp 1649977179
transform -1 0 38732 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1740_
timestamp 1649977179
transform 1 0 37904 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1741_
timestamp 1649977179
transform 1 0 37904 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1742_
timestamp 1649977179
transform 1 0 37904 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1743_
timestamp 1649977179
transform -1 0 38824 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1744_
timestamp 1649977179
transform -1 0 36432 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1745_
timestamp 1649977179
transform 1 0 33120 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1746_
timestamp 1649977179
transform -1 0 31004 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1747_
timestamp 1649977179
transform 1 0 27324 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1748_
timestamp 1649977179
transform 1 0 27232 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1749_
timestamp 1649977179
transform 1 0 30544 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1750_
timestamp 1649977179
transform 1 0 31188 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1751_
timestamp 1649977179
transform 1 0 32292 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1752_
timestamp 1649977179
transform -1 0 35972 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1753_
timestamp 1649977179
transform -1 0 36156 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1754_
timestamp 1649977179
transform 1 0 34868 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1755_
timestamp 1649977179
transform 1 0 35604 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1756_
timestamp 1649977179
transform 1 0 32660 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1757_
timestamp 1649977179
transform -1 0 34040 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1758_
timestamp 1649977179
transform 1 0 4508 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1759_
timestamp 1649977179
transform 1 0 2576 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1760_
timestamp 1649977179
transform 1 0 2576 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1761_
timestamp 1649977179
transform 1 0 6348 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1762_
timestamp 1649977179
transform -1 0 7820 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1763_
timestamp 1649977179
transform -1 0 21896 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1764_
timestamp 1649977179
transform 1 0 18492 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1765_
timestamp 1649977179
transform 1 0 19228 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1766_
timestamp 1649977179
transform -1 0 21712 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1767_
timestamp 1649977179
transform 1 0 18676 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1768_
timestamp 1649977179
transform -1 0 16560 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1769_
timestamp 1649977179
transform -1 0 15824 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1770_
timestamp 1649977179
transform 1 0 8372 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1771_
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1772_
timestamp 1649977179
transform -1 0 12972 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1773_
timestamp 1649977179
transform 1 0 12144 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1774_
timestamp 1649977179
transform 1 0 14352 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1775_
timestamp 1649977179
transform -1 0 26588 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1776_
timestamp 1649977179
transform 1 0 24932 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1777_
timestamp 1649977179
transform 1 0 24564 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1778_
timestamp 1649977179
transform -1 0 27232 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1779_
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1780_
timestamp 1649977179
transform -1 0 26864 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1781_
timestamp 1649977179
transform -1 0 27416 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1782_
timestamp 1649977179
transform -1 0 23368 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1783_
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1784_
timestamp 1649977179
transform 1 0 22632 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1785_
timestamp 1649977179
transform 1 0 24840 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1786_
timestamp 1649977179
transform 1 0 25024 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1787_
timestamp 1649977179
transform 1 0 30176 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1788_
timestamp 1649977179
transform -1 0 34224 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1789_
timestamp 1649977179
transform -1 0 33856 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1790_
timestamp 1649977179
transform 1 0 32384 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1791_
timestamp 1649977179
transform 1 0 28244 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1792_
timestamp 1649977179
transform 1 0 21620 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1793_
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1794_
timestamp 1649977179
transform -1 0 15640 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1795_
timestamp 1649977179
transform -1 0 15456 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1796_
timestamp 1649977179
transform -1 0 14628 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1797_
timestamp 1649977179
transform -1 0 18492 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1798_
timestamp 1649977179
transform -1 0 18492 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1799_
timestamp 1649977179
transform -1 0 29624 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1800_
timestamp 1649977179
transform -1 0 32384 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1801_
timestamp 1649977179
transform -1 0 30728 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1802_
timestamp 1649977179
transform 1 0 27692 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1803_
timestamp 1649977179
transform 1 0 25576 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1804_
timestamp 1649977179
transform -1 0 21344 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1805_
timestamp 1649977179
transform -1 0 22632 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1806_
timestamp 1649977179
transform 1 0 35052 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1807_
timestamp 1649977179
transform 1 0 38272 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1808_
timestamp 1649977179
transform 1 0 37352 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1809_
timestamp 1649977179
transform -1 0 39744 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1810_
timestamp 1649977179
transform 1 0 39836 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1811_
timestamp 1649977179
transform -1 0 37628 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1812_
timestamp 1649977179
transform -1 0 40204 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1813_
timestamp 1649977179
transform -1 0 40204 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1814_
timestamp 1649977179
transform -1 0 39376 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1815_
timestamp 1649977179
transform -1 0 39376 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1816_
timestamp 1649977179
transform 1 0 38824 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1817_
timestamp 1649977179
transform 1 0 35696 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1818_
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1819_
timestamp 1649977179
transform 1 0 35144 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1820_
timestamp 1649977179
transform -1 0 36156 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1821_
timestamp 1649977179
transform -1 0 39376 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1822_
timestamp 1649977179
transform 1 0 38548 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1823_
timestamp 1649977179
transform -1 0 37444 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1649977179
transform -1 0 40204 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1649977179
transform -1 0 40204 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1649977179
transform -1 0 40020 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1649977179
transform -1 0 40388 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1828_
timestamp 1649977179
transform 1 0 38824 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1649977179
transform 1 0 36064 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1649977179
transform 1 0 26864 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1831_
timestamp 1649977179
transform -1 0 26496 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1832_
timestamp 1649977179
transform -1 0 31096 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1833_
timestamp 1649977179
transform 1 0 29624 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1834_
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1835_
timestamp 1649977179
transform 1 0 32752 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1836_
timestamp 1649977179
transform 1 0 33580 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1837_
timestamp 1649977179
transform -1 0 34224 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1838_
timestamp 1649977179
transform -1 0 35052 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1839_
timestamp 1649977179
transform -1 0 33672 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1840_
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1841_
timestamp 1649977179
transform 1 0 24564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1842_
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1843_
timestamp 1649977179
transform 1 0 2392 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1844_
timestamp 1649977179
transform 1 0 1840 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1845_
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1846_
timestamp 1649977179
transform 1 0 6440 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1847_
timestamp 1649977179
transform -1 0 22448 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1848_
timestamp 1649977179
transform -1 0 25024 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1849_
timestamp 1649977179
transform 1 0 24380 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1850_
timestamp 1649977179
transform 1 0 22080 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1851_
timestamp 1649977179
transform 1 0 22264 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1852_
timestamp 1649977179
transform 1 0 17296 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1853_
timestamp 1649977179
transform 1 0 19412 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1854_
timestamp 1649977179
transform 1 0 16836 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1855_
timestamp 1649977179
transform 1 0 18308 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1856_
timestamp 1649977179
transform 1 0 15088 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1857_
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1858_
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1859_
timestamp 1649977179
transform 1 0 25024 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1860_
timestamp 1649977179
transform 1 0 25576 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1861_
timestamp 1649977179
transform 1 0 27876 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1862_
timestamp 1649977179
transform 1 0 26404 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1863_
timestamp 1649977179
transform 1 0 25576 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1864_
timestamp 1649977179
transform 1 0 22448 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1865_
timestamp 1649977179
transform 1 0 23000 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1866_
timestamp 1649977179
transform -1 0 8280 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1867_
timestamp 1649977179
transform -1 0 3956 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1868_
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1869_
timestamp 1649977179
transform -1 0 6808 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1870_
timestamp 1649977179
transform 1 0 6624 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1871_
timestamp 1649977179
transform 1 0 13156 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1872_
timestamp 1649977179
transform 1 0 15364 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1873_
timestamp 1649977179
transform 1 0 18400 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1874_
timestamp 1649977179
transform 1 0 17112 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1875_
timestamp 1649977179
transform -1 0 16928 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1876_
timestamp 1649977179
transform -1 0 14444 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1877_
timestamp 1649977179
transform 1 0 9108 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1878_
timestamp 1649977179
transform 1 0 2392 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1879_
timestamp 1649977179
transform 1 0 1840 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1880_
timestamp 1649977179
transform 1 0 2208 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1881_
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1882_
timestamp 1649977179
transform 1 0 5612 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1883_
timestamp 1649977179
transform 1 0 7360 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1884_
timestamp 1649977179
transform 1 0 9200 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1885_
timestamp 1649977179
transform 1 0 9200 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1886_
timestamp 1649977179
transform 1 0 10580 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1887_
timestamp 1649977179
transform 1 0 10120 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1888_
timestamp 1649977179
transform 1 0 9476 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1889_
timestamp 1649977179
transform 1 0 9200 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1890_
timestamp 1649977179
transform 1 0 9568 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1891_
timestamp 1649977179
transform 1 0 9568 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1892_
timestamp 1649977179
transform -1 0 13616 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1893_
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1894_
timestamp 1649977179
transform 1 0 12236 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1895_
timestamp 1649977179
transform 1 0 18676 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1896_
timestamp 1649977179
transform 1 0 19136 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1897_
timestamp 1649977179
transform -1 0 23000 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1898_
timestamp 1649977179
transform -1 0 23828 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1899_
timestamp 1649977179
transform 1 0 16928 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1900_
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1901_
timestamp 1649977179
transform 1 0 18216 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1902_
timestamp 1649977179
transform 1 0 14720 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1903_
timestamp 1649977179
transform 1 0 16008 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1904_
timestamp 1649977179
transform 1 0 14260 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1905_
timestamp 1649977179
transform 1 0 19504 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1906_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1907_
timestamp 1649977179
transform 1 0 30176 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1908_
timestamp 1649977179
transform 1 0 30728 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1909_
timestamp 1649977179
transform 1 0 31188 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1910_
timestamp 1649977179
transform 1 0 27232 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1911_
timestamp 1649977179
transform 1 0 27140 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1912_
timestamp 1649977179
transform 1 0 17296 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1913_
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1914_
timestamp 1649977179
transform 1 0 1840 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1915_
timestamp 1649977179
transform -1 0 9108 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1916_
timestamp 1649977179
transform -1 0 8464 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1917_
timestamp 1649977179
transform -1 0 8188 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1918_
timestamp 1649977179
transform -1 0 8464 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1919_
timestamp 1649977179
transform 1 0 7084 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1920_
timestamp 1649977179
transform -1 0 10948 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1921_
timestamp 1649977179
transform 1 0 10764 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1922_
timestamp 1649977179
transform -1 0 11960 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1923_
timestamp 1649977179
transform -1 0 13064 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1924_
timestamp 1649977179
transform 1 0 4232 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1925_
timestamp 1649977179
transform 1 0 8924 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1926_
timestamp 1649977179
transform 1 0 2392 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _2176_
timestamp 1649977179
transform -1 0 46368 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2177_
timestamp 1649977179
transform -1 0 22172 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2178_
timestamp 1649977179
transform -1 0 44068 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2179_
timestamp 1649977179
transform 1 0 19964 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2180_
timestamp 1649977179
transform 1 0 18492 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2181_
timestamp 1649977179
transform 1 0 18768 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2182_
timestamp 1649977179
transform 1 0 18124 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2183_
timestamp 1649977179
transform 1 0 19412 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2184_
timestamp 1649977179
transform 1 0 20056 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2185_
timestamp 1649977179
transform -1 0 24748 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2186_
timestamp 1649977179
transform -1 0 29440 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2187_
timestamp 1649977179
transform -1 0 32384 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2188_
timestamp 1649977179
transform -1 0 31372 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2189_
timestamp 1649977179
transform -1 0 28796 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2190_
timestamp 1649977179
transform -1 0 25392 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2191_
timestamp 1649977179
transform -1 0 27232 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2192_
timestamp 1649977179
transform -1 0 26496 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2193_
timestamp 1649977179
transform -1 0 24104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2194_
timestamp 1649977179
transform -1 0 22816 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2195_
timestamp 1649977179
transform -1 0 21344 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2196_
timestamp 1649977179
transform -1 0 19596 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2197_
timestamp 1649977179
transform -1 0 18768 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2198_
timestamp 1649977179
transform 1 0 17480 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2199_
timestamp 1649977179
transform 1 0 17480 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2200_
timestamp 1649977179
transform 1 0 15732 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2201_
timestamp 1649977179
transform 1 0 13524 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2202_
timestamp 1649977179
transform 1 0 19596 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2203_
timestamp 1649977179
transform -1 0 23460 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2204_
timestamp 1649977179
transform -1 0 30728 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2205_
timestamp 1649977179
transform -1 0 35788 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20516 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1649977179
transform -1 0 12236 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1649977179
transform -1 0 9660 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1649977179
transform 1 0 31188 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1649977179
transform -1 0 30452 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_wb_clk_i
timestamp 1649977179
transform 1 0 6624 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_wb_clk_i
timestamp 1649977179
transform -1 0 4508 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_wb_clk_i
timestamp 1649977179
transform 1 0 10580 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_wb_clk_i
timestamp 1649977179
transform -1 0 16836 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_wb_clk_i
timestamp 1649977179
transform 1 0 9292 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_wb_clk_i
timestamp 1649977179
transform 1 0 4140 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_wb_clk_i
timestamp 1649977179
transform 1 0 5888 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_wb_clk_i
timestamp 1649977179
transform -1 0 4968 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_wb_clk_i
timestamp 1649977179
transform 1 0 9292 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_wb_clk_i
timestamp 1649977179
transform 1 0 17020 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_wb_clk_i
timestamp 1649977179
transform 1 0 16744 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_wb_clk_i
timestamp 1649977179
transform -1 0 22816 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_12_wb_clk_i
timestamp 1649977179
transform 1 0 27232 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_13_wb_clk_i
timestamp 1649977179
transform 1 0 23644 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_14_wb_clk_i
timestamp 1649977179
transform 1 0 27784 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_15_wb_clk_i
timestamp 1649977179
transform 1 0 32384 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_16_wb_clk_i
timestamp 1649977179
transform 1 0 37628 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_17_wb_clk_i
timestamp 1649977179
transform 1 0 38272 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_18_wb_clk_i
timestamp 1649977179
transform 1 0 31004 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_19_wb_clk_i
timestamp 1649977179
transform -1 0 26496 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_20_wb_clk_i
timestamp 1649977179
transform 1 0 32476 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_21_wb_clk_i
timestamp 1649977179
transform 1 0 37996 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_22_wb_clk_i
timestamp 1649977179
transform 1 0 37628 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_23_wb_clk_i
timestamp 1649977179
transform 1 0 37628 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_24_wb_clk_i
timestamp 1649977179
transform 1 0 37076 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_25_wb_clk_i
timestamp 1649977179
transform 1 0 29992 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_26_wb_clk_i
timestamp 1649977179
transform -1 0 26036 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_27_wb_clk_i
timestamp 1649977179
transform 1 0 24288 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_28_wb_clk_i
timestamp 1649977179
transform 1 0 16928 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_29_wb_clk_i
timestamp 1649977179
transform 1 0 17296 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_30_wb_clk_i
timestamp 1649977179
transform 1 0 14352 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_31_wb_clk_i
timestamp 1649977179
transform -1 0 5980 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1649977179
transform 1 0 13248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1649977179
transform 1 0 15824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1649977179
transform 1 0 18400 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1649977179
transform -1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1649977179
transform -1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1649977179
transform -1 0 19136 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1649977179
transform -1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1649977179
transform -1 0 19872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1649977179
transform 1 0 20056 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1649977179
transform 1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1649977179
transform -1 0 20608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1649977179
transform 1 0 15640 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1649977179
transform -1 0 21252 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1649977179
transform -1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1649977179
transform -1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1649977179
transform -1 0 22080 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1649977179
transform 1 0 20976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1649977179
transform 1 0 22080 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1649977179
transform -1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1649977179
transform 1 0 22816 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1649977179
transform -1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1649977179
transform 1 0 23368 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1649977179
transform 1 0 14352 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input24
timestamp 1649977179
transform 1 0 14352 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1649977179
transform -1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1649977179
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input27
timestamp 1649977179
transform -1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input28
timestamp 1649977179
transform 1 0 17296 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input30
timestamp 1649977179
transform -1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1649977179
transform 1 0 6532 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform -1 0 13616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform -1 0 12328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1649977179
transform 1 0 6716 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform -1 0 14536 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform -1 0 13616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1649977179
transform 1 0 7268 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform 1 0 7268 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform -1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform -1 0 1840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform 1 0 5612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1649977179
transform -1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1649977179
transform -1 0 9752 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1649977179
transform -1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1649977179
transform 1 0 1656 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1649977179
transform -1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input50
timestamp 1649977179
transform 1 0 7544 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1649977179
transform -1 0 5060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input52
timestamp 1649977179
transform -1 0 6900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input53
timestamp 1649977179
transform -1 0 9844 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input54
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input55
timestamp 1649977179
transform 1 0 9384 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input56
timestamp 1649977179
transform 1 0 10304 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform -1 0 2668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1649977179
transform -1 0 4140 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1649977179
transform -1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform 1 0 47564 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform 1 0 40940 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform 1 0 45632 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform -1 0 10028 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform -1 0 8464 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform -1 0 6900 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform -1 0 5336 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform -1 0 4140 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform -1 0 2208 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform 1 0 37812 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform 1 0 36248 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform 1 0 34684 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform 1 0 33120 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform 1 0 32108 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform 1 0 29992 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform 1 0 28428 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform 1 0 26956 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform 1 0 25300 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform 1 0 24380 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform 1 0 22172 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform 1 0 20608 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform 1 0 19228 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform 1 0 17480 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform -1 0 17020 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform -1 0 14720 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform -1 0 13156 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform -1 0 11868 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform 1 0 42504 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 44068 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform 1 0 39836 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform 1 0 5520 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform 1 0 4784 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform 1 0 11316 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform -1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform -1 0 5612 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform -1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 9292 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform 1 0 12236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform -1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform -1 0 10948 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_103 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 1656 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_104
timestamp 1649977179
transform -1 0 1656 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_105
timestamp 1649977179
transform -1 0 1656 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_106
timestamp 1649977179
transform -1 0 1656 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_107
timestamp 1649977179
transform -1 0 1656 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_108
timestamp 1649977179
transform -1 0 1656 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_109
timestamp 1649977179
transform -1 0 1656 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_110
timestamp 1649977179
transform -1 0 1656 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_111
timestamp 1649977179
transform -1 0 1656 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_112
timestamp 1649977179
transform -1 0 58236 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_113
timestamp 1649977179
transform -1 0 56856 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_114
timestamp 1649977179
transform -1 0 55568 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_115
timestamp 1649977179
transform -1 0 53728 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_116
timestamp 1649977179
transform -1 0 52164 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_117
timestamp 1649977179
transform -1 0 49036 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_118
timestamp 1649977179
transform -1 0 50600 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_119
timestamp 1649977179
transform 1 0 57960 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_120
timestamp 1649977179
transform 1 0 57960 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_121
timestamp 1649977179
transform 1 0 57316 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_122
timestamp 1649977179
transform 1 0 57960 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_123
timestamp 1649977179
transform -1 0 52992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_124
timestamp 1649977179
transform -1 0 53636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_125
timestamp 1649977179
transform -1 0 51428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_126
timestamp 1649977179
transform -1 0 52440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_127
timestamp 1649977179
transform -1 0 54280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_128
timestamp 1649977179
transform -1 0 52072 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_129
timestamp 1649977179
transform -1 0 53084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_130
timestamp 1649977179
transform -1 0 53636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_131
timestamp 1649977179
transform -1 0 53728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_132
timestamp 1649977179
transform -1 0 54280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_133
timestamp 1649977179
transform -1 0 52992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_134
timestamp 1649977179
transform -1 0 54924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_135
timestamp 1649977179
transform -1 0 55568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_136
timestamp 1649977179
transform -1 0 52440 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_137
timestamp 1649977179
transform -1 0 53084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_138
timestamp 1649977179
transform -1 0 54372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_139
timestamp 1649977179
transform -1 0 56212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_140
timestamp 1649977179
transform -1 0 53636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_141
timestamp 1649977179
transform -1 0 55568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_142
timestamp 1649977179
transform -1 0 53728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_143
timestamp 1649977179
transform -1 0 54280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_144
timestamp 1649977179
transform -1 0 54924 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_145
timestamp 1649977179
transform -1 0 56856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_146
timestamp 1649977179
transform -1 0 55568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_147
timestamp 1649977179
transform -1 0 56212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_148
timestamp 1649977179
transform -1 0 54372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_149
timestamp 1649977179
transform -1 0 56212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_150
timestamp 1649977179
transform -1 0 56856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_151
timestamp 1649977179
transform -1 0 55568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_152
timestamp 1649977179
transform -1 0 58144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_153
timestamp 1649977179
transform -1 0 54004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_154
timestamp 1649977179
transform -1 0 54648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_155
timestamp 1649977179
transform -1 0 56856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_156
timestamp 1649977179
transform -1 0 55568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_157
timestamp 1649977179
transform -1 0 56212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_158
timestamp 1649977179
transform -1 0 55292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_159
timestamp 1649977179
transform -1 0 58144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_160
timestamp 1649977179
transform -1 0 56212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_161
timestamp 1649977179
transform 1 0 57960 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_162
timestamp 1649977179
transform 1 0 57316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_163
timestamp 1649977179
transform 1 0 57960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_164
timestamp 1649977179
transform 1 0 57960 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_165
timestamp 1649977179
transform 1 0 57960 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_166
timestamp 1649977179
transform 1 0 57960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_167
timestamp 1649977179
transform 1 0 57960 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_168
timestamp 1649977179
transform 1 0 57960 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_169
timestamp 1649977179
transform 1 0 57960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_170
timestamp 1649977179
transform 1 0 57960 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_171
timestamp 1649977179
transform 1 0 57960 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_172
timestamp 1649977179
transform 1 0 57960 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_173
timestamp 1649977179
transform 1 0 57960 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_174
timestamp 1649977179
transform 1 0 57960 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_175
timestamp 1649977179
transform 1 0 57960 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_176
timestamp 1649977179
transform 1 0 57960 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_177
timestamp 1649977179
transform 1 0 57960 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_178
timestamp 1649977179
transform 1 0 57960 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_179
timestamp 1649977179
transform 1 0 57960 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_180
timestamp 1649977179
transform 1 0 57960 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_181
timestamp 1649977179
transform 1 0 57960 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_182
timestamp 1649977179
transform 1 0 57960 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_183
timestamp 1649977179
transform 1 0 57960 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_184
timestamp 1649977179
transform 1 0 57960 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_185
timestamp 1649977179
transform 1 0 57960 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_186
timestamp 1649977179
transform 1 0 57960 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_187
timestamp 1649977179
transform 1 0 57960 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_188
timestamp 1649977179
transform 1 0 57960 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_189
timestamp 1649977179
transform 1 0 57960 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_190
timestamp 1649977179
transform 1 0 57960 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_191
timestamp 1649977179
transform 1 0 57960 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_192
timestamp 1649977179
transform 1 0 57960 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_193
timestamp 1649977179
transform 1 0 57960 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_194
timestamp 1649977179
transform 1 0 57960 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_195
timestamp 1649977179
transform 1 0 57960 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_196
timestamp 1649977179
transform 1 0 57960 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_197
timestamp 1649977179
transform 1 0 57960 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_198
timestamp 1649977179
transform 1 0 57960 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_199
timestamp 1649977179
transform -1 0 51704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_200
timestamp 1649977179
transform -1 0 51796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_201
timestamp 1649977179
transform -1 0 52992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_202
timestamp 1649977179
transform -1 0 15916 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_203
timestamp 1649977179
transform 1 0 13064 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_204
timestamp 1649977179
transform 1 0 14904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_205
timestamp 1649977179
transform 1 0 14996 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_206
timestamp 1649977179
transform 1 0 15548 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_207
timestamp 1649977179
transform -1 0 17112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_208
timestamp 1649977179
transform 1 0 12696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_209
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_210
timestamp 1649977179
transform -1 0 17848 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_211
timestamp 1649977179
transform 1 0 14352 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_212
timestamp 1649977179
transform 1 0 16192 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_213
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_214
timestamp 1649977179
transform 1 0 17848 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_215
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_216
timestamp 1649977179
transform -1 0 19596 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_217
timestamp 1649977179
transform 1 0 15364 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_218
timestamp 1649977179
transform 1 0 18492 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_219
timestamp 1649977179
transform -1 0 20424 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_220
timestamp 1649977179
transform 1 0 19136 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_221
timestamp 1649977179
transform 1 0 19780 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_222
timestamp 1649977179
transform -1 0 21252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_223
timestamp 1649977179
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_224
timestamp 1649977179
transform 1 0 20424 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_225
timestamp 1649977179
transform 1 0 21528 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_226
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_227
timestamp 1649977179
transform -1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_228
timestamp 1649977179
transform 1 0 22172 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_229
timestamp 1649977179
transform 1 0 21988 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_230
timestamp 1649977179
transform 1 0 22816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_231
timestamp 1649977179
transform -1 0 23736 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_232
timestamp 1649977179
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_233
timestamp 1649977179
transform -1 0 24748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_234
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_235
timestamp 1649977179
transform 1 0 23644 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_236
timestamp 1649977179
transform -1 0 25116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_237
timestamp 1649977179
transform 1 0 24288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_238
timestamp 1649977179
transform 1 0 24932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_239
timestamp 1649977179
transform -1 0 25944 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_240
timestamp 1649977179
transform 1 0 24932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_241
timestamp 1649977179
transform 1 0 25576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_242
timestamp 1649977179
transform 1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_243
timestamp 1649977179
transform -1 0 27048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_244
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_245
timestamp 1649977179
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_246
timestamp 1649977179
transform -1 0 27876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_247
timestamp 1649977179
transform 1 0 27416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_248
timestamp 1649977179
transform -1 0 28336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_249
timestamp 1649977179
transform 1 0 27508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_250
timestamp 1649977179
transform -1 0 28980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_251
timestamp 1649977179
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_252
timestamp 1649977179
transform 1 0 28704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_253
timestamp 1649977179
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_254
timestamp 1649977179
transform 1 0 29348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_255
timestamp 1649977179
transform -1 0 30268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_256
timestamp 1649977179
transform 1 0 29900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_257
timestamp 1649977179
transform -1 0 30912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_258
timestamp 1649977179
transform 1 0 30544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_259
timestamp 1649977179
transform -1 0 31464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_260
timestamp 1649977179
transform -1 0 32384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_261
timestamp 1649977179
transform -1 0 32384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_262
timestamp 1649977179
transform -1 0 33028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_263
timestamp 1649977179
transform -1 0 33028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_264
timestamp 1649977179
transform -1 0 33672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_265
timestamp 1649977179
transform -1 0 33672 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_266
timestamp 1649977179
transform -1 0 34960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_267
timestamp 1649977179
transform -1 0 34316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_268
timestamp 1649977179
transform -1 0 35604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_269
timestamp 1649977179
transform -1 0 34960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_270
timestamp 1649977179
transform -1 0 36248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_271
timestamp 1649977179
transform -1 0 35604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_272
timestamp 1649977179
transform -1 0 35052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_273
timestamp 1649977179
transform -1 0 35696 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_274
timestamp 1649977179
transform -1 0 36248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_275
timestamp 1649977179
transform -1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_276
timestamp 1649977179
transform -1 0 36340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_277
timestamp 1649977179
transform -1 0 38180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_278
timestamp 1649977179
transform -1 0 37536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_279
timestamp 1649977179
transform -1 0 36984 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_280
timestamp 1649977179
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_281
timestamp 1649977179
transform -1 0 38180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_282
timestamp 1649977179
transform -1 0 37812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_283
timestamp 1649977179
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_284
timestamp 1649977179
transform -1 0 40112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_285
timestamp 1649977179
transform -1 0 39468 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_286
timestamp 1649977179
transform -1 0 38916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_287
timestamp 1649977179
transform -1 0 40756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_288
timestamp 1649977179
transform -1 0 40112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_289
timestamp 1649977179
transform -1 0 41400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_290
timestamp 1649977179
transform -1 0 40756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_291
timestamp 1649977179
transform -1 0 40296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_292
timestamp 1649977179
transform -1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_293
timestamp 1649977179
transform -1 0 40940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_294
timestamp 1649977179
transform -1 0 42688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_295
timestamp 1649977179
transform -1 0 41584 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_296
timestamp 1649977179
transform -1 0 43332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_297
timestamp 1649977179
transform -1 0 42688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_298
timestamp 1649977179
transform -1 0 43976 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_299
timestamp 1649977179
transform -1 0 43332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_300
timestamp 1649977179
transform -1 0 42780 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_301
timestamp 1649977179
transform -1 0 43424 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_302
timestamp 1649977179
transform -1 0 43976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_303
timestamp 1649977179
transform -1 0 45264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_304
timestamp 1649977179
transform -1 0 44620 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_305
timestamp 1649977179
transform -1 0 45908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_306
timestamp 1649977179
transform -1 0 45264 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_307
timestamp 1649977179
transform -1 0 45264 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_308
timestamp 1649977179
transform -1 0 46552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_309
timestamp 1649977179
transform -1 0 45908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_310
timestamp 1649977179
transform -1 0 45908 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_311
timestamp 1649977179
transform -1 0 46552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_312
timestamp 1649977179
transform -1 0 47840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_313
timestamp 1649977179
transform -1 0 46552 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_314
timestamp 1649977179
transform -1 0 47196 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_315
timestamp 1649977179
transform -1 0 48484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_316
timestamp 1649977179
transform -1 0 47840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_317
timestamp 1649977179
transform -1 0 49128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_318
timestamp 1649977179
transform -1 0 48484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_319
timestamp 1649977179
transform -1 0 48024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_320
timestamp 1649977179
transform -1 0 49128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_321
timestamp 1649977179
transform -1 0 48668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_322
timestamp 1649977179
transform -1 0 50416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_323
timestamp 1649977179
transform -1 0 49772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_324
timestamp 1649977179
transform -1 0 51060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_325
timestamp 1649977179
transform -1 0 50416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_326
timestamp 1649977179
transform -1 0 51704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_327
timestamp 1649977179
transform -1 0 51060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_328
timestamp 1649977179
transform -1 0 50508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_329
timestamp 1649977179
transform -1 0 51152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_330
timestamp 1649977179
transform 1 0 57960 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_331
timestamp 1649977179
transform 1 0 57960 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_332
timestamp 1649977179
transform 1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_333
timestamp 1649977179
transform 1 0 9568 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_334
timestamp 1649977179
transform -1 0 11040 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_335
timestamp 1649977179
transform 1 0 10212 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_336
timestamp 1649977179
transform 1 0 10120 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_337
timestamp 1649977179
transform 1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_338
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_339
timestamp 1649977179
transform 1 0 11500 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_340
timestamp 1649977179
transform -1 0 12512 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_341
timestamp 1649977179
transform 1 0 12144 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_342
timestamp 1649977179
transform -1 0 13064 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_343
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_344
timestamp 1649977179
transform 1 0 12696 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_345
timestamp 1649977179
transform 1 0 13248 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_346
timestamp 1649977179
transform 1 0 11592 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_347
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_348
timestamp 1649977179
transform 1 0 13892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_349
timestamp 1649977179
transform 1 0 13064 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_350
timestamp 1649977179
transform 1 0 12420 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_351
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 314 592
<< labels >>
flabel metal2 s 47122 59200 47178 60000 0 FreeSans 224 90 0 0 CMP_out_c
port 0 nsew signal tristate
flabel metal2 s 40866 59200 40922 60000 0 FreeSans 224 90 0 0 OTA_out_c
port 1 nsew signal tristate
flabel metal2 s 45558 59200 45614 60000 0 FreeSans 224 90 0 0 OTA_sh_c
port 2 nsew signal tristate
flabel metal2 s 9586 59200 9642 60000 0 FreeSans 224 90 0 0 Pd10_a
port 3 nsew signal tristate
flabel metal2 s 8022 59200 8078 60000 0 FreeSans 224 90 0 0 Pd10_b
port 4 nsew signal tristate
flabel metal2 s 6458 59200 6514 60000 0 FreeSans 224 90 0 0 Pd11_a
port 5 nsew signal tristate
flabel metal2 s 4894 59200 4950 60000 0 FreeSans 224 90 0 0 Pd11_b
port 6 nsew signal tristate
flabel metal2 s 3330 59200 3386 60000 0 FreeSans 224 90 0 0 Pd12_a
port 7 nsew signal tristate
flabel metal2 s 1766 59200 1822 60000 0 FreeSans 224 90 0 0 Pd12_b
port 8 nsew signal tristate
flabel metal2 s 37738 59200 37794 60000 0 FreeSans 224 90 0 0 Pd1_a
port 9 nsew signal tristate
flabel metal2 s 36174 59200 36230 60000 0 FreeSans 224 90 0 0 Pd1_b
port 10 nsew signal tristate
flabel metal2 s 34610 59200 34666 60000 0 FreeSans 224 90 0 0 Pd2_a
port 11 nsew signal tristate
flabel metal2 s 33046 59200 33102 60000 0 FreeSans 224 90 0 0 Pd2_b
port 12 nsew signal tristate
flabel metal2 s 31482 59200 31538 60000 0 FreeSans 224 90 0 0 Pd3_a
port 13 nsew signal tristate
flabel metal2 s 29918 59200 29974 60000 0 FreeSans 224 90 0 0 Pd3_b
port 14 nsew signal tristate
flabel metal2 s 28354 59200 28410 60000 0 FreeSans 224 90 0 0 Pd4_a
port 15 nsew signal tristate
flabel metal2 s 26790 59200 26846 60000 0 FreeSans 224 90 0 0 Pd4_b
port 16 nsew signal tristate
flabel metal2 s 25226 59200 25282 60000 0 FreeSans 224 90 0 0 Pd5_a
port 17 nsew signal tristate
flabel metal2 s 23662 59200 23718 60000 0 FreeSans 224 90 0 0 Pd5_b
port 18 nsew signal tristate
flabel metal2 s 22098 59200 22154 60000 0 FreeSans 224 90 0 0 Pd6_a
port 19 nsew signal tristate
flabel metal2 s 20534 59200 20590 60000 0 FreeSans 224 90 0 0 Pd6_b
port 20 nsew signal tristate
flabel metal2 s 18970 59200 19026 60000 0 FreeSans 224 90 0 0 Pd7_a
port 21 nsew signal tristate
flabel metal2 s 17406 59200 17462 60000 0 FreeSans 224 90 0 0 Pd7_b
port 22 nsew signal tristate
flabel metal2 s 15842 59200 15898 60000 0 FreeSans 224 90 0 0 Pd8_a
port 23 nsew signal tristate
flabel metal2 s 14278 59200 14334 60000 0 FreeSans 224 90 0 0 Pd8_b
port 24 nsew signal tristate
flabel metal2 s 12714 59200 12770 60000 0 FreeSans 224 90 0 0 Pd9_a
port 25 nsew signal tristate
flabel metal2 s 11150 59200 11206 60000 0 FreeSans 224 90 0 0 Pd9_b
port 26 nsew signal tristate
flabel metal3 s 0 56584 800 56704 0 FreeSans 480 0 0 0 Pxl_done_i
port 27 nsew signal tristate
flabel metal3 s 0 50056 800 50176 0 FreeSans 480 0 0 0 Q1_1
port 28 nsew signal tristate
flabel metal3 s 0 48968 800 49088 0 FreeSans 480 0 0 0 Q1_2
port 29 nsew signal tristate
flabel metal3 s 0 47880 800 48000 0 FreeSans 480 0 0 0 Q1_3
port 30 nsew signal tristate
flabel metal3 s 0 52232 800 52352 0 FreeSans 480 0 0 0 Q2_1
port 31 nsew signal tristate
flabel metal3 s 0 51144 800 51264 0 FreeSans 480 0 0 0 Q2_3
port 32 nsew signal tristate
flabel metal3 s 0 55496 800 55616 0 FreeSans 480 0 0 0 Q3_1
port 33 nsew signal tristate
flabel metal3 s 0 54408 800 54528 0 FreeSans 480 0 0 0 Q3_2
port 34 nsew signal tristate
flabel metal3 s 0 53320 800 53440 0 FreeSans 480 0 0 0 Q3_3
port 35 nsew signal tristate
flabel metal2 s 42430 59200 42486 60000 0 FreeSans 224 90 0 0 SH_out_c
port 36 nsew signal tristate
flabel metal2 s 58070 59200 58126 60000 0 FreeSans 224 90 0 0 Sh
port 37 nsew signal tristate
flabel metal2 s 56506 59200 56562 60000 0 FreeSans 224 90 0 0 Sh_cmp
port 38 nsew signal tristate
flabel metal2 s 54942 59200 54998 60000 0 FreeSans 224 90 0 0 Sh_rst
port 39 nsew signal tristate
flabel metal2 s 53378 59200 53434 60000 0 FreeSans 224 90 0 0 Sw1
port 40 nsew signal tristate
flabel metal2 s 51814 59200 51870 60000 0 FreeSans 224 90 0 0 Sw2
port 41 nsew signal tristate
flabel metal2 s 48686 59200 48742 60000 0 FreeSans 224 90 0 0 Vd1
port 42 nsew signal tristate
flabel metal2 s 50250 59200 50306 60000 0 FreeSans 224 90 0 0 Vd2
port 43 nsew signal tristate
flabel metal2 s 43994 59200 44050 60000 0 FreeSans 224 90 0 0 Vref_cmp_c
port 44 nsew signal tristate
flabel metal2 s 39302 59200 39358 60000 0 FreeSans 224 90 0 0 Vref_sel_c
port 45 nsew signal tristate
flabel metal3 s 59200 52368 60000 52488 0 FreeSans 480 0 0 0 clk_o
port 46 nsew signal tristate
flabel metal3 s 59200 59168 60000 59288 0 FreeSans 480 0 0 0 counter_rst
port 47 nsew signal tristate
flabel metal3 s 59200 57808 60000 57928 0 FreeSans 480 0 0 0 data_o
port 48 nsew signal tristate
flabel metal3 s 59200 55088 60000 55208 0 FreeSans 480 0 0 0 done_o
port 49 nsew signal tristate
flabel metal3 s 0 44616 800 44736 0 FreeSans 480 0 0 0 ext_clk
port 50 nsew signal input
flabel metal3 s 0 46792 800 46912 0 FreeSans 480 0 0 0 ext_reset
port 51 nsew signal input
flabel metal3 s 0 45704 800 45824 0 FreeSans 480 0 0 0 ext_start
port 52 nsew signal input
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 io_in[0]
port 53 nsew signal input
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 io_in[10]
port 54 nsew signal input
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 io_in[11]
port 55 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 io_in[12]
port 56 nsew signal input
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 io_in[13]
port 57 nsew signal input
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 io_in[14]
port 58 nsew signal input
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 io_in[15]
port 59 nsew signal input
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 io_in[16]
port 60 nsew signal input
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 io_in[17]
port 61 nsew signal input
flabel metal3 s 0 22856 800 22976 0 FreeSans 480 0 0 0 io_in[18]
port 62 nsew signal input
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 io_in[19]
port 63 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 io_in[1]
port 64 nsew signal input
flabel metal3 s 0 25032 800 25152 0 FreeSans 480 0 0 0 io_in[20]
port 65 nsew signal input
flabel metal3 s 0 26120 800 26240 0 FreeSans 480 0 0 0 io_in[21]
port 66 nsew signal input
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 io_in[22]
port 67 nsew signal input
flabel metal3 s 0 28296 800 28416 0 FreeSans 480 0 0 0 io_in[23]
port 68 nsew signal input
flabel metal3 s 0 29384 800 29504 0 FreeSans 480 0 0 0 io_in[24]
port 69 nsew signal input
flabel metal3 s 0 30472 800 30592 0 FreeSans 480 0 0 0 io_in[25]
port 70 nsew signal input
flabel metal3 s 0 31560 800 31680 0 FreeSans 480 0 0 0 io_in[26]
port 71 nsew signal input
flabel metal3 s 0 32648 800 32768 0 FreeSans 480 0 0 0 io_in[27]
port 72 nsew signal input
flabel metal3 s 0 33736 800 33856 0 FreeSans 480 0 0 0 io_in[28]
port 73 nsew signal input
flabel metal3 s 0 34824 800 34944 0 FreeSans 480 0 0 0 io_in[29]
port 74 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 0 35912 800 36032 0 FreeSans 480 0 0 0 io_in[30]
port 76 nsew signal input
flabel metal3 s 0 37000 800 37120 0 FreeSans 480 0 0 0 io_in[31]
port 77 nsew signal input
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 io_in[32]
port 78 nsew signal input
flabel metal3 s 0 39176 800 39296 0 FreeSans 480 0 0 0 io_in[33]
port 79 nsew signal input
flabel metal3 s 0 40264 800 40384 0 FreeSans 480 0 0 0 io_in[34]
port 80 nsew signal input
flabel metal3 s 0 41352 800 41472 0 FreeSans 480 0 0 0 io_in[35]
port 81 nsew signal input
flabel metal3 s 0 42440 800 42560 0 FreeSans 480 0 0 0 io_in[36]
port 82 nsew signal input
flabel metal3 s 0 43528 800 43648 0 FreeSans 480 0 0 0 io_in[37]
port 83 nsew signal input
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 io_in[3]
port 84 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 io_in[4]
port 85 nsew signal input
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 io_in[5]
port 86 nsew signal input
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 io_in[6]
port 87 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 io_in[7]
port 88 nsew signal input
flabel metal3 s 0 11976 800 12096 0 FreeSans 480 0 0 0 io_in[8]
port 89 nsew signal input
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 io_in[9]
port 90 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 91 nsew signal tristate
flabel metal2 s 51814 0 51870 800 0 FreeSans 224 90 0 0 io_oeb[10]
port 92 nsew signal tristate
flabel metal2 s 51906 0 51962 800 0 FreeSans 224 90 0 0 io_oeb[11]
port 93 nsew signal tristate
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 io_oeb[12]
port 94 nsew signal tristate
flabel metal2 s 52090 0 52146 800 0 FreeSans 224 90 0 0 io_oeb[13]
port 95 nsew signal tristate
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 io_oeb[14]
port 96 nsew signal tristate
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 io_oeb[15]
port 97 nsew signal tristate
flabel metal2 s 52366 0 52422 800 0 FreeSans 224 90 0 0 io_oeb[16]
port 98 nsew signal tristate
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 io_oeb[17]
port 99 nsew signal tristate
flabel metal2 s 52550 0 52606 800 0 FreeSans 224 90 0 0 io_oeb[18]
port 100 nsew signal tristate
flabel metal2 s 52642 0 52698 800 0 FreeSans 224 90 0 0 io_oeb[19]
port 101 nsew signal tristate
flabel metal2 s 50986 0 51042 800 0 FreeSans 224 90 0 0 io_oeb[1]
port 102 nsew signal tristate
flabel metal2 s 52734 0 52790 800 0 FreeSans 224 90 0 0 io_oeb[20]
port 103 nsew signal tristate
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 io_oeb[21]
port 104 nsew signal tristate
flabel metal2 s 52918 0 52974 800 0 FreeSans 224 90 0 0 io_oeb[22]
port 105 nsew signal tristate
flabel metal2 s 53010 0 53066 800 0 FreeSans 224 90 0 0 io_oeb[23]
port 106 nsew signal tristate
flabel metal2 s 53102 0 53158 800 0 FreeSans 224 90 0 0 io_oeb[24]
port 107 nsew signal tristate
flabel metal2 s 53194 0 53250 800 0 FreeSans 224 90 0 0 io_oeb[25]
port 108 nsew signal tristate
flabel metal2 s 53286 0 53342 800 0 FreeSans 224 90 0 0 io_oeb[26]
port 109 nsew signal tristate
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 io_oeb[27]
port 110 nsew signal tristate
flabel metal2 s 53470 0 53526 800 0 FreeSans 224 90 0 0 io_oeb[28]
port 111 nsew signal tristate
flabel metal2 s 53562 0 53618 800 0 FreeSans 224 90 0 0 io_oeb[29]
port 112 nsew signal tristate
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 io_oeb[2]
port 113 nsew signal tristate
flabel metal2 s 53654 0 53710 800 0 FreeSans 224 90 0 0 io_oeb[30]
port 114 nsew signal tristate
flabel metal2 s 53746 0 53802 800 0 FreeSans 224 90 0 0 io_oeb[31]
port 115 nsew signal tristate
flabel metal2 s 53838 0 53894 800 0 FreeSans 224 90 0 0 io_oeb[32]
port 116 nsew signal tristate
flabel metal2 s 53930 0 53986 800 0 FreeSans 224 90 0 0 io_oeb[33]
port 117 nsew signal tristate
flabel metal2 s 54022 0 54078 800 0 FreeSans 224 90 0 0 io_oeb[34]
port 118 nsew signal tristate
flabel metal2 s 54114 0 54170 800 0 FreeSans 224 90 0 0 io_oeb[35]
port 119 nsew signal tristate
flabel metal2 s 54206 0 54262 800 0 FreeSans 224 90 0 0 io_oeb[36]
port 120 nsew signal tristate
flabel metal2 s 54298 0 54354 800 0 FreeSans 224 90 0 0 io_oeb[37]
port 121 nsew signal tristate
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 io_oeb[3]
port 122 nsew signal tristate
flabel metal2 s 51262 0 51318 800 0 FreeSans 224 90 0 0 io_oeb[4]
port 123 nsew signal tristate
flabel metal2 s 51354 0 51410 800 0 FreeSans 224 90 0 0 io_oeb[5]
port 124 nsew signal tristate
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 125 nsew signal tristate
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 io_oeb[7]
port 126 nsew signal tristate
flabel metal2 s 51630 0 51686 800 0 FreeSans 224 90 0 0 io_oeb[8]
port 127 nsew signal tristate
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 io_oeb[9]
port 128 nsew signal tristate
flabel metal3 s 59200 688 60000 808 0 FreeSans 480 0 0 0 io_out[0]
port 129 nsew signal tristate
flabel metal3 s 59200 14288 60000 14408 0 FreeSans 480 0 0 0 io_out[10]
port 130 nsew signal tristate
flabel metal3 s 59200 15648 60000 15768 0 FreeSans 480 0 0 0 io_out[11]
port 131 nsew signal tristate
flabel metal3 s 59200 17008 60000 17128 0 FreeSans 480 0 0 0 io_out[12]
port 132 nsew signal tristate
flabel metal3 s 59200 18368 60000 18488 0 FreeSans 480 0 0 0 io_out[13]
port 133 nsew signal tristate
flabel metal3 s 59200 19728 60000 19848 0 FreeSans 480 0 0 0 io_out[14]
port 134 nsew signal tristate
flabel metal3 s 59200 21088 60000 21208 0 FreeSans 480 0 0 0 io_out[15]
port 135 nsew signal tristate
flabel metal3 s 59200 22448 60000 22568 0 FreeSans 480 0 0 0 io_out[16]
port 136 nsew signal tristate
flabel metal3 s 59200 23808 60000 23928 0 FreeSans 480 0 0 0 io_out[17]
port 137 nsew signal tristate
flabel metal3 s 59200 25168 60000 25288 0 FreeSans 480 0 0 0 io_out[18]
port 138 nsew signal tristate
flabel metal3 s 59200 26528 60000 26648 0 FreeSans 480 0 0 0 io_out[19]
port 139 nsew signal tristate
flabel metal3 s 59200 2048 60000 2168 0 FreeSans 480 0 0 0 io_out[1]
port 140 nsew signal tristate
flabel metal3 s 59200 27888 60000 28008 0 FreeSans 480 0 0 0 io_out[20]
port 141 nsew signal tristate
flabel metal3 s 59200 29248 60000 29368 0 FreeSans 480 0 0 0 io_out[21]
port 142 nsew signal tristate
flabel metal3 s 59200 30608 60000 30728 0 FreeSans 480 0 0 0 io_out[22]
port 143 nsew signal tristate
flabel metal3 s 59200 31968 60000 32088 0 FreeSans 480 0 0 0 io_out[23]
port 144 nsew signal tristate
flabel metal3 s 59200 33328 60000 33448 0 FreeSans 480 0 0 0 io_out[24]
port 145 nsew signal tristate
flabel metal3 s 59200 34688 60000 34808 0 FreeSans 480 0 0 0 io_out[25]
port 146 nsew signal tristate
flabel metal3 s 59200 36048 60000 36168 0 FreeSans 480 0 0 0 io_out[26]
port 147 nsew signal tristate
flabel metal3 s 59200 37408 60000 37528 0 FreeSans 480 0 0 0 io_out[27]
port 148 nsew signal tristate
flabel metal3 s 59200 38768 60000 38888 0 FreeSans 480 0 0 0 io_out[28]
port 149 nsew signal tristate
flabel metal3 s 59200 40128 60000 40248 0 FreeSans 480 0 0 0 io_out[29]
port 150 nsew signal tristate
flabel metal3 s 59200 3408 60000 3528 0 FreeSans 480 0 0 0 io_out[2]
port 151 nsew signal tristate
flabel metal3 s 59200 41488 60000 41608 0 FreeSans 480 0 0 0 io_out[30]
port 152 nsew signal tristate
flabel metal3 s 59200 42848 60000 42968 0 FreeSans 480 0 0 0 io_out[31]
port 153 nsew signal tristate
flabel metal3 s 59200 44208 60000 44328 0 FreeSans 480 0 0 0 io_out[32]
port 154 nsew signal tristate
flabel metal3 s 59200 45568 60000 45688 0 FreeSans 480 0 0 0 io_out[33]
port 155 nsew signal tristate
flabel metal3 s 59200 46928 60000 47048 0 FreeSans 480 0 0 0 io_out[34]
port 156 nsew signal tristate
flabel metal3 s 59200 48288 60000 48408 0 FreeSans 480 0 0 0 io_out[35]
port 157 nsew signal tristate
flabel metal3 s 59200 49648 60000 49768 0 FreeSans 480 0 0 0 io_out[36]
port 158 nsew signal tristate
flabel metal3 s 59200 51008 60000 51128 0 FreeSans 480 0 0 0 io_out[37]
port 159 nsew signal tristate
flabel metal3 s 59200 4768 60000 4888 0 FreeSans 480 0 0 0 io_out[3]
port 160 nsew signal tristate
flabel metal3 s 59200 6128 60000 6248 0 FreeSans 480 0 0 0 io_out[4]
port 161 nsew signal tristate
flabel metal3 s 59200 7488 60000 7608 0 FreeSans 480 0 0 0 io_out[5]
port 162 nsew signal tristate
flabel metal3 s 59200 8848 60000 8968 0 FreeSans 480 0 0 0 io_out[6]
port 163 nsew signal tristate
flabel metal3 s 59200 10208 60000 10328 0 FreeSans 480 0 0 0 io_out[7]
port 164 nsew signal tristate
flabel metal3 s 59200 11568 60000 11688 0 FreeSans 480 0 0 0 io_out[8]
port 165 nsew signal tristate
flabel metal3 s 59200 12928 60000 13048 0 FreeSans 480 0 0 0 io_out[9]
port 166 nsew signal tristate
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 irq[0]
port 167 nsew signal tristate
flabel metal2 s 50710 0 50766 800 0 FreeSans 224 90 0 0 irq[1]
port 168 nsew signal tristate
flabel metal2 s 50802 0 50858 800 0 FreeSans 224 90 0 0 irq[2]
port 169 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 170 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 171 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 172 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 173 nsew signal input
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 174 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 175 nsew signal input
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 176 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 177 nsew signal input
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 178 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 179 nsew signal input
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 180 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 181 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 182 nsew signal input
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 183 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 184 nsew signal input
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 185 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 186 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 187 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 188 nsew signal input
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 189 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 190 nsew signal input
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 191 nsew signal input
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 192 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 193 nsew signal input
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 194 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 195 nsew signal input
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 196 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 197 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 198 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 199 nsew signal input
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 200 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 201 nsew signal input
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 202 nsew signal input
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 203 nsew signal input
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 204 nsew signal input
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 205 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 206 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 207 nsew signal input
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 208 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 209 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 210 nsew signal input
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 211 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 212 nsew signal input
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 213 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 214 nsew signal input
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 215 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 216 nsew signal input
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 217 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 218 nsew signal input
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 219 nsew signal input
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 220 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 221 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 222 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 223 nsew signal input
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 224 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 225 nsew signal input
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 226 nsew signal input
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 227 nsew signal input
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 228 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 229 nsew signal input
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 230 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 231 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 232 nsew signal input
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 233 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 234 nsew signal input
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 235 nsew signal input
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 236 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 237 nsew signal input
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 238 nsew signal input
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 239 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 240 nsew signal input
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 241 nsew signal input
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 242 nsew signal input
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 243 nsew signal input
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 244 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 245 nsew signal input
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 246 nsew signal input
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 247 nsew signal input
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 248 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 249 nsew signal input
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 250 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 251 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 252 nsew signal input
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 253 nsew signal input
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 254 nsew signal input
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 255 nsew signal input
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 256 nsew signal input
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 257 nsew signal input
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 258 nsew signal input
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 259 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 260 nsew signal input
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 261 nsew signal input
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 262 nsew signal input
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 263 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 264 nsew signal input
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 265 nsew signal input
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 266 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 267 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 268 nsew signal input
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 269 nsew signal input
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 270 nsew signal input
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 271 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 272 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 273 nsew signal input
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 274 nsew signal input
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 275 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 276 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 277 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 278 nsew signal input
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 279 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 280 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 281 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 282 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 283 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 284 nsew signal input
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 285 nsew signal input
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 286 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 287 nsew signal input
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 288 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 289 nsew signal input
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 290 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 291 nsew signal input
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 292 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 293 nsew signal input
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 294 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 295 nsew signal input
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 296 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 297 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 298 nsew signal tristate
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 299 nsew signal tristate
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 300 nsew signal tristate
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 301 nsew signal tristate
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 302 nsew signal tristate
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 303 nsew signal tristate
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 304 nsew signal tristate
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 305 nsew signal tristate
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 306 nsew signal tristate
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 307 nsew signal tristate
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 308 nsew signal tristate
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 309 nsew signal tristate
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 310 nsew signal tristate
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 311 nsew signal tristate
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 312 nsew signal tristate
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 313 nsew signal tristate
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 314 nsew signal tristate
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 315 nsew signal tristate
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 316 nsew signal tristate
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 317 nsew signal tristate
flabel metal2 s 47950 0 48006 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 318 nsew signal tristate
flabel metal2 s 48226 0 48282 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 319 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 320 nsew signal tristate
flabel metal2 s 48502 0 48558 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 321 nsew signal tristate
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 322 nsew signal tristate
flabel metal2 s 49054 0 49110 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 323 nsew signal tristate
flabel metal2 s 49330 0 49386 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 324 nsew signal tristate
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 325 nsew signal tristate
flabel metal2 s 49882 0 49938 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 326 nsew signal tristate
flabel metal2 s 50158 0 50214 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 327 nsew signal tristate
flabel metal2 s 50434 0 50490 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 328 nsew signal tristate
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 329 nsew signal tristate
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 330 nsew signal tristate
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 331 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 332 nsew signal tristate
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 333 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 334 nsew signal tristate
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 335 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 336 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 337 nsew signal tristate
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 338 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 339 nsew signal tristate
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 340 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 341 nsew signal tristate
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 342 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 343 nsew signal tristate
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 344 nsew signal tristate
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 345 nsew signal tristate
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 346 nsew signal tristate
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 347 nsew signal tristate
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 348 nsew signal tristate
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 349 nsew signal tristate
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 350 nsew signal tristate
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 351 nsew signal tristate
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 352 nsew signal tristate
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 353 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 354 nsew signal tristate
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 355 nsew signal tristate
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 356 nsew signal tristate
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 357 nsew signal tristate
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 358 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 359 nsew signal tristate
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 360 nsew signal tristate
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 361 nsew signal tristate
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 362 nsew signal tristate
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 363 nsew signal tristate
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 364 nsew signal tristate
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 365 nsew signal tristate
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 366 nsew signal tristate
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 367 nsew signal tristate
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 368 nsew signal tristate
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 369 nsew signal tristate
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 370 nsew signal tristate
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 371 nsew signal tristate
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 372 nsew signal tristate
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 373 nsew signal tristate
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 374 nsew signal tristate
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 375 nsew signal tristate
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 376 nsew signal tristate
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 377 nsew signal tristate
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 378 nsew signal tristate
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 379 nsew signal tristate
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 380 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 381 nsew signal tristate
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 382 nsew signal tristate
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 383 nsew signal tristate
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 384 nsew signal tristate
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 385 nsew signal tristate
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 386 nsew signal tristate
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 387 nsew signal tristate
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 388 nsew signal tristate
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 389 nsew signal tristate
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 390 nsew signal tristate
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 391 nsew signal tristate
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 392 nsew signal tristate
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 393 nsew signal tristate
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 394 nsew signal tristate
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 395 nsew signal tristate
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 396 nsew signal tristate
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 397 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 398 nsew signal tristate
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 399 nsew signal tristate
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 400 nsew signal tristate
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 401 nsew signal tristate
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 402 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 403 nsew signal tristate
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 404 nsew signal tristate
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 405 nsew signal tristate
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 406 nsew signal tristate
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 407 nsew signal tristate
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 408 nsew signal tristate
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 409 nsew signal tristate
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 410 nsew signal tristate
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 411 nsew signal tristate
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 412 nsew signal tristate
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 413 nsew signal tristate
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 414 nsew signal tristate
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 415 nsew signal tristate
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 416 nsew signal tristate
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 417 nsew signal tristate
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 418 nsew signal tristate
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 419 nsew signal tristate
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 420 nsew signal tristate
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 421 nsew signal tristate
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 422 nsew signal tristate
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 423 nsew signal tristate
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 424 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 425 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 426 nsew signal input
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 427 nsew signal input
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 428 nsew signal input
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 429 nsew signal input
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 430 nsew signal input
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 431 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 432 nsew signal input
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 433 nsew signal input
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 434 nsew signal input
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 435 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 436 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 437 nsew signal input
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 438 nsew signal input
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 439 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 440 nsew signal input
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 441 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 442 nsew signal input
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 443 nsew signal input
flabel metal2 s 47490 0 47546 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 444 nsew signal input
flabel metal2 s 47766 0 47822 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 445 nsew signal input
flabel metal2 s 48042 0 48098 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 446 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 447 nsew signal input
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 448 nsew signal input
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 449 nsew signal input
flabel metal2 s 48870 0 48926 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 450 nsew signal input
flabel metal2 s 49146 0 49202 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 451 nsew signal input
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 452 nsew signal input
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 453 nsew signal input
flabel metal2 s 49974 0 50030 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 454 nsew signal input
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 455 nsew signal input
flabel metal2 s 50526 0 50582 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 456 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 457 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 458 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 459 nsew signal input
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 460 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 461 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 462 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 463 nsew signal input
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 464 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 465 nsew signal input
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 466 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 467 nsew signal input
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 468 nsew signal input
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 469 nsew signal input
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 470 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 471 nsew signal input
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 472 nsew signal input
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 473 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 474 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 475 nsew signal input
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 476 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 477 nsew signal input
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 478 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 479 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 480 nsew signal input
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 481 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 482 nsew signal input
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 483 nsew signal input
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 484 nsew signal input
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 485 nsew signal input
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 486 nsew signal input
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 487 nsew signal input
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 488 nsew signal input
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 489 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 490 nsew signal input
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 491 nsew signal input
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 492 nsew signal input
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 493 nsew signal input
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 494 nsew signal input
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 495 nsew signal input
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 496 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 497 nsew signal input
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 498 nsew signal input
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 499 nsew signal input
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 500 nsew signal input
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 501 nsew signal input
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 502 nsew signal input
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 503 nsew signal input
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 504 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 505 nsew signal input
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 506 nsew signal input
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 507 nsew signal input
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 508 nsew signal input
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 509 nsew signal input
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 510 nsew signal input
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 511 nsew signal input
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 512 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 513 nsew signal input
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 514 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 515 nsew signal input
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 516 nsew signal input
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 517 nsew signal input
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 518 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 519 nsew signal input
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 520 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 521 nsew signal input
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 522 nsew signal input
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 523 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 524 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 525 nsew signal input
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 526 nsew signal input
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 527 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 528 nsew signal input
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 529 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 530 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 531 nsew signal input
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 532 nsew signal input
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 533 nsew signal input
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 534 nsew signal input
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 535 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 536 nsew signal input
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 537 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 538 nsew signal input
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 539 nsew signal input
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 540 nsew signal input
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 541 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 542 nsew signal input
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 543 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 544 nsew signal input
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 545 nsew signal input
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 546 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 547 nsew signal input
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 548 nsew signal input
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 549 nsew signal input
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 550 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 551 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 552 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 553 nsew signal input
flabel metal3 s 59200 53728 60000 53848 0 FreeSans 480 0 0 0 rst_o
port 554 nsew signal tristate
flabel metal3 s 59200 56448 60000 56568 0 FreeSans 480 0 0 0 start_o
port 555 nsew signal tristate
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 556 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 556 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 557 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 557 nsew ground bidirectional
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 wb_clk_i
port 558 nsew signal input
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 wb_rst_i
port 559 nsew signal input
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 560 nsew signal tristate
flabel metal2 s 6090 0 6146 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 561 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 562 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 563 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 564 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 565 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 566 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 567 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 568 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 569 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 570 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 571 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 572 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 573 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 574 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 575 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 576 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 577 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 578 nsew signal input
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 579 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 580 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 581 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 582 nsew signal input
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 583 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 584 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 585 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 586 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 587 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 588 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 589 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 590 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 591 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 592 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 593 nsew signal input
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 594 nsew signal input
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 595 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 596 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 597 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 598 nsew signal input
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 599 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 600 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 601 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 602 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 603 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 604 nsew signal input
flabel metal2 s 6550 0 6606 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 605 nsew signal input
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 606 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 607 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 608 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 609 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 610 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 611 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 612 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 613 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 614 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 615 nsew signal input
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 616 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 617 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 618 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 619 nsew signal input
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 620 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 621 nsew signal input
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 622 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 623 nsew signal input
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 624 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 625 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 626 nsew signal tristate
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 627 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 628 nsew signal tristate
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 629 nsew signal tristate
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 630 nsew signal tristate
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 631 nsew signal tristate
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 632 nsew signal tristate
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 633 nsew signal tristate
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 634 nsew signal tristate
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 635 nsew signal tristate
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 636 nsew signal tristate
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 637 nsew signal tristate
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 638 nsew signal tristate
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 639 nsew signal tristate
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 640 nsew signal tristate
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 641 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 642 nsew signal tristate
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 643 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 644 nsew signal tristate
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 645 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 646 nsew signal tristate
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 647 nsew signal tristate
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 648 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 649 nsew signal tristate
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 650 nsew signal tristate
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 651 nsew signal tristate
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 652 nsew signal tristate
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 653 nsew signal tristate
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 654 nsew signal tristate
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 655 nsew signal tristate
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 656 nsew signal tristate
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 657 nsew signal tristate
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 658 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 659 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 660 nsew signal input
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 661 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 662 nsew signal input
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 wbs_we_i
port 663 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
