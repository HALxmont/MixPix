magic
tech sky130A
magscale 1 2
timestamp 1669766749
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 410518 700408 410524 700460
rect 410576 700448 410582 700460
rect 429838 700448 429844 700460
rect 410576 700420 429844 700448
rect 410576 700408 410582 700420
rect 429838 700408 429844 700420
rect 429896 700408 429902 700460
rect 409138 700340 409144 700392
rect 409196 700380 409202 700392
rect 494790 700380 494796 700392
rect 409196 700352 494796 700380
rect 409196 700340 409202 700352
rect 494790 700340 494796 700352
rect 494848 700340 494854 700392
rect 155218 700272 155224 700324
rect 155276 700312 155282 700324
rect 202782 700312 202788 700324
rect 155276 700284 202788 700312
rect 155276 700272 155282 700284
rect 202782 700272 202788 700284
rect 202840 700272 202846 700324
rect 332502 700272 332508 700324
rect 332560 700312 332566 700324
rect 340138 700312 340144 700324
rect 332560 700284 340144 700312
rect 332560 700272 332566 700284
rect 340138 700272 340144 700284
rect 340196 700272 340202 700324
rect 407758 700272 407764 700324
rect 407816 700312 407822 700324
rect 559650 700312 559656 700324
rect 407816 700284 559656 700312
rect 407816 700272 407822 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 153010 699660 153016 699712
rect 153068 699700 153074 699712
rect 154114 699700 154120 699712
rect 153068 699672 154120 699700
rect 153068 699660 153074 699672
rect 154114 699660 154120 699672
rect 154172 699660 154178 699712
rect 149698 697688 149704 697740
rect 149756 697728 149762 697740
rect 153010 697728 153016 697740
rect 149756 697700 153016 697728
rect 149756 697688 149762 697700
rect 153010 697688 153016 697700
rect 153068 697688 153074 697740
rect 282178 696328 282184 696380
rect 282236 696368 282242 696380
rect 283834 696368 283840 696380
rect 282236 696340 283840 696368
rect 282236 696328 282242 696340
rect 283834 696328 283840 696340
rect 283892 696328 283898 696380
rect 348786 696192 348792 696244
rect 348844 696232 348850 696244
rect 359458 696232 359464 696244
rect 348844 696204 359464 696232
rect 348844 696192 348850 696204
rect 359458 696192 359464 696204
rect 359516 696192 359522 696244
rect 264238 695104 264244 695156
rect 264296 695144 264302 695156
rect 267642 695144 267648 695156
rect 264296 695116 267648 695144
rect 264296 695104 264302 695116
rect 267642 695104 267648 695116
rect 267700 695104 267706 695156
rect 299474 694764 299480 694816
rect 299532 694804 299538 694816
rect 309778 694804 309784 694816
rect 299532 694776 309784 694804
rect 299532 694764 299538 694776
rect 309778 694764 309784 694776
rect 309836 694764 309842 694816
rect 282178 687256 282184 687268
rect 280172 687228 282184 687256
rect 278682 687148 278688 687200
rect 278740 687188 278746 687200
rect 280172 687188 280200 687228
rect 282178 687216 282184 687228
rect 282236 687216 282242 687268
rect 278740 687160 280200 687188
rect 278740 687148 278746 687160
rect 359458 686468 359464 686520
rect 359516 686508 359522 686520
rect 371878 686508 371884 686520
rect 359516 686480 371884 686508
rect 359516 686468 359522 686480
rect 371878 686468 371884 686480
rect 371936 686468 371942 686520
rect 309778 685108 309784 685160
rect 309836 685148 309842 685160
rect 327718 685148 327724 685160
rect 309836 685120 327724 685148
rect 309836 685108 309842 685120
rect 327718 685108 327724 685120
rect 327776 685108 327782 685160
rect 276658 684496 276664 684548
rect 276716 684536 276722 684548
rect 278682 684536 278688 684548
rect 276716 684508 278688 684536
rect 276716 684496 276722 684508
rect 278682 684496 278688 684508
rect 278740 684496 278746 684548
rect 364334 683748 364340 683800
rect 364392 683788 364398 683800
rect 375374 683788 375380 683800
rect 364392 683760 375380 683788
rect 364392 683748 364398 683760
rect 375374 683748 375380 683760
rect 375432 683748 375438 683800
rect 371878 679600 371884 679652
rect 371936 679640 371942 679652
rect 381538 679640 381544 679652
rect 371936 679612 381544 679640
rect 371936 679600 371942 679612
rect 381538 679600 381544 679612
rect 381596 679600 381602 679652
rect 375374 678240 375380 678292
rect 375432 678280 375438 678292
rect 388438 678280 388444 678292
rect 375432 678252 388444 678280
rect 375432 678240 375438 678252
rect 388438 678240 388444 678252
rect 388496 678240 388502 678292
rect 140774 675452 140780 675504
rect 140832 675492 140838 675504
rect 155218 675492 155224 675504
rect 140832 675464 155224 675492
rect 140832 675452 140838 675464
rect 155218 675452 155224 675464
rect 155276 675452 155282 675504
rect 149698 673520 149704 673532
rect 146312 673492 149704 673520
rect 145558 673412 145564 673464
rect 145616 673452 145622 673464
rect 146312 673452 146340 673492
rect 149698 673480 149704 673492
rect 149756 673480 149762 673532
rect 217962 673520 217968 673532
rect 215312 673492 217968 673520
rect 145616 673424 146340 673452
rect 145616 673412 145622 673424
rect 212534 673412 212540 673464
rect 212592 673452 212598 673464
rect 215312 673452 215340 673492
rect 217962 673480 217968 673492
rect 218020 673480 218026 673532
rect 212592 673424 215340 673452
rect 212592 673412 212598 673424
rect 134518 672052 134524 672104
rect 134576 672092 134582 672104
rect 140774 672092 140780 672104
rect 134576 672064 140780 672092
rect 134576 672052 134582 672064
rect 140774 672052 140780 672064
rect 140832 672052 140838 672104
rect 388438 671100 388444 671152
rect 388496 671140 388502 671152
rect 391934 671140 391940 671152
rect 388496 671112 391940 671140
rect 388496 671100 388502 671112
rect 391934 671100 391940 671112
rect 391992 671100 391998 671152
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 15838 670732 15844 670744
rect 3568 670704 15844 670732
rect 3568 670692 3574 670704
rect 15838 670692 15844 670704
rect 15896 670692 15902 670744
rect 566458 670692 566464 670744
rect 566516 670732 566522 670744
rect 580166 670732 580172 670744
rect 566516 670704 580172 670732
rect 566516 670692 566522 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 212534 667944 212540 667956
rect 211172 667916 212540 667944
rect 211062 667836 211068 667888
rect 211120 667876 211126 667888
rect 211172 667876 211200 667916
rect 212534 667904 212540 667916
rect 212592 667904 212598 667956
rect 211120 667848 211200 667876
rect 211120 667836 211126 667848
rect 226978 665796 226984 665848
rect 227036 665836 227042 665848
rect 234614 665836 234620 665848
rect 227036 665808 234620 665836
rect 227036 665796 227042 665808
rect 234614 665796 234620 665808
rect 234672 665796 234678 665848
rect 391934 665184 391940 665236
rect 391992 665224 391998 665236
rect 395338 665224 395344 665236
rect 391992 665196 395344 665224
rect 391992 665184 391998 665196
rect 395338 665184 395344 665196
rect 395396 665184 395402 665236
rect 209038 663756 209044 663808
rect 209096 663796 209102 663808
rect 211062 663796 211068 663808
rect 209096 663768 211068 663796
rect 209096 663756 209102 663768
rect 211062 663756 211068 663768
rect 211120 663756 211126 663808
rect 258718 658180 258724 658232
rect 258776 658220 258782 658232
rect 264238 658220 264244 658232
rect 258776 658192 264244 658220
rect 258776 658180 258782 658192
rect 264238 658180 264244 658192
rect 264296 658180 264302 658232
rect 143166 658112 143172 658164
rect 143224 658152 143230 658164
rect 145558 658152 145564 658164
rect 143224 658124 145564 658152
rect 143224 658112 143230 658124
rect 145558 658112 145564 658124
rect 145616 658112 145622 658164
rect 141418 655528 141424 655580
rect 141476 655568 141482 655580
rect 143166 655568 143172 655580
rect 141476 655540 143172 655568
rect 141476 655528 141482 655540
rect 143166 655528 143172 655540
rect 143224 655528 143230 655580
rect 327718 655460 327724 655512
rect 327776 655500 327782 655512
rect 332686 655500 332692 655512
rect 327776 655472 332692 655500
rect 327776 655460 327782 655472
rect 332686 655460 332692 655472
rect 332744 655460 332750 655512
rect 131758 651856 131764 651908
rect 131816 651896 131822 651908
rect 134518 651896 134524 651908
rect 131816 651868 134524 651896
rect 131816 651856 131822 651868
rect 134518 651856 134524 651868
rect 134576 651856 134582 651908
rect 332686 649952 332692 650004
rect 332744 649992 332750 650004
rect 337378 649992 337384 650004
rect 332744 649964 337384 649992
rect 332744 649952 332750 649964
rect 337378 649952 337384 649964
rect 337436 649952 337442 650004
rect 381538 646484 381544 646536
rect 381596 646524 381602 646536
rect 395522 646524 395528 646536
rect 381596 646496 395528 646524
rect 381596 646484 381602 646496
rect 395522 646484 395528 646496
rect 395580 646484 395586 646536
rect 209038 644484 209044 644496
rect 205652 644456 209044 644484
rect 204898 644376 204904 644428
rect 204956 644416 204962 644428
rect 205652 644416 205680 644456
rect 209038 644444 209044 644456
rect 209096 644444 209102 644496
rect 204956 644388 205680 644416
rect 204956 644376 204962 644388
rect 337378 642132 337384 642184
rect 337436 642172 337442 642184
rect 343634 642172 343640 642184
rect 337436 642144 343640 642172
rect 337436 642132 337442 642144
rect 343634 642132 343640 642144
rect 343692 642132 343698 642184
rect 139394 641724 139400 641776
rect 139452 641764 139458 641776
rect 141418 641764 141424 641776
rect 139452 641736 141424 641764
rect 139452 641724 139458 641736
rect 141418 641724 141424 641736
rect 141476 641724 141482 641776
rect 340138 640976 340144 641028
rect 340196 641016 340202 641028
rect 352558 641016 352564 641028
rect 340196 640988 352564 641016
rect 340196 640976 340202 640988
rect 352558 640976 352564 640988
rect 352616 640976 352622 641028
rect 224218 640296 224224 640348
rect 224276 640336 224282 640348
rect 226978 640336 226984 640348
rect 224276 640308 226984 640336
rect 224276 640296 224282 640308
rect 226978 640296 226984 640308
rect 227036 640296 227042 640348
rect 343634 639548 343640 639600
rect 343692 639588 343698 639600
rect 349154 639588 349160 639600
rect 343692 639560 349160 639588
rect 343692 639548 343698 639560
rect 349154 639548 349160 639560
rect 349212 639548 349218 639600
rect 139394 638976 139400 638988
rect 136652 638948 139400 638976
rect 136542 638868 136548 638920
rect 136600 638908 136606 638920
rect 136652 638908 136680 638948
rect 139394 638936 139400 638948
rect 139452 638936 139458 638988
rect 136600 638880 136680 638908
rect 136600 638868 136606 638880
rect 349154 637508 349160 637560
rect 349212 637548 349218 637560
rect 352650 637548 352656 637560
rect 349212 637520 352656 637548
rect 349212 637508 349218 637520
rect 352650 637508 352656 637520
rect 352708 637508 352714 637560
rect 134518 635536 134524 635588
rect 134576 635576 134582 635588
rect 136542 635576 136548 635588
rect 134576 635548 136548 635576
rect 134576 635536 134582 635548
rect 136542 635536 136548 635548
rect 136600 635536 136606 635588
rect 211798 634040 211804 634092
rect 211856 634080 211862 634092
rect 224218 634080 224224 634092
rect 211856 634052 224224 634080
rect 211856 634040 211862 634052
rect 224218 634040 224224 634052
rect 224276 634040 224282 634092
rect 247034 634040 247040 634092
rect 247092 634080 247098 634092
rect 258718 634080 258724 634092
rect 247092 634052 258724 634080
rect 247092 634040 247098 634052
rect 258718 634040 258724 634052
rect 258776 634040 258782 634092
rect 203518 630640 203524 630692
rect 203576 630680 203582 630692
rect 204898 630680 204904 630692
rect 203576 630652 204904 630680
rect 203576 630640 203582 630652
rect 204898 630640 204904 630652
rect 204956 630640 204962 630692
rect 275370 630640 275376 630692
rect 275428 630680 275434 630692
rect 276658 630680 276664 630692
rect 275428 630652 276664 630680
rect 275428 630640 275434 630652
rect 276658 630640 276664 630652
rect 276716 630640 276722 630692
rect 243538 629620 243544 629672
rect 243596 629660 243602 629672
rect 247034 629660 247040 629672
rect 243596 629632 247040 629660
rect 243596 629620 243602 629632
rect 247034 629620 247040 629632
rect 247092 629620 247098 629672
rect 273898 628736 273904 628788
rect 273956 628776 273962 628788
rect 275370 628776 275376 628788
rect 273956 628748 275376 628776
rect 273956 628736 273962 628748
rect 275370 628736 275376 628748
rect 275428 628736 275434 628788
rect 352650 624384 352656 624436
rect 352708 624424 352714 624436
rect 370498 624424 370504 624436
rect 352708 624396 370504 624424
rect 352708 624384 352714 624396
rect 370498 624384 370504 624396
rect 370556 624384 370562 624436
rect 209038 623772 209044 623824
rect 209096 623812 209102 623824
rect 211798 623812 211804 623824
rect 209096 623784 211804 623812
rect 209096 623772 209102 623784
rect 211798 623772 211804 623784
rect 211856 623772 211862 623824
rect 352558 623024 352564 623076
rect 352616 623064 352622 623076
rect 360194 623064 360200 623076
rect 352616 623036 360200 623064
rect 352616 623024 352622 623036
rect 360194 623024 360200 623036
rect 360252 623024 360258 623076
rect 271138 622412 271144 622464
rect 271196 622452 271202 622464
rect 273898 622452 273904 622464
rect 271196 622424 273904 622452
rect 271196 622412 271202 622424
rect 273898 622412 273904 622424
rect 273956 622412 273962 622464
rect 123478 620984 123484 621036
rect 123536 621024 123542 621036
rect 131758 621024 131764 621036
rect 123536 620996 131764 621024
rect 123536 620984 123542 620996
rect 131758 620984 131764 620996
rect 131816 620984 131822 621036
rect 360194 619556 360200 619608
rect 360252 619596 360258 619608
rect 362954 619596 362960 619608
rect 360252 619568 362960 619596
rect 360252 619556 360258 619568
rect 362954 619556 362960 619568
rect 363012 619556 363018 619608
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 37918 618304 37924 618316
rect 3568 618276 37924 618304
rect 3568 618264 3574 618276
rect 37918 618264 37924 618276
rect 37976 618264 37982 618316
rect 406378 616836 406384 616888
rect 406436 616876 406442 616888
rect 579982 616876 579988 616888
rect 406436 616848 579988 616876
rect 406436 616836 406442 616848
rect 579982 616836 579988 616848
rect 580040 616836 580046 616888
rect 362954 616088 362960 616140
rect 363012 616128 363018 616140
rect 373258 616128 373264 616140
rect 363012 616100 373264 616128
rect 363012 616088 363018 616100
rect 373258 616088 373264 616100
rect 373316 616088 373322 616140
rect 233142 613368 233148 613420
rect 233200 613408 233206 613420
rect 243538 613408 243544 613420
rect 233200 613380 243544 613408
rect 233200 613368 233206 613380
rect 243538 613368 243544 613380
rect 243596 613368 243602 613420
rect 268378 612756 268384 612808
rect 268436 612796 268442 612808
rect 271138 612796 271144 612808
rect 268436 612768 271144 612796
rect 268436 612756 268442 612768
rect 271138 612756 271144 612768
rect 271196 612756 271202 612808
rect 200758 610512 200764 610564
rect 200816 610552 200822 610564
rect 203518 610552 203524 610564
rect 200816 610524 203524 610552
rect 200816 610512 200822 610524
rect 203518 610512 203524 610524
rect 203576 610512 203582 610564
rect 59262 609220 59268 609272
rect 59320 609260 59326 609272
rect 123478 609260 123484 609272
rect 59320 609232 123484 609260
rect 59320 609220 59326 609232
rect 123478 609220 123484 609232
rect 123536 609220 123542 609272
rect 224218 609220 224224 609272
rect 224276 609260 224282 609272
rect 233142 609260 233148 609272
rect 224276 609232 233148 609260
rect 224276 609220 224282 609232
rect 233142 609220 233148 609232
rect 233200 609220 233206 609272
rect 53098 606432 53104 606484
rect 53156 606472 53162 606484
rect 59262 606472 59268 606484
rect 53156 606444 59268 606472
rect 53156 606432 53162 606444
rect 59262 606432 59268 606444
rect 59320 606432 59326 606484
rect 266998 604460 267004 604512
rect 267056 604500 267062 604512
rect 268378 604500 268384 604512
rect 267056 604472 268384 604500
rect 267056 604460 267062 604472
rect 268378 604460 268384 604472
rect 268436 604460 268442 604512
rect 370498 602352 370504 602404
rect 370556 602392 370562 602404
rect 387058 602392 387064 602404
rect 370556 602364 387064 602392
rect 370556 602352 370562 602364
rect 387058 602352 387064 602364
rect 387116 602352 387122 602404
rect 373258 599564 373264 599616
rect 373316 599604 373322 599616
rect 397546 599604 397552 599616
rect 373316 599576 397552 599604
rect 373316 599564 373322 599576
rect 397546 599564 397552 599576
rect 397604 599564 397610 599616
rect 131758 597524 131764 597576
rect 131816 597564 131822 597576
rect 134518 597564 134524 597576
rect 131816 597536 134524 597564
rect 131816 597524 131822 597536
rect 134518 597524 134524 597536
rect 134576 597524 134582 597576
rect 195238 593308 195244 593360
rect 195296 593348 195302 593360
rect 200758 593348 200764 593360
rect 195296 593320 200764 593348
rect 195296 593308 195302 593320
rect 200758 593308 200764 593320
rect 200816 593308 200822 593360
rect 214558 591268 214564 591320
rect 214616 591308 214622 591320
rect 224218 591308 224224 591320
rect 214616 591280 224224 591308
rect 214616 591268 214622 591280
rect 224218 591268 224224 591280
rect 224276 591268 224282 591320
rect 211798 585148 211804 585200
rect 211856 585188 211862 585200
rect 214558 585188 214564 585200
rect 211856 585160 214564 585188
rect 211856 585148 211862 585160
rect 214558 585148 214564 585160
rect 214616 585148 214622 585200
rect 200758 583720 200764 583772
rect 200816 583760 200822 583772
rect 209038 583760 209044 583772
rect 200816 583732 209044 583760
rect 200816 583720 200822 583732
rect 209038 583720 209044 583732
rect 209096 583720 209102 583772
rect 387058 573996 387064 574048
rect 387116 574036 387122 574048
rect 393958 574036 393964 574048
rect 387116 574008 393964 574036
rect 387116 573996 387122 574008
rect 393958 573996 393964 574008
rect 394016 573996 394022 574048
rect 265710 572704 265716 572756
rect 265768 572744 265774 572756
rect 266998 572744 267004 572756
rect 265768 572716 267004 572744
rect 265768 572704 265774 572716
rect 266998 572704 267004 572716
rect 267056 572704 267062 572756
rect 264238 570664 264244 570716
rect 264296 570704 264302 570716
rect 265710 570704 265716 570716
rect 264296 570676 265716 570704
rect 264296 570664 264302 570676
rect 265710 570664 265716 570676
rect 265768 570664 265774 570716
rect 3326 565836 3332 565888
rect 3384 565876 3390 565888
rect 29638 565876 29644 565888
rect 3384 565848 29644 565876
rect 3384 565836 3390 565848
rect 29638 565836 29644 565848
rect 29696 565836 29702 565888
rect 197998 564952 198004 565004
rect 198056 564992 198062 565004
rect 200758 564992 200764 565004
rect 198056 564964 200764 564992
rect 198056 564952 198062 564964
rect 200758 564952 200764 564964
rect 200816 564952 200822 565004
rect 404998 563048 405004 563100
rect 405056 563088 405062 563100
rect 580166 563088 580172 563100
rect 405056 563060 580172 563088
rect 405056 563048 405062 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 393958 562640 393964 562692
rect 394016 562680 394022 562692
rect 395430 562680 395436 562692
rect 394016 562652 395436 562680
rect 394016 562640 394022 562652
rect 395430 562640 395436 562652
rect 395488 562640 395494 562692
rect 193950 560260 193956 560312
rect 194008 560300 194014 560312
rect 195238 560300 195244 560312
rect 194008 560272 195244 560300
rect 194008 560260 194014 560272
rect 195238 560260 195244 560272
rect 195296 560260 195302 560312
rect 46198 559716 46204 559768
rect 46256 559756 46262 559768
rect 53098 559756 53104 559768
rect 46256 559728 53104 559756
rect 46256 559716 46262 559728
rect 53098 559716 53104 559728
rect 53156 559716 53162 559768
rect 192478 558560 192484 558612
rect 192536 558600 192542 558612
rect 193950 558600 193956 558612
rect 192536 558572 193956 558600
rect 192536 558560 192542 558572
rect 193950 558560 193956 558572
rect 194008 558560 194014 558612
rect 2774 553800 2780 553852
rect 2832 553840 2838 553852
rect 4798 553840 4804 553852
rect 2832 553812 4804 553840
rect 2832 553800 2838 553812
rect 4798 553800 4804 553812
rect 4856 553800 4862 553852
rect 261478 553392 261484 553444
rect 261536 553432 261542 553444
rect 264238 553432 264244 553444
rect 261536 553404 264244 553432
rect 261536 553392 261542 553404
rect 264238 553392 264244 553404
rect 264296 553392 264302 553444
rect 206278 549244 206284 549296
rect 206336 549284 206342 549296
rect 211798 549284 211804 549296
rect 206336 549256 211804 549284
rect 206336 549244 206342 549256
rect 211798 549244 211804 549256
rect 211856 549244 211862 549296
rect 191098 546456 191104 546508
rect 191156 546496 191162 546508
rect 192478 546496 192484 546508
rect 191156 546468 192484 546496
rect 191156 546456 191162 546468
rect 192478 546456 192484 546468
rect 192536 546456 192542 546508
rect 189718 538840 189724 538892
rect 189776 538880 189782 538892
rect 197998 538880 198004 538892
rect 189776 538852 198004 538880
rect 189776 538840 189782 538852
rect 197998 538840 198004 538852
rect 198056 538840 198062 538892
rect 62666 537480 62672 537532
rect 62724 537520 62730 537532
rect 169754 537520 169760 537532
rect 62724 537492 169760 537520
rect 62724 537480 62730 537492
rect 169754 537480 169760 537492
rect 169812 537480 169818 537532
rect 188338 535100 188344 535152
rect 188396 535140 188402 535152
rect 191098 535140 191104 535152
rect 188396 535112 191104 535140
rect 188396 535100 188402 535112
rect 191098 535100 191104 535112
rect 191156 535100 191162 535152
rect 130378 533332 130384 533384
rect 130436 533372 130442 533384
rect 131758 533372 131764 533384
rect 130436 533344 131764 533372
rect 130436 533332 130442 533344
rect 131758 533332 131764 533344
rect 131816 533332 131822 533384
rect 61378 532992 61384 533044
rect 61436 533032 61442 533044
rect 62666 533032 62672 533044
rect 61436 533004 62672 533032
rect 61436 532992 61442 533004
rect 62666 532992 62672 533004
rect 62724 532992 62730 533044
rect 260098 531224 260104 531276
rect 260156 531264 260162 531276
rect 261478 531264 261484 531276
rect 260156 531236 261484 531264
rect 260156 531224 260162 531236
rect 261478 531224 261484 531236
rect 261536 531224 261542 531276
rect 128998 527144 129004 527196
rect 129056 527184 129062 527196
rect 130378 527184 130384 527196
rect 129056 527156 130384 527184
rect 129056 527144 129062 527156
rect 130378 527144 130384 527156
rect 130436 527144 130442 527196
rect 200758 524424 200764 524476
rect 200816 524464 200822 524476
rect 206278 524464 206284 524476
rect 200816 524436 206284 524464
rect 200816 524424 200822 524436
rect 206278 524424 206284 524436
rect 206336 524424 206342 524476
rect 257338 518916 257344 518968
rect 257396 518956 257402 518968
rect 260098 518956 260104 518968
rect 257396 518928 260104 518956
rect 257396 518916 257402 518928
rect 260098 518916 260104 518928
rect 260156 518916 260162 518968
rect 45094 517488 45100 517540
rect 45152 517528 45158 517540
rect 46198 517528 46204 517540
rect 45152 517500 46204 517528
rect 45152 517488 45158 517500
rect 46198 517488 46204 517500
rect 46256 517488 46262 517540
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 33778 514808 33784 514820
rect 3384 514780 33784 514808
rect 3384 514768 3390 514780
rect 33778 514768 33784 514780
rect 33836 514768 33842 514820
rect 153194 511232 153200 511284
rect 153252 511272 153258 511284
rect 189718 511272 189724 511284
rect 153252 511244 189724 511272
rect 153252 511232 153258 511244
rect 189718 511232 189724 511244
rect 189776 511232 189782 511284
rect 403618 510620 403624 510672
rect 403676 510660 403682 510672
rect 579798 510660 579804 510672
rect 403676 510632 579804 510660
rect 403676 510620 403682 510632
rect 579798 510620 579804 510632
rect 579856 510620 579862 510672
rect 117958 508512 117964 508564
rect 118016 508552 118022 508564
rect 136634 508552 136640 508564
rect 118016 508524 136640 508552
rect 118016 508512 118022 508524
rect 136634 508512 136640 508524
rect 136692 508512 136698 508564
rect 150434 507832 150440 507884
rect 150492 507872 150498 507884
rect 153194 507872 153200 507884
rect 150492 507844 153200 507872
rect 150492 507832 150498 507844
rect 153194 507832 153200 507844
rect 153252 507832 153258 507884
rect 192478 505724 192484 505776
rect 192536 505764 192542 505776
rect 200758 505764 200764 505776
rect 192536 505736 200764 505764
rect 192536 505724 192542 505736
rect 200758 505724 200764 505736
rect 200816 505724 200822 505776
rect 257338 502364 257344 502376
rect 255332 502336 257344 502364
rect 253934 502256 253940 502308
rect 253992 502296 253998 502308
rect 255332 502296 255360 502336
rect 257338 502324 257344 502336
rect 257396 502324 257402 502376
rect 253992 502268 255360 502296
rect 253992 502256 253998 502268
rect 143534 501712 143540 501764
rect 143592 501752 143598 501764
rect 150434 501752 150440 501764
rect 143592 501724 150440 501752
rect 143592 501712 143598 501724
rect 150434 501712 150440 501724
rect 150492 501712 150498 501764
rect 2774 501032 2780 501084
rect 2832 501072 2838 501084
rect 4890 501072 4896 501084
rect 2832 501044 4896 501072
rect 2832 501032 2838 501044
rect 4890 501032 4896 501044
rect 4948 501032 4954 501084
rect 126974 500896 126980 500948
rect 127032 500936 127038 500948
rect 128998 500936 129004 500948
rect 127032 500908 129004 500936
rect 127032 500896 127038 500908
rect 128998 500896 129004 500908
rect 129056 500896 129062 500948
rect 180058 498788 180064 498840
rect 180116 498828 180122 498840
rect 192478 498828 192484 498840
rect 180116 498800 192484 498828
rect 180116 498788 180122 498800
rect 192478 498788 192484 498800
rect 192536 498788 192542 498840
rect 253934 498216 253940 498228
rect 252572 498188 253940 498216
rect 249518 498108 249524 498160
rect 249576 498148 249582 498160
rect 252572 498148 252600 498188
rect 253934 498176 253940 498188
rect 253992 498176 253998 498228
rect 249576 498120 252600 498148
rect 249576 498108 249582 498120
rect 126974 496856 126980 496868
rect 125612 496828 126980 496856
rect 124858 496748 124864 496800
rect 124916 496788 124922 496800
rect 125612 496788 125640 496828
rect 126974 496816 126980 496828
rect 127032 496816 127038 496868
rect 124916 496760 125640 496788
rect 124916 496748 124922 496760
rect 140038 496680 140044 496732
rect 140096 496720 140102 496732
rect 143534 496720 143540 496732
rect 140096 496692 143540 496720
rect 140096 496680 140102 496692
rect 143534 496680 143540 496692
rect 143592 496680 143598 496732
rect 246298 495456 246304 495508
rect 246356 495496 246362 495508
rect 249518 495496 249524 495508
rect 246356 495468 249524 495496
rect 246356 495456 246362 495468
rect 249518 495456 249524 495468
rect 249576 495456 249582 495508
rect 116578 487160 116584 487212
rect 116636 487200 116642 487212
rect 117958 487200 117964 487212
rect 116636 487172 117964 487200
rect 116636 487160 116642 487172
rect 117958 487160 117964 487172
rect 118016 487160 118022 487212
rect 136450 487160 136456 487212
rect 136508 487200 136514 487212
rect 140038 487200 140044 487212
rect 136508 487172 140044 487200
rect 136508 487160 136514 487172
rect 140038 487160 140044 487172
rect 140096 487160 140102 487212
rect 175918 481992 175924 482044
rect 175976 482032 175982 482044
rect 180058 482032 180064 482044
rect 175976 482004 180064 482032
rect 175976 481992 175982 482004
rect 180058 481992 180064 482004
rect 180116 481992 180122 482044
rect 133138 481448 133144 481500
rect 133196 481488 133202 481500
rect 136450 481488 136456 481500
rect 133196 481460 136456 481488
rect 133196 481448 133202 481460
rect 136450 481448 136456 481460
rect 136508 481448 136514 481500
rect 123478 473968 123484 474020
rect 123536 474008 123542 474020
rect 124858 474008 124864 474020
rect 123536 473980 124864 474008
rect 123536 473968 123542 473980
rect 124858 473968 124864 473980
rect 124916 473968 124922 474020
rect 115198 472948 115204 473000
rect 115256 472988 115262 473000
rect 116578 472988 116584 473000
rect 115256 472960 116584 472988
rect 115256 472948 115262 472960
rect 116578 472948 116584 472960
rect 116636 472948 116642 473000
rect 246298 472036 246304 472048
rect 240152 472008 246304 472036
rect 239398 471928 239404 471980
rect 239456 471968 239462 471980
rect 240152 471968 240180 472008
rect 246298 471996 246304 472008
rect 246356 471996 246362 472048
rect 239456 471940 240180 471968
rect 239456 471928 239462 471940
rect 122098 464992 122104 465044
rect 122156 465032 122162 465044
rect 123478 465032 123484 465044
rect 122156 465004 123484 465032
rect 122156 464992 122162 465004
rect 123478 464992 123484 465004
rect 123536 464992 123542 465044
rect 2774 462544 2780 462596
rect 2832 462584 2838 462596
rect 5074 462584 5080 462596
rect 2832 462556 5080 462584
rect 2832 462544 2838 462556
rect 5074 462544 5080 462556
rect 5132 462544 5138 462596
rect 163498 460164 163504 460216
rect 163556 460204 163562 460216
rect 175918 460204 175924 460216
rect 163556 460176 175924 460204
rect 163556 460164 163562 460176
rect 175918 460164 175924 460176
rect 175976 460164 175982 460216
rect 400858 456764 400864 456816
rect 400916 456804 400922 456816
rect 579982 456804 579988 456816
rect 400916 456776 579988 456804
rect 400916 456764 400922 456776
rect 579982 456764 579988 456776
rect 580040 456764 580046 456816
rect 188338 455444 188344 455456
rect 186332 455416 188344 455444
rect 182818 455336 182824 455388
rect 182876 455376 182882 455388
rect 186332 455376 186360 455416
rect 188338 455404 188344 455416
rect 188396 455404 188402 455456
rect 182876 455348 186360 455376
rect 182876 455336 182882 455348
rect 238018 451256 238024 451308
rect 238076 451296 238082 451308
rect 239398 451296 239404 451308
rect 238076 451268 239404 451296
rect 238076 451256 238082 451268
rect 239398 451256 239404 451268
rect 239456 451256 239462 451308
rect 127618 449896 127624 449948
rect 127676 449936 127682 449948
rect 133138 449936 133144 449948
rect 127676 449908 133144 449936
rect 127676 449896 127682 449908
rect 133138 449896 133144 449908
rect 133196 449896 133202 449948
rect 2774 448808 2780 448860
rect 2832 448848 2838 448860
rect 4982 448848 4988 448860
rect 2832 448820 4988 448848
rect 2832 448808 2838 448820
rect 4982 448808 4988 448820
rect 5040 448808 5046 448860
rect 160738 446972 160744 447024
rect 160796 447012 160802 447024
rect 163498 447012 163504 447024
rect 160796 446984 163504 447012
rect 160796 446972 160802 446984
rect 163498 446972 163504 446984
rect 163556 446972 163562 447024
rect 119430 446156 119436 446208
rect 119488 446196 119494 446208
rect 122098 446196 122104 446208
rect 119488 446168 122104 446196
rect 119488 446156 119494 446168
rect 122098 446156 122104 446168
rect 122156 446156 122162 446208
rect 399478 444388 399484 444440
rect 399536 444428 399542 444440
rect 579982 444428 579988 444440
rect 399536 444400 579988 444428
rect 399536 444388 399542 444400
rect 579982 444388 579988 444400
rect 580040 444388 580046 444440
rect 181438 438880 181444 438932
rect 181496 438920 181502 438932
rect 182818 438920 182824 438932
rect 181496 438892 182824 438920
rect 181496 438880 181502 438892
rect 182818 438880 182824 438892
rect 182876 438880 182882 438932
rect 117958 433236 117964 433288
rect 118016 433276 118022 433288
rect 119430 433276 119436 433288
rect 118016 433248 119436 433276
rect 118016 433236 118022 433248
rect 119430 433236 119436 433248
rect 119488 433236 119494 433288
rect 119338 432556 119344 432608
rect 119396 432596 119402 432608
rect 127618 432596 127624 432608
rect 119396 432568 127624 432596
rect 119396 432556 119402 432568
rect 127618 432556 127624 432568
rect 127676 432556 127682 432608
rect 236638 427796 236644 427848
rect 236696 427836 236702 427848
rect 238018 427836 238024 427848
rect 236696 427808 238024 427836
rect 236696 427796 236702 427808
rect 238018 427796 238024 427808
rect 238076 427796 238082 427848
rect 116578 416712 116584 416764
rect 116636 416752 116642 416764
rect 117958 416752 117964 416764
rect 116636 416724 117964 416752
rect 116636 416712 116642 416724
rect 117958 416712 117964 416724
rect 118016 416712 118022 416764
rect 179322 413992 179328 414044
rect 179380 414032 179386 414044
rect 181438 414032 181444 414044
rect 179380 414004 181444 414032
rect 179380 413992 179386 414004
rect 181438 413992 181444 414004
rect 181496 413992 181502 414044
rect 3142 410048 3148 410100
rect 3200 410088 3206 410100
rect 8938 410088 8944 410100
rect 3200 410060 8944 410088
rect 3200 410048 3206 410060
rect 8938 410048 8944 410060
rect 8996 410048 9002 410100
rect 177298 409844 177304 409896
rect 177356 409884 177362 409896
rect 179322 409884 179328 409896
rect 177356 409856 179328 409884
rect 177356 409844 177362 409856
rect 179322 409844 179328 409856
rect 179380 409844 179386 409896
rect 115290 407192 115296 407244
rect 115348 407232 115354 407244
rect 116578 407232 116584 407244
rect 115348 407204 116584 407232
rect 115348 407192 115354 407204
rect 116578 407192 116584 407204
rect 116636 407192 116642 407244
rect 113910 405424 113916 405476
rect 113968 405464 113974 405476
rect 115290 405464 115296 405476
rect 113968 405436 115296 405464
rect 113968 405424 113974 405436
rect 115290 405424 115296 405436
rect 115348 405424 115354 405476
rect 417418 404336 417424 404388
rect 417476 404376 417482 404388
rect 579982 404376 579988 404388
rect 417476 404348 579988 404376
rect 417476 404336 417482 404348
rect 579982 404336 579988 404348
rect 580040 404336 580046 404388
rect 233878 404268 233884 404320
rect 233936 404308 233942 404320
rect 236638 404308 236644 404320
rect 233936 404280 236644 404308
rect 233936 404268 233942 404280
rect 236638 404268 236644 404280
rect 236696 404268 236702 404320
rect 112438 398488 112444 398540
rect 112496 398528 112502 398540
rect 113910 398528 113916 398540
rect 112496 398500 113916 398528
rect 112496 398488 112502 398500
rect 113910 398488 113916 398500
rect 113968 398488 113974 398540
rect 2774 397468 2780 397520
rect 2832 397508 2838 397520
rect 5166 397508 5172 397520
rect 2832 397480 5172 397508
rect 2832 397468 2838 397480
rect 5166 397468 5172 397480
rect 5224 397468 5230 397520
rect 110414 391960 110420 392012
rect 110472 392000 110478 392012
rect 112438 392000 112444 392012
rect 110472 391972 112444 392000
rect 110472 391960 110478 391972
rect 112438 391960 112444 391972
rect 112496 391960 112502 392012
rect 112438 385636 112444 385688
rect 112496 385676 112502 385688
rect 119338 385676 119344 385688
rect 112496 385648 119344 385676
rect 112496 385636 112502 385648
rect 119338 385636 119344 385648
rect 119396 385636 119402 385688
rect 106918 384616 106924 384668
rect 106976 384656 106982 384668
rect 110414 384656 110420 384668
rect 106976 384628 110420 384656
rect 106976 384616 106982 384628
rect 110414 384616 110420 384628
rect 110472 384616 110478 384668
rect 157978 379516 157984 379568
rect 158036 379556 158042 379568
rect 160738 379556 160744 379568
rect 158036 379528 160744 379556
rect 158036 379516 158042 379528
rect 160738 379516 160744 379528
rect 160796 379516 160802 379568
rect 396718 378156 396724 378208
rect 396776 378196 396782 378208
rect 579982 378196 579988 378208
rect 396776 378168 579988 378196
rect 396776 378156 396782 378168
rect 579982 378156 579988 378168
rect 580040 378156 580046 378208
rect 58618 376592 58624 376644
rect 58676 376632 58682 376644
rect 61378 376632 61384 376644
rect 58676 376604 61384 376632
rect 58676 376592 58682 376604
rect 61378 376592 61384 376604
rect 61436 376592 61442 376644
rect 175274 375300 175280 375352
rect 175332 375340 175338 375352
rect 177298 375340 177304 375352
rect 175332 375312 177304 375340
rect 175332 375300 175338 375312
rect 177298 375300 177304 375312
rect 177356 375300 177362 375352
rect 175274 371260 175280 371272
rect 173912 371232 175280 371260
rect 173158 371152 173164 371204
rect 173216 371192 173222 371204
rect 173912 371192 173940 371232
rect 175274 371220 175280 371232
rect 175332 371220 175338 371272
rect 173216 371164 173940 371192
rect 173216 371152 173222 371164
rect 103514 365644 103520 365696
rect 103572 365684 103578 365696
rect 112438 365684 112444 365696
rect 103572 365656 112444 365684
rect 103572 365644 103578 365656
rect 112438 365644 112444 365656
rect 112496 365644 112502 365696
rect 396902 364352 396908 364404
rect 396960 364392 396966 364404
rect 579982 364392 579988 364404
rect 396960 364364 579988 364392
rect 396960 364352 396966 364364
rect 579982 364352 579988 364364
rect 580040 364352 580046 364404
rect 78582 362176 78588 362228
rect 78640 362216 78646 362228
rect 103514 362216 103520 362228
rect 78640 362188 103520 362216
rect 78640 362176 78646 362188
rect 103514 362176 103520 362188
rect 103572 362176 103578 362228
rect 75178 357756 75184 357808
rect 75236 357796 75242 357808
rect 78582 357796 78588 357808
rect 75236 357768 78588 357796
rect 75236 357756 75242 357768
rect 78582 357756 78588 357768
rect 78640 357756 78646 357808
rect 105262 357552 105268 357604
rect 105320 357592 105326 357604
rect 106918 357592 106924 357604
rect 105320 357564 106924 357592
rect 105320 357552 105326 357564
rect 106918 357552 106924 357564
rect 106976 357552 106982 357604
rect 3326 357416 3332 357468
rect 3384 357456 3390 357468
rect 10318 357456 10324 357468
rect 3384 357428 10324 357456
rect 3384 357416 3390 357428
rect 10318 357416 10324 357428
rect 10376 357416 10382 357468
rect 69658 356668 69664 356720
rect 69716 356708 69722 356720
rect 115198 356708 115204 356720
rect 69716 356680 115204 356708
rect 69716 356668 69722 356680
rect 115198 356668 115204 356680
rect 115256 356668 115262 356720
rect 103514 355784 103520 355836
rect 103572 355824 103578 355836
rect 105262 355824 105268 355836
rect 103572 355796 105268 355824
rect 103572 355784 103578 355796
rect 105262 355784 105268 355796
rect 105320 355784 105326 355836
rect 414658 351908 414664 351960
rect 414716 351948 414722 351960
rect 579982 351948 579988 351960
rect 414716 351920 579988 351948
rect 414716 351908 414722 351920
rect 579982 351908 579988 351920
rect 580040 351908 580046 351960
rect 98638 351840 98644 351892
rect 98696 351880 98702 351892
rect 103514 351880 103520 351892
rect 98696 351852 103520 351880
rect 98696 351840 98702 351852
rect 103514 351840 103520 351852
rect 103572 351840 103578 351892
rect 231118 349460 231124 349512
rect 231176 349500 231182 349512
rect 233878 349500 233884 349512
rect 231176 349472 233884 349500
rect 231176 349460 231182 349472
rect 233878 349460 233884 349472
rect 233936 349460 233942 349512
rect 172146 349120 172152 349172
rect 172204 349160 172210 349172
rect 173158 349160 173164 349172
rect 172204 349132 173164 349160
rect 172204 349120 172210 349132
rect 173158 349120 173164 349132
rect 173216 349120 173222 349172
rect 56870 346332 56876 346384
rect 56928 346372 56934 346384
rect 58618 346372 58624 346384
rect 56928 346344 58624 346372
rect 56928 346332 56934 346344
rect 58618 346332 58624 346344
rect 58676 346332 58682 346384
rect 2774 345176 2780 345228
rect 2832 345216 2838 345228
rect 5258 345216 5264 345228
rect 2832 345188 5264 345216
rect 2832 345176 2838 345188
rect 5258 345176 5264 345188
rect 5316 345176 5322 345228
rect 170398 345040 170404 345092
rect 170456 345080 170462 345092
rect 172146 345080 172152 345092
rect 170456 345052 172152 345080
rect 170456 345040 170462 345052
rect 172146 345040 172152 345052
rect 172204 345040 172210 345092
rect 94498 340892 94504 340944
rect 94556 340932 94562 340944
rect 98638 340932 98644 340944
rect 94556 340904 98644 340932
rect 94556 340892 94562 340904
rect 98638 340892 98644 340904
rect 98696 340892 98702 340944
rect 68278 339668 68284 339720
rect 68336 339708 68342 339720
rect 69658 339708 69664 339720
rect 68336 339680 69664 339708
rect 68336 339668 68342 339680
rect 69658 339668 69664 339680
rect 69716 339668 69722 339720
rect 55858 338240 55864 338292
rect 55916 338280 55922 338292
rect 56870 338280 56876 338292
rect 55916 338252 56876 338280
rect 55916 338240 55922 338252
rect 56870 338240 56876 338252
rect 56928 338240 56934 338292
rect 566550 338104 566556 338156
rect 566608 338144 566614 338156
rect 579982 338144 579988 338156
rect 566608 338116 579988 338144
rect 566608 338104 566614 338116
rect 579982 338104 579988 338116
rect 580040 338104 580046 338156
rect 66254 335996 66260 336048
rect 66312 336036 66318 336048
rect 75178 336036 75184 336048
rect 66312 336008 75184 336036
rect 66312 335996 66318 336008
rect 75178 335996 75184 336008
rect 75236 335996 75242 336048
rect 48958 331848 48964 331900
rect 49016 331888 49022 331900
rect 66254 331888 66260 331900
rect 49016 331860 66260 331888
rect 49016 331848 49022 331860
rect 66254 331848 66260 331860
rect 66312 331848 66318 331900
rect 167638 330352 167644 330404
rect 167696 330392 167702 330404
rect 170398 330392 170404 330404
rect 167696 330364 170404 330392
rect 167696 330352 167702 330364
rect 170398 330352 170404 330364
rect 170456 330352 170462 330404
rect 396810 324300 396816 324352
rect 396868 324340 396874 324352
rect 579798 324340 579804 324352
rect 396868 324312 579804 324340
rect 396868 324300 396874 324312
rect 579798 324300 579804 324312
rect 579856 324300 579862 324352
rect 53098 323348 53104 323400
rect 53156 323388 53162 323400
rect 55858 323388 55864 323400
rect 53156 323360 55864 323388
rect 53156 323348 53162 323360
rect 55858 323348 55864 323360
rect 55916 323348 55922 323400
rect 165614 322940 165620 322992
rect 165672 322980 165678 322992
rect 167638 322980 167644 322992
rect 165672 322952 167644 322980
rect 165672 322940 165678 322952
rect 167638 322940 167644 322952
rect 167696 322940 167702 322992
rect 231118 321620 231124 321632
rect 229066 321592 231124 321620
rect 228358 321512 228364 321564
rect 228416 321552 228422 321564
rect 229066 321552 229094 321592
rect 231118 321580 231124 321592
rect 231176 321580 231182 321632
rect 228416 321524 229094 321552
rect 228416 321512 228422 321524
rect 162118 320424 162124 320476
rect 162176 320464 162182 320476
rect 165614 320464 165620 320476
rect 162176 320436 165620 320464
rect 162176 320424 162182 320436
rect 165614 320424 165620 320436
rect 165672 320424 165678 320476
rect 85574 318112 85580 318164
rect 85632 318152 85638 318164
rect 88334 318152 88340 318164
rect 85632 318124 88340 318152
rect 85632 318112 85638 318124
rect 88334 318112 88340 318124
rect 88392 318112 88398 318164
rect 62758 313896 62764 313948
rect 62816 313936 62822 313948
rect 104894 313936 104900 313948
rect 62816 313908 104900 313936
rect 62816 313896 62822 313908
rect 104894 313896 104900 313908
rect 104952 313896 104958 313948
rect 79318 313352 79324 313404
rect 79376 313392 79382 313404
rect 85574 313392 85580 313404
rect 79376 313364 85580 313392
rect 79376 313352 79382 313364
rect 85574 313352 85580 313364
rect 85632 313352 85638 313404
rect 397086 311856 397092 311908
rect 397144 311896 397150 311908
rect 561950 311896 561956 311908
rect 397144 311868 561956 311896
rect 397144 311856 397150 311868
rect 561950 311856 561956 311868
rect 562008 311856 562014 311908
rect 562226 311856 562232 311908
rect 562284 311896 562290 311908
rect 579982 311896 579988 311908
rect 562284 311868 579988 311896
rect 562284 311856 562290 311868
rect 579982 311856 579988 311868
rect 580040 311856 580046 311908
rect 93118 311516 93124 311568
rect 93176 311556 93182 311568
rect 94498 311556 94504 311568
rect 93176 311528 94504 311556
rect 93176 311516 93182 311528
rect 94498 311516 94504 311528
rect 94556 311516 94562 311568
rect 160094 307776 160100 307828
rect 160152 307816 160158 307828
rect 162118 307816 162124 307828
rect 160152 307788 162124 307816
rect 160152 307776 160158 307788
rect 162118 307776 162124 307788
rect 162176 307776 162182 307828
rect 228358 307816 228364 307828
rect 222212 307788 228364 307816
rect 221458 307708 221464 307760
rect 221516 307748 221522 307760
rect 222212 307748 222240 307788
rect 228358 307776 228364 307788
rect 228416 307776 228422 307828
rect 221516 307720 222240 307748
rect 221516 307708 221522 307720
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 24118 305028 24124 305040
rect 3292 305000 24124 305028
rect 3292 304988 3298 305000
rect 24118 304988 24124 305000
rect 24176 304988 24182 305040
rect 51718 304988 51724 305040
rect 51776 305028 51782 305040
rect 53098 305028 53104 305040
rect 51776 305000 53104 305028
rect 51776 304988 51782 305000
rect 53098 304988 53104 305000
rect 53156 304988 53162 305040
rect 157334 304988 157340 305040
rect 157392 305028 157398 305040
rect 160094 305028 160100 305040
rect 157392 305000 160100 305028
rect 157392 304988 157398 305000
rect 160094 304988 160100 305000
rect 160152 304988 160158 305040
rect 155954 302268 155960 302320
rect 156012 302308 156018 302320
rect 157334 302308 157340 302320
rect 156012 302280 157340 302308
rect 156012 302268 156018 302280
rect 157334 302268 157340 302280
rect 157392 302268 157398 302320
rect 46198 302200 46204 302252
rect 46256 302240 46262 302252
rect 48958 302240 48964 302252
rect 46256 302212 48964 302240
rect 46256 302200 46262 302212
rect 48958 302200 48964 302212
rect 49016 302200 49022 302252
rect 155218 302200 155224 302252
rect 155276 302240 155282 302252
rect 157978 302240 157984 302252
rect 155276 302212 157984 302240
rect 155276 302200 155282 302212
rect 157978 302200 157984 302212
rect 158036 302200 158042 302252
rect 57238 301452 57244 301504
rect 57296 301492 57302 301504
rect 79318 301492 79324 301504
rect 57296 301464 79324 301492
rect 57296 301452 57302 301464
rect 79318 301452 79324 301464
rect 79376 301452 79382 301504
rect 61378 301044 61384 301096
rect 61436 301084 61442 301096
rect 62758 301084 62764 301096
rect 61436 301056 62764 301084
rect 61436 301044 61442 301056
rect 62758 301044 62764 301056
rect 62816 301044 62822 301096
rect 556062 300840 556068 300892
rect 556120 300880 556126 300892
rect 566550 300880 566556 300892
rect 556120 300852 566556 300880
rect 556120 300840 556126 300852
rect 566550 300840 566556 300852
rect 566608 300840 566614 300892
rect 66898 300160 66904 300212
rect 66956 300200 66962 300212
rect 68278 300200 68284 300212
rect 66956 300172 68284 300200
rect 66956 300160 66962 300172
rect 68278 300160 68284 300172
rect 68336 300160 68342 300212
rect 220078 299412 220084 299464
rect 220136 299452 220142 299464
rect 221458 299452 221464 299464
rect 220136 299424 221464 299452
rect 220136 299412 220142 299424
rect 221458 299412 221464 299424
rect 221516 299412 221522 299464
rect 552658 298732 552664 298784
rect 552716 298772 552722 298784
rect 579982 298772 579988 298784
rect 552716 298744 579988 298772
rect 552716 298732 552722 298744
rect 579982 298732 579988 298744
rect 580040 298732 580046 298784
rect 151998 298528 152004 298580
rect 152056 298568 152062 298580
rect 155862 298568 155868 298580
rect 152056 298540 155868 298568
rect 152056 298528 152062 298540
rect 155862 298528 155868 298540
rect 155920 298528 155926 298580
rect 150434 295944 150440 295996
rect 150492 295984 150498 295996
rect 155218 295984 155224 295996
rect 150492 295956 155224 295984
rect 150492 295944 150498 295956
rect 155218 295944 155224 295956
rect 155276 295944 155282 295996
rect 151078 294040 151084 294092
rect 151136 294080 151142 294092
rect 151998 294080 152004 294092
rect 151136 294052 152004 294080
rect 151136 294040 151142 294052
rect 151998 294040 152004 294052
rect 152056 294040 152062 294092
rect 3234 292544 3240 292596
rect 3292 292584 3298 292596
rect 29730 292584 29736 292596
rect 3292 292556 29736 292584
rect 3292 292544 3298 292556
rect 29730 292544 29736 292556
rect 29788 292544 29794 292596
rect 146938 292544 146944 292596
rect 146996 292584 147002 292596
rect 150434 292584 150440 292596
rect 146996 292556 150440 292584
rect 146996 292544 147002 292556
rect 150434 292544 150440 292556
rect 150492 292544 150498 292596
rect 91830 289756 91836 289808
rect 91888 289796 91894 289808
rect 93118 289796 93124 289808
rect 91888 289768 93124 289796
rect 91888 289756 91894 289768
rect 93118 289756 93124 289768
rect 93176 289756 93182 289808
rect 55858 288328 55864 288380
rect 55916 288368 55922 288380
rect 57238 288368 57244 288380
rect 55916 288340 57244 288368
rect 55916 288328 55922 288340
rect 57238 288328 57244 288340
rect 57296 288328 57302 288380
rect 556154 285608 556160 285660
rect 556212 285648 556218 285660
rect 579982 285648 579988 285660
rect 556212 285620 579988 285648
rect 556212 285608 556218 285620
rect 579982 285608 579988 285620
rect 580040 285608 580046 285660
rect 135898 282140 135904 282192
rect 135956 282180 135962 282192
rect 146938 282180 146944 282192
rect 135956 282152 146944 282180
rect 135956 282140 135962 282152
rect 146938 282140 146944 282152
rect 146996 282140 147002 282192
rect 59998 280780 60004 280832
rect 60056 280820 60062 280832
rect 61378 280820 61384 280832
rect 60056 280792 61384 280820
rect 60056 280780 60062 280792
rect 61378 280780 61384 280792
rect 61436 280780 61442 280832
rect 91830 280208 91836 280220
rect 89732 280180 91836 280208
rect 88978 280100 88984 280152
rect 89036 280140 89042 280152
rect 89732 280140 89760 280180
rect 91830 280168 91836 280180
rect 91888 280168 91894 280220
rect 89036 280112 89760 280140
rect 89036 280100 89042 280112
rect 218054 274728 218060 274780
rect 218112 274768 218118 274780
rect 220078 274768 220084 274780
rect 218112 274740 220084 274768
rect 218112 274728 218118 274740
rect 220078 274728 220084 274740
rect 220136 274728 220142 274780
rect 57974 274660 57980 274712
rect 58032 274700 58038 274712
rect 59998 274700 60004 274712
rect 58032 274672 60004 274700
rect 58032 274660 58038 274672
rect 59998 274660 60004 274672
rect 60056 274660 60062 274712
rect 45370 273164 45376 273216
rect 45428 273204 45434 273216
rect 46198 273204 46204 273216
rect 45428 273176 46204 273204
rect 45428 273164 45434 273176
rect 46198 273164 46204 273176
rect 46256 273164 46262 273216
rect 54478 272892 54484 272944
rect 54536 272932 54542 272944
rect 55858 272932 55864 272944
rect 54536 272904 55864 272932
rect 54536 272892 54542 272904
rect 55858 272892 55864 272904
rect 55916 272892 55922 272944
rect 396994 271872 397000 271924
rect 397052 271912 397058 271924
rect 579982 271912 579988 271924
rect 397052 271884 579988 271912
rect 397052 271872 397058 271884
rect 579982 271872 579988 271884
rect 580040 271872 580046 271924
rect 215938 271056 215944 271108
rect 215996 271096 216002 271108
rect 218054 271096 218060 271108
rect 215996 271068 218060 271096
rect 215996 271056 216002 271068
rect 218054 271056 218060 271068
rect 218112 271056 218118 271108
rect 52362 269084 52368 269136
rect 52420 269124 52426 269136
rect 57882 269124 57888 269136
rect 52420 269096 57888 269124
rect 52420 269084 52426 269096
rect 57882 269084 57888 269096
rect 57940 269084 57946 269136
rect 149054 269016 149060 269068
rect 149112 269056 149118 269068
rect 151078 269056 151084 269068
rect 149112 269028 151084 269056
rect 149112 269016 149118 269028
rect 151078 269016 151084 269028
rect 151136 269016 151142 269068
rect 51074 266364 51080 266416
rect 51132 266404 51138 266416
rect 54478 266404 54484 266416
rect 51132 266376 54484 266404
rect 51132 266364 51138 266376
rect 54478 266364 54484 266376
rect 54536 266364 54542 266416
rect 63494 266364 63500 266416
rect 63552 266404 63558 266416
rect 66898 266404 66904 266416
rect 63552 266376 66904 266404
rect 63552 266364 63558 266376
rect 66898 266364 66904 266376
rect 66956 266364 66962 266416
rect 146938 262896 146944 262948
rect 146996 262936 147002 262948
rect 149054 262936 149060 262948
rect 146996 262908 149060 262936
rect 146996 262896 147002 262908
rect 149054 262896 149060 262908
rect 149112 262896 149118 262948
rect 50338 262828 50344 262880
rect 50396 262868 50402 262880
rect 63494 262868 63500 262880
rect 50396 262840 63500 262868
rect 50396 262828 50402 262840
rect 63494 262828 63500 262840
rect 63552 262828 63558 262880
rect 121454 262828 121460 262880
rect 121512 262868 121518 262880
rect 135898 262868 135904 262880
rect 121512 262840 135904 262868
rect 121512 262828 121518 262840
rect 135898 262828 135904 262840
rect 135956 262828 135962 262880
rect 50890 261196 50896 261248
rect 50948 261236 50954 261248
rect 52362 261236 52368 261248
rect 50948 261208 52368 261236
rect 50948 261196 50954 261208
rect 52362 261196 52368 261208
rect 52420 261196 52426 261248
rect 47578 260448 47584 260500
rect 47636 260488 47642 260500
rect 51074 260488 51080 260500
rect 47636 260460 51080 260488
rect 47636 260448 47642 260460
rect 51074 260448 51080 260460
rect 51132 260448 51138 260500
rect 49234 258952 49240 259004
rect 49292 258992 49298 259004
rect 50890 258992 50896 259004
rect 49292 258964 50896 258992
rect 49292 258952 49298 258964
rect 50890 258952 50896 258964
rect 50948 258952 50954 259004
rect 81710 258680 81716 258732
rect 81768 258720 81774 258732
rect 88978 258720 88984 258732
rect 81768 258692 88984 258720
rect 81768 258680 81774 258692
rect 88978 258680 88984 258692
rect 89036 258680 89042 258732
rect 117222 258680 117228 258732
rect 117280 258720 117286 258732
rect 121454 258720 121460 258732
rect 117280 258692 121460 258720
rect 117280 258680 117286 258692
rect 121454 258680 121460 258692
rect 121512 258680 121518 258732
rect 397178 258068 397184 258120
rect 397236 258108 397242 258120
rect 579982 258108 579988 258120
rect 397236 258080 579988 258108
rect 397236 258068 397242 258080
rect 579982 258068 579988 258080
rect 580040 258068 580046 258120
rect 47486 256708 47492 256760
rect 47544 256748 47550 256760
rect 49234 256748 49240 256760
rect 47544 256720 49240 256748
rect 47544 256708 47550 256720
rect 49234 256708 49240 256720
rect 49292 256708 49298 256760
rect 215938 256748 215944 256760
rect 212552 256720 215944 256748
rect 210418 256640 210424 256692
rect 210476 256680 210482 256692
rect 212552 256680 212580 256720
rect 215938 256708 215944 256720
rect 215996 256708 216002 256760
rect 210476 256652 212580 256680
rect 210476 256640 210482 256652
rect 3142 253920 3148 253972
rect 3200 253960 3206 253972
rect 22738 253960 22744 253972
rect 3200 253932 22744 253960
rect 3200 253920 3206 253932
rect 22738 253920 22744 253932
rect 22796 253920 22802 253972
rect 45830 253920 45836 253972
rect 45888 253960 45894 253972
rect 47486 253960 47492 253972
rect 45888 253932 47492 253960
rect 45888 253920 45894 253932
rect 47486 253920 47492 253932
rect 47544 253920 47550 253972
rect 79318 253920 79324 253972
rect 79376 253960 79382 253972
rect 81710 253960 81716 253972
rect 79376 253932 81716 253960
rect 79376 253920 79382 253932
rect 81710 253920 81716 253932
rect 81768 253920 81774 253972
rect 113818 253920 113824 253972
rect 113876 253960 113882 253972
rect 117222 253960 117228 253972
rect 113876 253932 117228 253960
rect 113876 253920 113882 253932
rect 117222 253920 117228 253932
rect 117280 253920 117286 253972
rect 145558 253920 145564 253972
rect 145616 253960 145622 253972
rect 146938 253960 146944 253972
rect 145616 253932 146944 253960
rect 145616 253920 145622 253932
rect 146938 253920 146944 253932
rect 146996 253920 147002 253972
rect 209038 253920 209044 253972
rect 209096 253960 209102 253972
rect 210418 253960 210424 253972
rect 209096 253932 210424 253960
rect 209096 253920 209102 253932
rect 210418 253920 210424 253932
rect 210476 253920 210482 253972
rect 48682 252560 48688 252612
rect 48740 252600 48746 252612
rect 50338 252600 50344 252612
rect 48740 252572 50344 252600
rect 48740 252560 48746 252572
rect 50338 252560 50344 252572
rect 50396 252560 50402 252612
rect 47670 251812 47676 251864
rect 47728 251852 47734 251864
rect 71774 251852 71780 251864
rect 47728 251824 71780 251852
rect 47728 251812 47734 251824
rect 71774 251812 71780 251824
rect 71832 251812 71838 251864
rect 46934 249432 46940 249484
rect 46992 249472 46998 249484
rect 48682 249472 48688 249484
rect 46992 249444 48688 249472
rect 46992 249432 46998 249444
rect 48682 249432 48688 249444
rect 48740 249432 48746 249484
rect 97258 247664 97264 247716
rect 97316 247704 97322 247716
rect 113818 247704 113824 247716
rect 97316 247676 113824 247704
rect 97316 247664 97322 247676
rect 113818 247664 113824 247676
rect 113876 247664 113882 247716
rect 76190 247052 76196 247104
rect 76248 247092 76254 247104
rect 79318 247092 79324 247104
rect 76248 247064 79324 247092
rect 76248 247052 76254 247064
rect 79318 247052 79324 247064
rect 79376 247052 79382 247104
rect 143166 247052 143172 247104
rect 143224 247092 143230 247104
rect 145558 247092 145564 247104
rect 143224 247064 145564 247092
rect 143224 247052 143230 247064
rect 145558 247052 145564 247064
rect 145616 247052 145622 247104
rect 49694 245624 49700 245676
rect 49752 245664 49758 245676
rect 51718 245664 51724 245676
rect 49752 245636 51724 245664
rect 49752 245624 49758 245636
rect 51718 245624 51724 245636
rect 51776 245624 51782 245676
rect 413278 244264 413284 244316
rect 413336 244304 413342 244316
rect 579982 244304 579988 244316
rect 413336 244276 579988 244304
rect 413336 244264 413342 244276
rect 579982 244264 579988 244276
rect 580040 244264 580046 244316
rect 143166 242944 143172 242956
rect 138032 242916 143172 242944
rect 136082 242836 136088 242888
rect 136140 242876 136146 242888
rect 138032 242876 138060 242916
rect 143166 242904 143172 242916
rect 143224 242904 143230 242956
rect 136140 242848 138060 242876
rect 136140 242836 136146 242848
rect 45186 242224 45192 242276
rect 45244 242264 45250 242276
rect 46934 242264 46940 242276
rect 45244 242236 46940 242264
rect 45244 242224 45250 242236
rect 46934 242224 46940 242236
rect 46992 242224 46998 242276
rect 45830 241408 45836 241460
rect 45888 241448 45894 241460
rect 49602 241448 49608 241460
rect 45888 241420 49608 241448
rect 45888 241408 45894 241420
rect 49602 241408 49608 241420
rect 49660 241408 49666 241460
rect 45554 241340 45560 241392
rect 45612 241380 45618 241392
rect 47670 241380 47676 241392
rect 45612 241352 47676 241380
rect 45612 241340 45618 241352
rect 47670 241340 47676 241352
rect 47728 241340 47734 241392
rect 45646 241272 45652 241324
rect 45704 241312 45710 241324
rect 47578 241312 47584 241324
rect 45704 241284 47584 241312
rect 45704 241272 45710 241284
rect 47578 241272 47584 241284
rect 47636 241272 47642 241324
rect 46842 240864 46848 240916
rect 46900 240904 46906 240916
rect 76190 240904 76196 240916
rect 46900 240876 76196 240904
rect 46900 240864 46906 240876
rect 76190 240864 76196 240876
rect 76248 240864 76254 240916
rect 45370 240796 45376 240848
rect 45428 240836 45434 240848
rect 136082 240836 136088 240848
rect 45428 240808 136088 240836
rect 45428 240796 45434 240808
rect 136082 240796 136088 240808
rect 136140 240796 136146 240848
rect 45002 240728 45008 240780
rect 45060 240768 45066 240780
rect 209038 240768 209044 240780
rect 45060 240740 209044 240768
rect 45060 240728 45066 240740
rect 209038 240728 209044 240740
rect 209096 240728 209102 240780
rect 3050 240116 3056 240168
rect 3108 240156 3114 240168
rect 44818 240156 44824 240168
rect 3108 240128 44824 240156
rect 3108 240116 3114 240128
rect 44818 240116 44824 240128
rect 44876 240116 44882 240168
rect 395430 240048 395436 240100
rect 395488 240088 395494 240100
rect 396534 240088 396540 240100
rect 395488 240060 396540 240088
rect 395488 240048 395494 240060
rect 396534 240048 396540 240060
rect 396592 240048 396598 240100
rect 44726 239708 44732 239760
rect 44784 239748 44790 239760
rect 46842 239748 46848 239760
rect 44784 239720 46848 239748
rect 44784 239708 44790 239720
rect 46842 239708 46848 239720
rect 46900 239708 46906 239760
rect 45462 239368 45468 239420
rect 45520 239408 45526 239420
rect 97258 239408 97264 239420
rect 45520 239380 97264 239408
rect 45520 239368 45526 239380
rect 97258 239368 97264 239380
rect 97316 239368 97322 239420
rect 396534 238824 396540 238876
rect 396592 238824 396598 238876
rect 44910 238756 44916 238808
rect 44968 238796 44974 238808
rect 45738 238796 45744 238808
rect 44968 238768 45744 238796
rect 44968 238756 44974 238768
rect 45738 238756 45744 238768
rect 45796 238756 45802 238808
rect 396552 238796 396580 238824
rect 396046 238768 396580 238796
rect 396046 238728 396074 238768
rect 396534 238728 396540 238740
rect 396046 238700 396540 238728
rect 396534 238688 396540 238700
rect 396592 238688 396598 238740
rect 54864 233056 60734 233084
rect 44910 232908 44916 232960
rect 44968 232948 44974 232960
rect 54864 232948 54892 233056
rect 60706 233016 60734 233056
rect 60706 232988 64874 233016
rect 44968 232920 54892 232948
rect 54956 232920 57284 232948
rect 44968 232908 44974 232920
rect 45830 232840 45836 232892
rect 45888 232880 45894 232892
rect 54956 232880 54984 232920
rect 45888 232852 54984 232880
rect 57256 232880 57284 232920
rect 57256 232852 64184 232880
rect 45888 232840 45894 232852
rect 45002 232772 45008 232824
rect 45060 232812 45066 232824
rect 45738 232812 45744 232824
rect 45060 232784 45744 232812
rect 45060 232772 45066 232784
rect 45738 232772 45744 232784
rect 45796 232772 45802 232824
rect 64156 232416 64184 232852
rect 64138 232364 64144 232416
rect 64196 232364 64202 232416
rect 64846 232404 64874 232988
rect 85758 232404 85764 232416
rect 64846 232376 85764 232404
rect 85758 232364 85764 232376
rect 85816 232364 85822 232416
rect 394694 232092 394700 232144
rect 394752 232132 394758 232144
rect 396534 232132 396540 232144
rect 394752 232104 396540 232132
rect 394752 232092 394758 232104
rect 396534 232092 396540 232104
rect 396592 232092 396598 232144
rect 45278 231888 45284 231940
rect 45336 231928 45342 231940
rect 46842 231928 46848 231940
rect 45336 231900 46848 231928
rect 45336 231888 45342 231900
rect 46842 231888 46848 231900
rect 46900 231888 46906 231940
rect 45370 231820 45376 231872
rect 45428 231820 45434 231872
rect 45462 231820 45468 231872
rect 45520 231860 45526 231872
rect 46658 231860 46664 231872
rect 45520 231832 46664 231860
rect 45520 231820 45526 231832
rect 46658 231820 46664 231832
rect 46716 231820 46722 231872
rect 520918 231820 520924 231872
rect 520976 231860 520982 231872
rect 579798 231860 579804 231872
rect 520976 231832 579804 231860
rect 520976 231820 520982 231832
rect 579798 231820 579804 231832
rect 579856 231820 579862 231872
rect 45388 231792 45416 231820
rect 48314 231792 48320 231804
rect 45388 231764 48320 231792
rect 48314 231752 48320 231764
rect 48372 231752 48378 231804
rect 45186 231072 45192 231124
rect 45244 231112 45250 231124
rect 60734 231112 60740 231124
rect 45244 231084 60740 231112
rect 45244 231072 45250 231084
rect 60734 231072 60740 231084
rect 60792 231072 60798 231124
rect 85758 230664 85764 230716
rect 85816 230704 85822 230716
rect 93762 230704 93768 230716
rect 85816 230676 93768 230704
rect 85816 230664 85822 230676
rect 93762 230664 93768 230676
rect 93820 230664 93826 230716
rect 390830 230460 390836 230512
rect 390888 230500 390894 230512
rect 394694 230500 394700 230512
rect 390888 230472 394700 230500
rect 390888 230460 390894 230472
rect 394694 230460 394700 230472
rect 394752 230460 394758 230512
rect 45738 230392 45744 230444
rect 45796 230432 45802 230444
rect 51902 230432 51908 230444
rect 45796 230404 51908 230432
rect 45796 230392 45802 230404
rect 51902 230392 51908 230404
rect 51960 230392 51966 230444
rect 60734 230120 60740 230172
rect 60792 230160 60798 230172
rect 62758 230160 62764 230172
rect 60792 230132 62764 230160
rect 60792 230120 60798 230132
rect 62758 230120 62764 230132
rect 62816 230120 62822 230172
rect 167638 229712 167644 229764
rect 167696 229752 167702 229764
rect 176654 229752 176660 229764
rect 167696 229724 176660 229752
rect 167696 229712 167702 229724
rect 176654 229712 176660 229724
rect 176712 229712 176718 229764
rect 48314 229100 48320 229152
rect 48372 229140 48378 229152
rect 48372 229112 51074 229140
rect 48372 229100 48378 229112
rect 46658 229032 46664 229084
rect 46716 229072 46722 229084
rect 48222 229072 48228 229084
rect 46716 229044 48228 229072
rect 46716 229032 46722 229044
rect 48222 229032 48228 229044
rect 48280 229032 48286 229084
rect 51046 229072 51074 229112
rect 55858 229072 55864 229084
rect 51046 229044 55864 229072
rect 55858 229032 55864 229044
rect 55916 229032 55922 229084
rect 157978 228420 157984 228472
rect 158036 228460 158042 228472
rect 266538 228460 266544 228472
rect 158036 228432 266544 228460
rect 158036 228420 158042 228432
rect 266538 228420 266544 228432
rect 266596 228420 266602 228472
rect 297358 228420 297364 228472
rect 297416 228460 297422 228472
rect 327074 228460 327080 228472
rect 297416 228432 327080 228460
rect 297416 228420 297422 228432
rect 327074 228420 327080 228432
rect 327132 228420 327138 228472
rect 366358 228420 366364 228472
rect 366416 228460 366422 228472
rect 380158 228460 380164 228472
rect 366416 228432 380164 228460
rect 366416 228420 366422 228432
rect 380158 228420 380164 228432
rect 380216 228420 380222 228472
rect 117222 228352 117228 228404
rect 117280 228392 117286 228404
rect 138658 228392 138664 228404
rect 117280 228364 138664 228392
rect 117280 228352 117286 228364
rect 138658 228352 138664 228364
rect 138716 228352 138722 228404
rect 236638 228352 236644 228404
rect 236696 228392 236702 228404
rect 386506 228392 386512 228404
rect 236696 228364 386512 228392
rect 236696 228352 236702 228364
rect 386506 228352 386512 228364
rect 386564 228352 386570 228404
rect 51902 227740 51908 227792
rect 51960 227780 51966 227792
rect 51960 227752 52500 227780
rect 51960 227740 51966 227752
rect 44726 227672 44732 227724
rect 44784 227712 44790 227724
rect 46198 227712 46204 227724
rect 44784 227684 46204 227712
rect 44784 227672 44790 227684
rect 46198 227672 46204 227684
rect 46256 227672 46262 227724
rect 52472 227712 52500 227752
rect 387058 227740 387064 227792
rect 387116 227780 387122 227792
rect 392578 227780 392584 227792
rect 387116 227752 392584 227780
rect 387116 227740 387122 227752
rect 392578 227740 392584 227752
rect 392636 227740 392642 227792
rect 59998 227712 60004 227724
rect 52472 227684 60004 227712
rect 59998 227672 60004 227684
rect 60056 227672 60062 227724
rect 64138 227060 64144 227112
rect 64196 227100 64202 227112
rect 95878 227100 95884 227112
rect 64196 227072 95884 227100
rect 64196 227060 64202 227072
rect 95878 227060 95884 227072
rect 95936 227060 95942 227112
rect 3970 226992 3976 227044
rect 4028 227032 4034 227044
rect 176654 227032 176660 227044
rect 4028 227004 176660 227032
rect 4028 226992 4034 227004
rect 176654 226992 176660 227004
rect 176712 226992 176718 227044
rect 93854 226448 93860 226500
rect 93912 226488 93918 226500
rect 97994 226488 98000 226500
rect 93912 226460 98000 226488
rect 93912 226448 93918 226460
rect 97994 226448 98000 226460
rect 98052 226448 98058 226500
rect 390830 226352 390836 226364
rect 386432 226324 390836 226352
rect 384942 226244 384948 226296
rect 385000 226284 385006 226296
rect 386432 226284 386460 226324
rect 390830 226312 390836 226324
rect 390888 226312 390894 226364
rect 385000 226256 386460 226284
rect 385000 226244 385006 226256
rect 46934 224340 46940 224392
rect 46992 224380 46998 224392
rect 50338 224380 50344 224392
rect 46992 224352 50344 224380
rect 46992 224340 46998 224352
rect 50338 224340 50344 224352
rect 50396 224340 50402 224392
rect 55858 224136 55864 224188
rect 55916 224176 55922 224188
rect 57238 224176 57244 224188
rect 55916 224148 57244 224176
rect 55916 224136 55922 224148
rect 57238 224136 57244 224148
rect 57296 224136 57302 224188
rect 59998 224136 60004 224188
rect 60056 224176 60062 224188
rect 62114 224176 62120 224188
rect 60056 224148 62120 224176
rect 60056 224136 60062 224148
rect 62114 224136 62120 224148
rect 62172 224136 62178 224188
rect 97994 224136 98000 224188
rect 98052 224176 98058 224188
rect 100018 224176 100024 224188
rect 98052 224148 100024 224176
rect 98052 224136 98058 224148
rect 100018 224136 100024 224148
rect 100076 224136 100082 224188
rect 384942 223632 384948 223644
rect 383626 223604 384948 223632
rect 380894 223524 380900 223576
rect 380952 223564 380958 223576
rect 383626 223564 383654 223604
rect 384942 223592 384948 223604
rect 385000 223592 385006 223644
rect 380952 223536 383654 223564
rect 380952 223524 380958 223536
rect 46198 223252 46204 223304
rect 46256 223292 46262 223304
rect 47670 223292 47676 223304
rect 46256 223264 47676 223292
rect 46256 223252 46262 223264
rect 47670 223252 47676 223264
rect 47728 223252 47734 223304
rect 48222 222096 48228 222148
rect 48280 222136 48286 222148
rect 51442 222136 51448 222148
rect 48280 222108 51448 222136
rect 48280 222096 48286 222108
rect 51442 222096 51448 222108
rect 51500 222096 51506 222148
rect 62758 221416 62764 221468
rect 62816 221456 62822 221468
rect 69014 221456 69020 221468
rect 62816 221428 69020 221456
rect 62816 221416 62822 221428
rect 69014 221416 69020 221428
rect 69072 221416 69078 221468
rect 372614 221416 372620 221468
rect 372672 221456 372678 221468
rect 380894 221456 380900 221468
rect 372672 221428 380900 221456
rect 372672 221416 372678 221428
rect 380894 221416 380900 221428
rect 380952 221416 380958 221468
rect 62114 221212 62120 221264
rect 62172 221252 62178 221264
rect 66254 221252 66260 221264
rect 62172 221224 66260 221252
rect 62172 221212 62178 221224
rect 66254 221212 66260 221224
rect 66312 221212 66318 221264
rect 45094 221076 45100 221128
rect 45152 221116 45158 221128
rect 46934 221116 46940 221128
rect 45152 221088 46940 221116
rect 45152 221076 45158 221088
rect 46934 221076 46940 221088
rect 46992 221076 46998 221128
rect 369854 220396 369860 220448
rect 369912 220436 369918 220448
rect 372614 220436 372620 220448
rect 369912 220408 372620 220436
rect 369912 220396 369918 220408
rect 372614 220396 372620 220408
rect 372672 220396 372678 220448
rect 69014 219444 69020 219496
rect 69072 219484 69078 219496
rect 69072 219456 70440 219484
rect 69072 219444 69078 219456
rect 70412 219416 70440 219456
rect 72418 219416 72424 219428
rect 70412 219388 72424 219416
rect 72418 219376 72424 219388
rect 72476 219376 72482 219428
rect 95878 218696 95884 218748
rect 95936 218736 95942 218748
rect 106182 218736 106188 218748
rect 95936 218708 106188 218736
rect 95936 218696 95942 218708
rect 106182 218696 106188 218708
rect 106240 218696 106246 218748
rect 379514 218696 379520 218748
rect 379572 218736 379578 218748
rect 387058 218736 387064 218748
rect 379572 218708 387064 218736
rect 379572 218696 379578 218708
rect 387058 218696 387064 218708
rect 387116 218696 387122 218748
rect 47670 218016 47676 218068
rect 47728 218056 47734 218068
rect 47728 218028 48360 218056
rect 47728 218016 47734 218028
rect 48332 217988 48360 218028
rect 115842 218016 115848 218068
rect 115900 218056 115906 218068
rect 579798 218056 579804 218068
rect 115900 218028 579804 218056
rect 115900 218016 115906 218028
rect 579798 218016 579804 218028
rect 579856 218016 579862 218068
rect 53834 217988 53840 218000
rect 48332 217960 53840 217988
rect 53834 217948 53840 217960
rect 53892 217948 53898 218000
rect 100018 217948 100024 218000
rect 100076 217988 100082 218000
rect 105998 217988 106004 218000
rect 100076 217960 106004 217988
rect 100076 217948 100082 217960
rect 105998 217948 106004 217960
rect 106056 217948 106062 218000
rect 45646 217268 45652 217320
rect 45704 217308 45710 217320
rect 58250 217308 58256 217320
rect 45704 217280 58256 217308
rect 45704 217268 45710 217280
rect 58250 217268 58256 217280
rect 58308 217268 58314 217320
rect 46934 216656 46940 216708
rect 46992 216696 46998 216708
rect 51718 216696 51724 216708
rect 46992 216668 51724 216696
rect 46992 216656 46998 216668
rect 51718 216656 51724 216668
rect 51776 216656 51782 216708
rect 66254 216656 66260 216708
rect 66312 216696 66318 216708
rect 68278 216696 68284 216708
rect 66312 216668 68284 216696
rect 66312 216656 66318 216668
rect 68278 216656 68284 216668
rect 68336 216656 68342 216708
rect 369854 216696 369860 216708
rect 368492 216668 369860 216696
rect 366450 216588 366456 216640
rect 366508 216628 366514 216640
rect 368492 216628 368520 216668
rect 369854 216656 369860 216668
rect 369912 216656 369918 216708
rect 366508 216600 368520 216628
rect 366508 216588 366514 216600
rect 57238 215772 57244 215824
rect 57296 215812 57302 215824
rect 58710 215812 58716 215824
rect 57296 215784 58716 215812
rect 57296 215772 57302 215784
rect 58710 215772 58716 215784
rect 58768 215772 58774 215824
rect 105998 215296 106004 215348
rect 106056 215336 106062 215348
rect 106056 215308 107700 215336
rect 106056 215296 106062 215308
rect 72418 215228 72424 215280
rect 72476 215268 72482 215280
rect 75178 215268 75184 215280
rect 72476 215240 75184 215268
rect 72476 215228 72482 215240
rect 75178 215228 75184 215240
rect 75236 215228 75242 215280
rect 107672 215268 107700 215308
rect 110414 215268 110420 215280
rect 107672 215240 110420 215268
rect 110414 215228 110420 215240
rect 110472 215228 110478 215280
rect 106182 214616 106188 214668
rect 106240 214656 106246 214668
rect 107838 214656 107844 214668
rect 106240 214628 107844 214656
rect 106240 214616 106246 214628
rect 107838 214616 107844 214628
rect 107896 214616 107902 214668
rect 3142 213936 3148 213988
rect 3200 213976 3206 213988
rect 176746 213976 176752 213988
rect 3200 213948 176752 213976
rect 3200 213936 3206 213948
rect 176746 213936 176752 213948
rect 176804 213936 176810 213988
rect 51442 213868 51448 213920
rect 51500 213908 51506 213920
rect 54478 213908 54484 213920
rect 51500 213880 54484 213908
rect 51500 213868 51506 213880
rect 54478 213868 54484 213880
rect 54536 213868 54542 213920
rect 58710 213868 58716 213920
rect 58768 213908 58774 213920
rect 59998 213908 60004 213920
rect 58768 213880 60004 213908
rect 58768 213868 58774 213880
rect 59998 213868 60004 213880
rect 60056 213868 60062 213920
rect 58250 212440 58256 212492
rect 58308 212480 58314 212492
rect 61930 212480 61936 212492
rect 58308 212452 61936 212480
rect 58308 212440 58314 212452
rect 61930 212440 61936 212452
rect 61988 212440 61994 212492
rect 375282 211896 375288 211948
rect 375340 211936 375346 211948
rect 379422 211936 379428 211948
rect 375340 211908 379428 211936
rect 375340 211896 375346 211908
rect 379422 211896 379428 211908
rect 379480 211896 379486 211948
rect 53834 211148 53840 211200
rect 53892 211188 53898 211200
rect 53892 211160 55214 211188
rect 53892 211148 53898 211160
rect 55186 211120 55214 211160
rect 56686 211120 56692 211132
rect 55186 211092 56692 211120
rect 56686 211080 56692 211092
rect 56744 211080 56750 211132
rect 110414 210468 110420 210520
rect 110472 210508 110478 210520
rect 113174 210508 113180 210520
rect 110472 210480 113180 210508
rect 110472 210468 110478 210480
rect 113174 210468 113180 210480
rect 113232 210468 113238 210520
rect 107838 210400 107844 210452
rect 107896 210440 107902 210452
rect 116578 210440 116584 210452
rect 107896 210412 116584 210440
rect 107896 210400 107902 210412
rect 116578 210400 116584 210412
rect 116636 210400 116642 210452
rect 371142 209788 371148 209840
rect 371200 209828 371206 209840
rect 375282 209828 375288 209840
rect 371200 209800 375288 209828
rect 371200 209788 371206 209800
rect 375282 209788 375288 209800
rect 375340 209788 375346 209840
rect 382918 209040 382924 209092
rect 382976 209080 382982 209092
rect 397546 209080 397552 209092
rect 382976 209052 397552 209080
rect 382976 209040 382982 209052
rect 397546 209040 397552 209052
rect 397604 209040 397610 209092
rect 54478 208156 54484 208208
rect 54536 208196 54542 208208
rect 55858 208196 55864 208208
rect 54536 208168 55864 208196
rect 54536 208156 54542 208168
rect 55858 208156 55864 208168
rect 55916 208156 55922 208208
rect 56686 207748 56692 207800
rect 56744 207788 56750 207800
rect 62022 207788 62028 207800
rect 56744 207760 62028 207788
rect 56744 207748 56750 207760
rect 62022 207748 62028 207760
rect 62080 207748 62086 207800
rect 59998 206932 60004 206984
rect 60056 206972 60062 206984
rect 66162 206972 66168 206984
rect 60056 206944 66168 206972
rect 60056 206932 60062 206944
rect 66162 206932 66168 206944
rect 66220 206932 66226 206984
rect 113174 205980 113180 206032
rect 113232 206020 113238 206032
rect 115106 206020 115112 206032
rect 113232 205992 115112 206020
rect 113232 205980 113238 205992
rect 115106 205980 115112 205992
rect 115164 205980 115170 206032
rect 364978 205708 364984 205760
rect 365036 205748 365042 205760
rect 366450 205748 366456 205760
rect 365036 205720 366456 205748
rect 365036 205708 365042 205720
rect 366450 205708 366456 205720
rect 366508 205708 366514 205760
rect 188338 205640 188344 205692
rect 188396 205680 188402 205692
rect 579982 205680 579988 205692
rect 188396 205652 579988 205680
rect 188396 205640 188402 205652
rect 579982 205640 579988 205652
rect 580040 205640 580046 205692
rect 61930 204892 61936 204944
rect 61988 204932 61994 204944
rect 71038 204932 71044 204944
rect 61988 204904 71044 204932
rect 61988 204892 61994 204904
rect 71038 204892 71044 204904
rect 71096 204892 71102 204944
rect 367738 204756 367744 204808
rect 367796 204796 367802 204808
rect 371142 204796 371148 204808
rect 367796 204768 371148 204796
rect 367796 204756 367802 204768
rect 371142 204756 371148 204768
rect 371200 204756 371206 204808
rect 62114 204212 62120 204264
rect 62172 204252 62178 204264
rect 64138 204252 64144 204264
rect 62172 204224 64144 204252
rect 62172 204212 62178 204224
rect 64138 204212 64144 204224
rect 64196 204212 64202 204264
rect 75178 202852 75184 202904
rect 75236 202892 75242 202904
rect 75236 202864 78720 202892
rect 75236 202852 75242 202864
rect 78692 202824 78720 202864
rect 80698 202824 80704 202836
rect 78692 202796 80704 202824
rect 80698 202784 80704 202796
rect 80756 202784 80762 202836
rect 2958 201492 2964 201544
rect 3016 201532 3022 201544
rect 22830 201532 22836 201544
rect 3016 201504 22836 201532
rect 3016 201492 3022 201504
rect 22830 201492 22836 201504
rect 22888 201492 22894 201544
rect 362954 201492 362960 201544
rect 363012 201532 363018 201544
rect 366358 201532 366364 201544
rect 363012 201504 366364 201532
rect 363012 201492 363018 201504
rect 366358 201492 366364 201504
rect 366416 201492 366422 201544
rect 115106 201424 115112 201476
rect 115164 201464 115170 201476
rect 116854 201464 116860 201476
rect 115164 201436 116860 201464
rect 115164 201424 115170 201436
rect 116854 201424 116860 201436
rect 116912 201424 116918 201476
rect 51718 200744 51724 200796
rect 51776 200784 51782 200796
rect 73154 200784 73160 200796
rect 51776 200756 73160 200784
rect 51776 200744 51782 200756
rect 73154 200744 73160 200756
rect 73212 200744 73218 200796
rect 66438 199384 66444 199436
rect 66496 199424 66502 199436
rect 75454 199424 75460 199436
rect 66496 199396 75460 199424
rect 66496 199384 66502 199396
rect 75454 199384 75460 199396
rect 75512 199384 75518 199436
rect 155954 199384 155960 199436
rect 156012 199424 156018 199436
rect 296714 199424 296720 199436
rect 156012 199396 296720 199424
rect 156012 199384 156018 199396
rect 296714 199384 296720 199396
rect 296772 199384 296778 199436
rect 377398 198704 377404 198756
rect 377456 198744 377462 198756
rect 382918 198744 382924 198756
rect 377456 198716 382924 198744
rect 377456 198704 377462 198716
rect 382918 198704 382924 198716
rect 382976 198704 382982 198756
rect 362218 198024 362224 198076
rect 362276 198064 362282 198076
rect 364978 198064 364984 198076
rect 362276 198036 364984 198064
rect 362276 198024 362282 198036
rect 364978 198024 364984 198036
rect 365036 198024 365042 198076
rect 50338 197956 50344 198008
rect 50396 197996 50402 198008
rect 53834 197996 53840 198008
rect 50396 197968 53840 197996
rect 50396 197956 50402 197968
rect 53834 197956 53840 197968
rect 53892 197956 53898 198008
rect 73154 197956 73160 198008
rect 73212 197996 73218 198008
rect 77938 197996 77944 198008
rect 73212 197968 77944 197996
rect 73212 197956 73218 197968
rect 77938 197956 77944 197968
rect 77996 197956 78002 198008
rect 148962 197956 148968 198008
rect 149020 197996 149026 198008
rect 207014 197996 207020 198008
rect 149020 197968 207020 197996
rect 149020 197956 149026 197968
rect 207014 197956 207020 197968
rect 207072 197956 207078 198008
rect 116854 197820 116860 197872
rect 116912 197860 116918 197872
rect 119982 197860 119988 197872
rect 116912 197832 119988 197860
rect 116912 197820 116918 197832
rect 119982 197820 119988 197832
rect 120040 197820 120046 197872
rect 154482 197412 154488 197464
rect 154540 197452 154546 197464
rect 155954 197452 155960 197464
rect 154540 197424 155960 197452
rect 154540 197412 154546 197424
rect 155954 197412 155960 197424
rect 156012 197412 156018 197464
rect 68278 197344 68284 197396
rect 68336 197384 68342 197396
rect 68336 197356 69060 197384
rect 68336 197344 68342 197356
rect 69032 197316 69060 197356
rect 355318 197344 355324 197396
rect 355376 197384 355382 197396
rect 362954 197384 362960 197396
rect 355376 197356 362960 197384
rect 355376 197344 355382 197356
rect 362954 197344 362960 197356
rect 363012 197344 363018 197396
rect 71774 197316 71780 197328
rect 69032 197288 71780 197316
rect 71774 197276 71780 197288
rect 71832 197276 71838 197328
rect 152734 197276 152740 197328
rect 152792 197316 152798 197328
rect 157978 197316 157984 197328
rect 152792 197288 157984 197316
rect 152792 197276 152798 197288
rect 157978 197276 157984 197288
rect 158036 197276 158042 197328
rect 147950 196732 147956 196784
rect 148008 196772 148014 196784
rect 167638 196772 167644 196784
rect 148008 196744 167644 196772
rect 148008 196732 148014 196744
rect 167638 196732 167644 196744
rect 167696 196732 167702 196784
rect 160830 196664 160836 196716
rect 160888 196704 160894 196716
rect 236638 196704 236644 196716
rect 160888 196676 236644 196704
rect 160888 196664 160894 196676
rect 236638 196664 236644 196676
rect 236696 196664 236702 196716
rect 151170 196596 151176 196648
rect 151228 196636 151234 196648
rect 235994 196636 236000 196648
rect 151228 196608 236000 196636
rect 151228 196596 151234 196608
rect 235994 196596 236000 196608
rect 236052 196596 236058 196648
rect 64138 195916 64144 195968
rect 64196 195956 64202 195968
rect 65518 195956 65524 195968
rect 64196 195928 65524 195956
rect 64196 195916 64202 195928
rect 65518 195916 65524 195928
rect 65576 195916 65582 195968
rect 138658 195916 138664 195968
rect 138716 195956 138722 195968
rect 141418 195956 141424 195968
rect 138716 195928 141424 195956
rect 138716 195916 138722 195928
rect 141418 195916 141424 195928
rect 141476 195916 141482 195968
rect 157518 195916 157524 195968
rect 157576 195956 157582 195968
rect 356054 195956 356060 195968
rect 157576 195928 356060 195956
rect 157576 195916 157582 195928
rect 356054 195916 356060 195928
rect 356112 195916 356118 195968
rect 86954 195848 86960 195900
rect 87012 195888 87018 195900
rect 139394 195888 139400 195900
rect 87012 195860 139400 195888
rect 87012 195848 87018 195860
rect 139394 195848 139400 195860
rect 139452 195848 139458 195900
rect 157426 195848 157432 195900
rect 157484 195888 157490 195900
rect 297358 195888 297364 195900
rect 157484 195860 297364 195888
rect 157484 195848 157490 195860
rect 297358 195848 297364 195860
rect 297416 195848 297422 195900
rect 56594 195780 56600 195832
rect 56652 195820 56658 195832
rect 138106 195820 138112 195832
rect 56652 195792 138112 195820
rect 56652 195780 56658 195792
rect 138106 195780 138112 195792
rect 138164 195780 138170 195832
rect 71774 194488 71780 194540
rect 71832 194528 71838 194540
rect 75178 194528 75184 194540
rect 71832 194500 75184 194528
rect 71832 194488 71838 194500
rect 75178 194488 75184 194500
rect 75236 194488 75242 194540
rect 75454 194488 75460 194540
rect 75512 194528 75518 194540
rect 76558 194528 76564 194540
rect 75512 194500 76564 194528
rect 75512 194488 75518 194500
rect 76558 194488 76564 194500
rect 76616 194488 76622 194540
rect 116578 194488 116584 194540
rect 116636 194528 116642 194540
rect 124858 194528 124864 194540
rect 116636 194500 124864 194528
rect 116636 194488 116642 194500
rect 124858 194488 124864 194500
rect 124916 194488 124922 194540
rect 217318 193808 217324 193860
rect 217376 193848 217382 193860
rect 580166 193848 580172 193860
rect 217376 193820 580172 193848
rect 217376 193808 217382 193820
rect 580166 193808 580172 193820
rect 580224 193808 580230 193860
rect 53834 192448 53840 192500
rect 53892 192488 53898 192500
rect 60366 192488 60372 192500
rect 53892 192460 60372 192488
rect 53892 192448 53898 192460
rect 60366 192448 60372 192460
rect 60424 192448 60430 192500
rect 120074 192448 120080 192500
rect 120132 192488 120138 192500
rect 128354 192488 128360 192500
rect 120132 192460 128360 192488
rect 120132 192448 120138 192460
rect 128354 192448 128360 192460
rect 128412 192448 128418 192500
rect 341518 189728 341524 189780
rect 341576 189768 341582 189780
rect 355318 189768 355324 189780
rect 341576 189740 355324 189768
rect 341576 189728 341582 189740
rect 355318 189728 355324 189740
rect 355376 189728 355382 189780
rect 60366 189048 60372 189100
rect 60424 189088 60430 189100
rect 62758 189088 62764 189100
rect 60424 189060 62764 189088
rect 60424 189048 60430 189060
rect 62758 189048 62764 189060
rect 62816 189048 62822 189100
rect 128354 189048 128360 189100
rect 128412 189088 128418 189100
rect 130378 189088 130384 189100
rect 128412 189060 130384 189088
rect 128412 189048 128418 189060
rect 130378 189048 130384 189060
rect 130436 189048 130442 189100
rect 359458 189048 359464 189100
rect 359516 189088 359522 189100
rect 362218 189088 362224 189100
rect 359516 189060 362224 189088
rect 359516 189048 359522 189060
rect 362218 189048 362224 189060
rect 362276 189048 362282 189100
rect 76558 188572 76564 188624
rect 76616 188612 76622 188624
rect 79962 188612 79968 188624
rect 76616 188584 79968 188612
rect 76616 188572 76622 188584
rect 79962 188572 79968 188584
rect 80020 188572 80026 188624
rect 80698 187892 80704 187944
rect 80756 187932 80762 187944
rect 82170 187932 82176 187944
rect 80756 187904 82176 187932
rect 80756 187892 80762 187904
rect 82170 187892 82176 187904
rect 82228 187892 82234 187944
rect 3142 187688 3148 187740
rect 3200 187728 3206 187740
rect 112438 187728 112444 187740
rect 3200 187700 112444 187728
rect 3200 187688 3206 187700
rect 112438 187688 112444 187700
rect 112496 187688 112502 187740
rect 366358 187688 366364 187740
rect 366416 187728 366422 187740
rect 367738 187728 367744 187740
rect 366416 187700 367744 187728
rect 366416 187688 366422 187700
rect 367738 187688 367744 187700
rect 367796 187688 367802 187740
rect 166166 187620 166172 187672
rect 166224 187660 166230 187672
rect 399478 187660 399484 187672
rect 166224 187632 399484 187660
rect 166224 187620 166230 187632
rect 399478 187620 399484 187632
rect 399536 187620 399542 187672
rect 79962 186328 79968 186380
rect 80020 186368 80026 186380
rect 80020 186340 80100 186368
rect 80020 186328 80026 186340
rect 80072 186300 80100 186340
rect 86218 186300 86224 186312
rect 80072 186272 86224 186300
rect 86218 186260 86224 186272
rect 86276 186260 86282 186312
rect 159542 185852 159548 185904
rect 159600 185852 159606 185904
rect 159560 185552 159588 185852
rect 159910 185552 159916 185564
rect 159560 185524 159916 185552
rect 159910 185512 159916 185524
rect 159968 185512 159974 185564
rect 142430 184260 142436 184272
rect 137986 184232 142436 184260
rect 135254 184152 135260 184204
rect 135312 184192 135318 184204
rect 137986 184192 138014 184232
rect 142430 184220 142436 184232
rect 142488 184220 142494 184272
rect 135312 184164 138014 184192
rect 135312 184152 135318 184164
rect 371878 184152 371884 184204
rect 371936 184192 371942 184204
rect 377398 184192 377404 184204
rect 371936 184164 377404 184192
rect 371936 184152 371942 184164
rect 377398 184152 377404 184164
rect 377456 184152 377462 184204
rect 82170 183472 82176 183524
rect 82228 183512 82234 183524
rect 83550 183512 83556 183524
rect 82228 183484 83556 183512
rect 82228 183472 82234 183484
rect 83550 183472 83556 183484
rect 83608 183472 83614 183524
rect 65518 182112 65524 182164
rect 65576 182152 65582 182164
rect 66898 182152 66904 182164
rect 65576 182124 66904 182152
rect 65576 182112 65582 182124
rect 66898 182112 66904 182124
rect 66956 182112 66962 182164
rect 144638 181500 144644 181552
rect 144696 181540 144702 181552
rect 145190 181540 145196 181552
rect 144696 181512 145196 181540
rect 144696 181500 144702 181512
rect 145190 181500 145196 181512
rect 145248 181500 145254 181552
rect 157242 181160 157248 181212
rect 157300 181200 157306 181212
rect 159910 181200 159916 181212
rect 157300 181172 159916 181200
rect 157300 181160 157306 181172
rect 159910 181160 159916 181172
rect 159968 181160 159974 181212
rect 144730 181092 144736 181144
rect 144788 181092 144794 181144
rect 144748 181064 144776 181092
rect 150894 181064 150900 181076
rect 144748 181036 150900 181064
rect 150894 181024 150900 181036
rect 150952 181024 150958 181076
rect 157242 180616 157248 180668
rect 157300 180616 157306 180668
rect 157260 180124 157288 180616
rect 71038 180072 71044 180124
rect 71096 180112 71102 180124
rect 81434 180112 81440 180124
rect 71096 180084 81440 180112
rect 71096 180072 71102 180084
rect 81434 180072 81440 180084
rect 81492 180072 81498 180124
rect 117314 180072 117320 180124
rect 117372 180112 117378 180124
rect 136358 180112 136364 180124
rect 117372 180084 136364 180112
rect 117372 180072 117378 180084
rect 136358 180072 136364 180084
rect 136416 180072 136422 180124
rect 150894 180072 150900 180124
rect 150952 180112 150958 180124
rect 153930 180112 153936 180124
rect 150952 180084 153936 180112
rect 150952 180072 150958 180084
rect 153930 180072 153936 180084
rect 153988 180072 153994 180124
rect 157242 180072 157248 180124
rect 157300 180072 157306 180124
rect 62758 180004 62764 180056
rect 62816 180044 62822 180056
rect 63770 180044 63776 180056
rect 62816 180016 63776 180044
rect 62816 180004 62822 180016
rect 63770 180004 63776 180016
rect 63828 180004 63834 180056
rect 158622 179596 158628 179648
rect 158680 179636 158686 179648
rect 166534 179636 166540 179648
rect 158680 179608 166540 179636
rect 158680 179596 158686 179608
rect 166534 179596 166540 179608
rect 166592 179596 166598 179648
rect 154390 179528 154396 179580
rect 154448 179568 154454 179580
rect 157794 179568 157800 179580
rect 154448 179540 157800 179568
rect 154448 179528 154454 179540
rect 157794 179528 157800 179540
rect 157852 179528 157858 179580
rect 130378 179392 130384 179444
rect 130436 179432 130442 179444
rect 130436 179404 131160 179432
rect 130436 179392 130442 179404
rect 131132 179364 131160 179404
rect 336550 179392 336556 179444
rect 336608 179432 336614 179444
rect 341518 179432 341524 179444
rect 336608 179404 341524 179432
rect 336608 179392 336614 179404
rect 341518 179392 341524 179404
rect 341576 179392 341582 179444
rect 135162 179364 135168 179376
rect 131132 179336 135168 179364
rect 135162 179324 135168 179336
rect 135220 179324 135226 179376
rect 136726 178780 136732 178832
rect 136784 178780 136790 178832
rect 120718 178644 120724 178696
rect 120776 178684 120782 178696
rect 136450 178684 136456 178696
rect 120776 178656 136456 178684
rect 120776 178644 120782 178656
rect 136450 178644 136456 178656
rect 136508 178644 136514 178696
rect 136744 178616 136772 178780
rect 136376 178588 136772 178616
rect 136376 178424 136404 178588
rect 154390 178508 154396 178560
rect 154448 178548 154454 178560
rect 157242 178548 157248 178560
rect 154448 178520 157248 178548
rect 154448 178508 154454 178520
rect 157242 178508 157248 178520
rect 157300 178508 157306 178560
rect 153102 178440 153108 178492
rect 153160 178480 153166 178492
rect 153930 178480 153936 178492
rect 153160 178452 153936 178480
rect 153160 178440 153166 178452
rect 153930 178440 153936 178452
rect 153988 178440 153994 178492
rect 136358 178372 136364 178424
rect 136416 178372 136422 178424
rect 114462 178032 114468 178084
rect 114520 178072 114526 178084
rect 153930 178072 153936 178084
rect 114520 178044 153936 178072
rect 114520 178032 114526 178044
rect 153930 178032 153936 178044
rect 153988 178032 153994 178084
rect 154390 178032 154396 178084
rect 154448 178072 154454 178084
rect 157794 178072 157800 178084
rect 154448 178044 157800 178072
rect 154448 178032 154454 178044
rect 157794 178032 157800 178044
rect 157852 178032 157858 178084
rect 158622 178032 158628 178084
rect 158680 178072 158686 178084
rect 579982 178072 579988 178084
rect 158680 178044 579988 178072
rect 158680 178032 158686 178044
rect 579982 178032 579988 178044
rect 580040 178032 580046 178084
rect 63770 177964 63776 178016
rect 63828 178004 63834 178016
rect 65518 178004 65524 178016
rect 63828 177976 65524 178004
rect 63828 177964 63834 177976
rect 65518 177964 65524 177976
rect 65576 177964 65582 178016
rect 134702 177760 134708 177812
rect 134760 177800 134766 177812
rect 136634 177800 136640 177812
rect 134760 177772 136640 177800
rect 134760 177760 134766 177772
rect 136634 177760 136640 177772
rect 136692 177760 136698 177812
rect 120074 177284 120080 177336
rect 120132 177324 120138 177336
rect 136450 177324 136456 177336
rect 120132 177296 136456 177324
rect 120132 177284 120138 177296
rect 136450 177284 136456 177296
rect 136508 177284 136514 177336
rect 144454 177216 144460 177268
rect 144512 177256 144518 177268
rect 148042 177256 148048 177268
rect 144512 177228 148048 177256
rect 144512 177216 144518 177228
rect 148042 177216 148048 177228
rect 148100 177216 148106 177268
rect 55858 177148 55864 177200
rect 55916 177188 55922 177200
rect 56870 177188 56876 177200
rect 55916 177160 56876 177188
rect 55916 177148 55922 177160
rect 56870 177148 56876 177160
rect 56928 177148 56934 177200
rect 368474 176672 368480 176724
rect 368532 176712 368538 176724
rect 371878 176712 371884 176724
rect 368532 176684 371884 176712
rect 368532 176672 368538 176684
rect 371878 176672 371884 176684
rect 371936 176672 371942 176724
rect 83550 176604 83556 176656
rect 83608 176644 83614 176656
rect 84930 176644 84936 176656
rect 83608 176616 84936 176644
rect 83608 176604 83614 176616
rect 84930 176604 84936 176616
rect 84988 176604 84994 176656
rect 153102 176400 153108 176452
rect 153160 176400 153166 176452
rect 122834 176060 122840 176112
rect 122892 176100 122898 176112
rect 134702 176100 134708 176112
rect 122892 176072 134708 176100
rect 122892 176060 122898 176072
rect 134702 176060 134708 176072
rect 134760 176060 134766 176112
rect 121454 175924 121460 175976
rect 121512 175964 121518 175976
rect 136358 175964 136364 175976
rect 121512 175936 136364 175964
rect 121512 175924 121518 175936
rect 136358 175924 136364 175936
rect 136416 175924 136422 175976
rect 153120 175432 153148 176400
rect 153102 175380 153108 175432
rect 153160 175380 153166 175432
rect 141602 175312 141608 175364
rect 141660 175352 141666 175364
rect 153930 175352 153936 175364
rect 141660 175324 153936 175352
rect 141660 175312 141666 175324
rect 153930 175312 153936 175324
rect 153988 175312 153994 175364
rect 56870 175244 56876 175296
rect 56928 175284 56934 175296
rect 56928 175256 58020 175284
rect 56928 175244 56934 175256
rect 57992 175216 58020 175256
rect 154390 175244 154396 175296
rect 154448 175284 154454 175296
rect 156506 175284 156512 175296
rect 154448 175256 156512 175284
rect 154448 175244 154454 175256
rect 156506 175244 156512 175256
rect 156564 175244 156570 175296
rect 62114 175216 62120 175228
rect 57992 175188 62120 175216
rect 62114 175176 62120 175188
rect 62172 175176 62178 175228
rect 81434 175176 81440 175228
rect 81492 175216 81498 175228
rect 84838 175216 84844 175228
rect 81492 175188 84844 175216
rect 81492 175176 81498 175188
rect 84838 175176 84844 175188
rect 84896 175176 84902 175228
rect 153102 174836 153108 174888
rect 153160 174836 153166 174888
rect 144086 174700 144092 174752
rect 144144 174740 144150 174752
rect 145466 174740 145472 174752
rect 144144 174712 145472 174740
rect 144144 174700 144150 174712
rect 145466 174700 145472 174712
rect 145524 174700 145530 174752
rect 153120 174740 153148 174836
rect 152936 174712 153148 174740
rect 140056 174644 144914 174672
rect 125594 174496 125600 174548
rect 125652 174536 125658 174548
rect 136450 174536 136456 174548
rect 125652 174508 136456 174536
rect 125652 174496 125658 174508
rect 136450 174496 136456 174508
rect 136508 174496 136514 174548
rect 134518 174428 134524 174480
rect 134576 174468 134582 174480
rect 140056 174468 140084 174644
rect 144886 174604 144914 174644
rect 152936 174604 152964 174712
rect 329098 174632 329104 174684
rect 329156 174672 329162 174684
rect 336550 174672 336556 174684
rect 329156 174644 336556 174672
rect 329156 174632 329162 174644
rect 336550 174632 336556 174644
rect 336608 174632 336614 174684
rect 364978 174632 364984 174684
rect 365036 174672 365042 174684
rect 368474 174672 368480 174684
rect 365036 174644 368480 174672
rect 365036 174632 365042 174644
rect 368474 174632 368480 174644
rect 368532 174632 368538 174684
rect 144886 174576 152964 174604
rect 162486 174536 162492 174548
rect 134576 174440 140084 174468
rect 143276 174508 162492 174536
rect 134576 174428 134582 174440
rect 140498 174360 140504 174412
rect 140556 174400 140562 174412
rect 143276 174400 143304 174508
rect 162486 174496 162492 174508
rect 162544 174496 162550 174548
rect 145466 174428 145472 174480
rect 145524 174468 145530 174480
rect 155494 174468 155500 174480
rect 145524 174440 155500 174468
rect 145524 174428 145530 174440
rect 155494 174428 155500 174440
rect 155552 174428 155558 174480
rect 140556 174372 143304 174400
rect 140556 174360 140562 174372
rect 115750 174292 115756 174344
rect 115808 174332 115814 174344
rect 580442 174332 580448 174344
rect 115808 174304 138014 174332
rect 115808 174292 115814 174304
rect 137986 174264 138014 174304
rect 154546 174304 580448 174332
rect 154546 174264 154574 174304
rect 580442 174292 580448 174304
rect 580500 174292 580506 174344
rect 137986 174236 154574 174264
rect 129734 173884 129740 173936
rect 129792 173924 129798 173936
rect 137370 173924 137376 173936
rect 129792 173896 137376 173924
rect 129792 173884 129798 173896
rect 137370 173884 137376 173896
rect 137428 173884 137434 173936
rect 155494 173884 155500 173936
rect 155552 173924 155558 173936
rect 155552 173896 159496 173924
rect 155552 173884 155558 173896
rect 124858 173816 124864 173868
rect 124916 173856 124922 173868
rect 128262 173856 128268 173868
rect 124916 173828 128268 173856
rect 124916 173816 124922 173828
rect 128262 173816 128268 173828
rect 128320 173816 128326 173868
rect 126974 173204 126980 173256
rect 127032 173244 127038 173256
rect 136542 173244 136548 173256
rect 127032 173216 136548 173244
rect 127032 173204 127038 173216
rect 136542 173204 136548 173216
rect 136600 173204 136606 173256
rect 135162 173136 135168 173188
rect 135220 173176 135226 173188
rect 135220 173148 138014 173176
rect 135220 173136 135226 173148
rect 62114 173000 62120 173052
rect 62172 173040 62178 173052
rect 65242 173040 65248 173052
rect 62172 173012 65248 173040
rect 62172 173000 62178 173012
rect 65242 173000 65248 173012
rect 65300 173000 65306 173052
rect 137986 172972 138014 173148
rect 159468 173052 159496 173896
rect 159450 173000 159456 173052
rect 159508 173000 159514 173052
rect 162854 172972 162860 172984
rect 137986 172944 162860 172972
rect 162854 172932 162860 172944
rect 162912 172932 162918 172984
rect 143442 172864 143448 172916
rect 143500 172904 143506 172916
rect 145650 172904 145656 172916
rect 143500 172876 145656 172904
rect 143500 172864 143506 172876
rect 145650 172864 145656 172876
rect 145708 172864 145714 172916
rect 146478 172864 146484 172916
rect 146536 172904 146542 172916
rect 148594 172904 148600 172916
rect 146536 172876 148600 172904
rect 146536 172864 146542 172876
rect 148594 172864 148600 172876
rect 148652 172864 148658 172916
rect 156506 172864 156512 172916
rect 156564 172904 156570 172916
rect 158438 172904 158444 172916
rect 156564 172876 158444 172904
rect 156564 172864 156570 172876
rect 158438 172864 158444 172876
rect 158496 172864 158502 172916
rect 143534 172796 143540 172848
rect 143592 172836 143598 172848
rect 146662 172836 146668 172848
rect 143592 172808 146668 172836
rect 143592 172796 143598 172808
rect 146662 172796 146668 172808
rect 146720 172796 146726 172848
rect 142430 172728 142436 172780
rect 142488 172768 142494 172780
rect 147582 172768 147588 172780
rect 142488 172740 147588 172768
rect 142488 172728 142494 172740
rect 147582 172728 147588 172740
rect 147640 172728 147646 172780
rect 45554 172456 45560 172508
rect 45612 172496 45618 172508
rect 46934 172496 46940 172508
rect 45612 172468 46940 172496
rect 45612 172456 45618 172468
rect 46934 172456 46940 172468
rect 46992 172456 46998 172508
rect 133874 172116 133880 172168
rect 133932 172156 133938 172168
rect 140774 172156 140780 172168
rect 133932 172128 140780 172156
rect 133932 172116 133938 172128
rect 140774 172116 140780 172128
rect 140832 172116 140838 172168
rect 131114 171844 131120 171896
rect 131172 171884 131178 171896
rect 138658 171884 138664 171896
rect 131172 171856 138664 171884
rect 131172 171844 131178 171856
rect 138658 171844 138664 171856
rect 138716 171844 138722 171896
rect 132494 171504 132500 171556
rect 132552 171544 132558 171556
rect 139670 171544 139676 171556
rect 132552 171516 139676 171544
rect 132552 171504 132558 171516
rect 139670 171504 139676 171516
rect 139728 171504 139734 171556
rect 128354 171096 128360 171148
rect 128412 171136 128418 171148
rect 136726 171136 136732 171148
rect 128412 171108 136732 171136
rect 128412 171096 128418 171108
rect 136726 171096 136732 171108
rect 136784 171096 136790 171148
rect 140774 171096 140780 171148
rect 140832 171136 140838 171148
rect 144914 171136 144920 171148
rect 140832 171108 144920 171136
rect 140832 171096 140838 171108
rect 144914 171096 144920 171108
rect 144972 171096 144978 171148
rect 84930 170076 84936 170128
rect 84988 170116 84994 170128
rect 88242 170116 88248 170128
rect 84988 170088 88248 170116
rect 84988 170076 84994 170088
rect 88242 170076 88248 170088
rect 88300 170076 88306 170128
rect 162854 169668 162860 169720
rect 162912 169708 162918 169720
rect 164970 169708 164976 169720
rect 162912 169680 164976 169708
rect 162912 169668 162918 169680
rect 164970 169668 164976 169680
rect 165028 169668 165034 169720
rect 46934 168988 46940 169040
rect 46992 169028 46998 169040
rect 50982 169028 50988 169040
rect 46992 169000 50988 169028
rect 46992 168988 46998 169000
rect 50982 168988 50988 169000
rect 51040 168988 51046 169040
rect 362218 168512 362224 168564
rect 362276 168552 362282 168564
rect 366358 168552 366364 168564
rect 362276 168524 366364 168552
rect 362276 168512 362282 168524
rect 366358 168512 366364 168524
rect 366416 168512 366422 168564
rect 84838 167628 84844 167680
rect 84896 167668 84902 167680
rect 87690 167668 87696 167680
rect 84896 167640 87696 167668
rect 84896 167628 84902 167640
rect 87690 167628 87696 167640
rect 87748 167628 87754 167680
rect 88242 167016 88248 167068
rect 88300 167056 88306 167068
rect 88300 167028 89760 167056
rect 88300 167016 88306 167028
rect 89732 166988 89760 167028
rect 91094 166988 91100 167000
rect 89732 166960 91100 166988
rect 91094 166948 91100 166960
rect 91152 166948 91158 167000
rect 164970 166268 164976 166320
rect 165028 166308 165034 166320
rect 167638 166308 167644 166320
rect 165028 166280 167644 166308
rect 165028 166268 165034 166280
rect 167638 166268 167644 166280
rect 167696 166268 167702 166320
rect 359366 166268 359372 166320
rect 359424 166308 359430 166320
rect 364978 166308 364984 166320
rect 359424 166280 364984 166308
rect 359424 166268 359430 166280
rect 364978 166268 364984 166280
rect 365036 166268 365042 166320
rect 185578 165588 185584 165640
rect 185636 165628 185642 165640
rect 579798 165628 579804 165640
rect 185636 165600 579804 165628
rect 185636 165588 185642 165600
rect 579798 165588 579804 165600
rect 579856 165588 579862 165640
rect 65242 165520 65248 165572
rect 65300 165560 65306 165572
rect 68278 165560 68284 165572
rect 65300 165532 68284 165560
rect 65300 165520 65306 165532
rect 68278 165520 68284 165532
rect 68336 165520 68342 165572
rect 86218 165520 86224 165572
rect 86276 165560 86282 165572
rect 88978 165560 88984 165572
rect 86276 165532 88984 165560
rect 86276 165520 86282 165532
rect 88978 165520 88984 165532
rect 89036 165520 89042 165572
rect 65518 165452 65524 165504
rect 65576 165492 65582 165504
rect 73798 165492 73804 165504
rect 65576 165464 73804 165492
rect 65576 165452 65582 165464
rect 73798 165452 73804 165464
rect 73856 165452 73862 165504
rect 128262 164840 128268 164892
rect 128320 164880 128326 164892
rect 137278 164880 137284 164892
rect 128320 164852 137284 164880
rect 128320 164840 128326 164852
rect 137278 164840 137284 164852
rect 137336 164840 137342 164892
rect 87690 164160 87696 164212
rect 87748 164200 87754 164212
rect 90358 164200 90364 164212
rect 87748 164172 90364 164200
rect 87748 164160 87754 164172
rect 90358 164160 90364 164172
rect 90416 164160 90422 164212
rect 91094 164160 91100 164212
rect 91152 164200 91158 164212
rect 93118 164200 93124 164212
rect 91152 164172 93124 164200
rect 91152 164160 91158 164172
rect 93118 164160 93124 164172
rect 93176 164160 93182 164212
rect 314654 163480 314660 163532
rect 314712 163520 314718 163532
rect 329098 163520 329104 163532
rect 314712 163492 329104 163520
rect 314712 163480 314718 163492
rect 329098 163480 329104 163492
rect 329156 163480 329162 163532
rect 3142 162868 3148 162920
rect 3200 162908 3206 162920
rect 175366 162908 175372 162920
rect 3200 162880 175372 162908
rect 3200 162868 3206 162880
rect 175366 162868 175372 162880
rect 175424 162868 175430 162920
rect 50982 162120 50988 162172
rect 51040 162160 51046 162172
rect 60550 162160 60556 162172
rect 51040 162132 60556 162160
rect 51040 162120 51046 162132
rect 60550 162120 60556 162132
rect 60608 162120 60614 162172
rect 338758 162120 338764 162172
rect 338816 162160 338822 162172
rect 359366 162160 359372 162172
rect 338816 162132 359372 162160
rect 338816 162120 338822 162132
rect 359366 162120 359372 162132
rect 359424 162120 359430 162172
rect 167638 160080 167644 160132
rect 167696 160120 167702 160132
rect 169018 160120 169024 160132
rect 167696 160092 169024 160120
rect 167696 160080 167702 160092
rect 169018 160080 169024 160092
rect 169076 160080 169082 160132
rect 360194 160080 360200 160132
rect 360252 160120 360258 160132
rect 362218 160120 362224 160132
rect 360252 160092 362224 160120
rect 360252 160080 360258 160092
rect 362218 160080 362224 160092
rect 362276 160080 362282 160132
rect 147490 159264 147496 159316
rect 147548 159304 147554 159316
rect 149698 159304 149704 159316
rect 147548 159276 149704 159304
rect 147548 159264 147554 159276
rect 149698 159264 149704 159276
rect 149756 159264 149762 159316
rect 60550 158992 60556 159044
rect 60608 159032 60614 159044
rect 66990 159032 66996 159044
rect 60608 159004 66996 159032
rect 60608 158992 60614 159004
rect 66990 158992 66996 159004
rect 67048 158992 67054 159044
rect 73798 158652 73804 158704
rect 73856 158692 73862 158704
rect 76742 158692 76748 158704
rect 73856 158664 76748 158692
rect 73856 158652 73862 158664
rect 76742 158652 76748 158664
rect 76800 158652 76806 158704
rect 309778 156544 309784 156596
rect 309836 156584 309842 156596
rect 314654 156584 314660 156596
rect 309836 156556 314660 156584
rect 309836 156544 309842 156556
rect 314654 156544 314660 156556
rect 314712 156544 314718 156596
rect 76742 155932 76748 155984
rect 76800 155972 76806 155984
rect 359458 155972 359464 155984
rect 76800 155944 81480 155972
rect 76800 155932 76806 155944
rect 81452 155904 81480 155944
rect 357452 155944 359464 155972
rect 84838 155904 84844 155916
rect 81452 155876 84844 155904
rect 84838 155864 84844 155876
rect 84896 155864 84902 155916
rect 129826 155864 129832 155916
rect 129884 155904 129890 155916
rect 134518 155904 134524 155916
rect 129884 155876 134524 155904
rect 129884 155864 129890 155876
rect 134518 155864 134524 155876
rect 134576 155864 134582 155916
rect 356698 155864 356704 155916
rect 356756 155904 356762 155916
rect 357452 155904 357480 155944
rect 359458 155932 359464 155944
rect 359516 155932 359522 155984
rect 356756 155876 357480 155904
rect 356756 155864 356762 155876
rect 137278 154504 137284 154556
rect 137336 154544 137342 154556
rect 140682 154544 140688 154556
rect 137336 154516 140688 154544
rect 137336 154504 137342 154516
rect 140682 154504 140688 154516
rect 140740 154504 140746 154556
rect 357986 154164 357992 154216
rect 358044 154204 358050 154216
rect 360194 154204 360200 154216
rect 358044 154176 360200 154204
rect 358044 154164 358050 154176
rect 360194 154164 360200 154176
rect 360252 154164 360258 154216
rect 84838 153212 84844 153264
rect 84896 153252 84902 153264
rect 129826 153252 129832 153264
rect 84896 153224 85620 153252
rect 84896 153212 84902 153224
rect 66990 153144 66996 153196
rect 67048 153184 67054 153196
rect 71038 153184 71044 153196
rect 67048 153156 71044 153184
rect 67048 153144 67054 153156
rect 71038 153144 71044 153156
rect 71096 153144 71102 153196
rect 85592 153184 85620 153224
rect 128372 153224 129832 153252
rect 87598 153184 87604 153196
rect 85592 153156 87604 153184
rect 87598 153144 87604 153156
rect 87656 153144 87662 153196
rect 127618 153144 127624 153196
rect 127676 153184 127682 153196
rect 128372 153184 128400 153224
rect 129826 153212 129832 153224
rect 129884 153212 129890 153264
rect 127676 153156 128400 153184
rect 127676 153144 127682 153156
rect 93118 151784 93124 151836
rect 93176 151824 93182 151836
rect 93176 151796 93900 151824
rect 93176 151784 93182 151796
rect 93872 151756 93900 151796
rect 95234 151756 95240 151768
rect 93872 151728 95240 151756
rect 95234 151716 95240 151728
rect 95292 151716 95298 151768
rect 88978 151512 88984 151564
rect 89036 151552 89042 151564
rect 90450 151552 90456 151564
rect 89036 151524 90456 151552
rect 89036 151512 89042 151524
rect 90450 151512 90456 151524
rect 90508 151512 90514 151564
rect 77938 151036 77944 151088
rect 77996 151076 78002 151088
rect 81434 151076 81440 151088
rect 77996 151048 81440 151076
rect 77996 151036 78002 151048
rect 81434 151036 81440 151048
rect 81492 151036 81498 151088
rect 169018 149676 169024 149728
rect 169076 149716 169082 149728
rect 170122 149716 170128 149728
rect 169076 149688 170128 149716
rect 169076 149676 169082 149688
rect 170122 149676 170128 149688
rect 170180 149676 170186 149728
rect 3142 149064 3148 149116
rect 3200 149104 3206 149116
rect 25498 149104 25504 149116
rect 3200 149076 25504 149104
rect 3200 149064 3206 149076
rect 25498 149064 25504 149076
rect 25556 149064 25562 149116
rect 307662 149064 307668 149116
rect 307720 149104 307726 149116
rect 309778 149104 309784 149116
rect 307720 149076 309784 149104
rect 307720 149064 307726 149076
rect 309778 149064 309784 149076
rect 309836 149064 309842 149116
rect 140682 148316 140688 148368
rect 140740 148356 140746 148368
rect 162118 148356 162124 148368
rect 140740 148328 162124 148356
rect 140740 148316 140746 148328
rect 162118 148316 162124 148328
rect 162176 148316 162182 148368
rect 170122 147568 170128 147620
rect 170180 147608 170186 147620
rect 172422 147608 172428 147620
rect 170180 147580 172428 147608
rect 170180 147568 170186 147580
rect 172422 147568 172428 147580
rect 172480 147568 172486 147620
rect 68278 146208 68284 146260
rect 68336 146248 68342 146260
rect 69658 146248 69664 146260
rect 68336 146220 69664 146248
rect 68336 146208 68342 146220
rect 69658 146208 69664 146220
rect 69716 146208 69722 146260
rect 95234 146208 95240 146260
rect 95292 146248 95298 146260
rect 97258 146248 97264 146260
rect 95292 146220 97264 146248
rect 95292 146208 95298 146220
rect 97258 146208 97264 146220
rect 97316 146208 97322 146260
rect 149698 146208 149704 146260
rect 149756 146248 149762 146260
rect 152642 146248 152648 146260
rect 149756 146220 152648 146248
rect 149756 146208 149762 146220
rect 152642 146208 152648 146220
rect 152700 146208 152706 146260
rect 81434 145528 81440 145580
rect 81492 145568 81498 145580
rect 91738 145568 91744 145580
rect 81492 145540 91744 145568
rect 81492 145528 81498 145540
rect 91738 145528 91744 145540
rect 91796 145528 91802 145580
rect 351914 145528 351920 145580
rect 351972 145568 351978 145580
rect 357986 145568 357992 145580
rect 351972 145540 357992 145568
rect 351972 145528 351978 145540
rect 357986 145528 357992 145540
rect 358044 145528 358050 145580
rect 303614 143556 303620 143608
rect 303672 143596 303678 143608
rect 307662 143596 307668 143608
rect 303672 143568 307668 143596
rect 303672 143556 303678 143568
rect 307662 143556 307668 143568
rect 307720 143556 307726 143608
rect 351914 143596 351920 143608
rect 347792 143568 351920 143596
rect 69658 143488 69664 143540
rect 69716 143528 69722 143540
rect 71130 143528 71136 143540
rect 69716 143500 71136 143528
rect 69716 143488 69722 143500
rect 71130 143488 71136 143500
rect 71188 143488 71194 143540
rect 75178 143488 75184 143540
rect 75236 143528 75242 143540
rect 76558 143528 76564 143540
rect 75236 143500 76564 143528
rect 75236 143488 75242 143500
rect 76558 143488 76564 143500
rect 76616 143488 76622 143540
rect 152642 143488 152648 143540
rect 152700 143528 152706 143540
rect 154850 143528 154856 143540
rect 152700 143500 154856 143528
rect 152700 143488 152706 143500
rect 154850 143488 154856 143500
rect 154908 143488 154914 143540
rect 347038 143488 347044 143540
rect 347096 143528 347102 143540
rect 347792 143528 347820 143568
rect 351914 143556 351920 143568
rect 351972 143556 351978 143608
rect 347096 143500 347820 143528
rect 347096 143488 347102 143500
rect 71038 143012 71044 143064
rect 71096 143052 71102 143064
rect 76650 143052 76656 143064
rect 71096 143024 76656 143052
rect 71096 143012 71102 143024
rect 76650 143012 76656 143024
rect 76708 143012 76714 143064
rect 115658 142808 115664 142860
rect 115716 142848 115722 142860
rect 580534 142848 580540 142860
rect 115716 142820 580540 142848
rect 115716 142808 115722 142820
rect 580534 142808 580540 142820
rect 580592 142808 580598 142860
rect 91738 141516 91744 141568
rect 91796 141556 91802 141568
rect 94038 141556 94044 141568
rect 91796 141528 94044 141556
rect 91796 141516 91802 141528
rect 94038 141516 94044 141528
rect 94096 141516 94102 141568
rect 66898 141244 66904 141296
rect 66956 141284 66962 141296
rect 68370 141284 68376 141296
rect 66956 141256 68376 141284
rect 66956 141244 66962 141256
rect 68370 141244 68376 141256
rect 68428 141244 68434 141296
rect 172514 138388 172520 138440
rect 172572 138428 172578 138440
rect 174354 138428 174360 138440
rect 172572 138400 174360 138428
rect 172572 138388 172578 138400
rect 174354 138388 174360 138400
rect 174412 138388 174418 138440
rect 3418 138320 3424 138372
rect 3476 138360 3482 138372
rect 4062 138360 4068 138372
rect 3476 138332 4068 138360
rect 3476 138320 3482 138332
rect 4062 138320 4068 138332
rect 4120 138320 4126 138372
rect 300854 138048 300860 138100
rect 300912 138088 300918 138100
rect 303614 138088 303620 138100
rect 300912 138060 303620 138088
rect 300912 138048 300918 138060
rect 303614 138048 303620 138060
rect 303672 138048 303678 138100
rect 90358 137980 90364 138032
rect 90416 138020 90422 138032
rect 93118 138020 93124 138032
rect 90416 137992 93124 138020
rect 90416 137980 90422 137992
rect 93118 137980 93124 137992
rect 93176 137980 93182 138032
rect 114370 137980 114376 138032
rect 114428 138020 114434 138032
rect 579982 138020 579988 138032
rect 114428 137992 579988 138020
rect 114428 137980 114434 137992
rect 579982 137980 579988 137992
rect 580040 137980 580046 138032
rect 90450 137912 90456 137964
rect 90508 137952 90514 137964
rect 94682 137952 94688 137964
rect 90508 137924 94688 137952
rect 90508 137912 90514 137924
rect 94682 137912 94688 137924
rect 94740 137912 94746 137964
rect 119338 137912 119344 137964
rect 119396 137952 119402 137964
rect 120718 137952 120724 137964
rect 119396 137924 120724 137952
rect 119396 137912 119402 137924
rect 120718 137912 120724 137924
rect 120776 137912 120782 137964
rect 142430 137912 142436 137964
rect 142488 137952 142494 137964
rect 145926 137952 145932 137964
rect 142488 137924 145932 137952
rect 142488 137912 142494 137924
rect 145926 137912 145932 137924
rect 145984 137912 145990 137964
rect 150526 137912 150532 137964
rect 150584 137952 150590 137964
rect 152182 137952 152188 137964
rect 150584 137924 152188 137952
rect 150584 137912 150590 137924
rect 152182 137912 152188 137924
rect 152240 137912 152246 137964
rect 164510 137912 164516 137964
rect 164568 137952 164574 137964
rect 172514 137952 172520 137964
rect 164568 137924 172520 137952
rect 164568 137912 164574 137924
rect 172514 137912 172520 137924
rect 172572 137912 172578 137964
rect 68370 137844 68376 137896
rect 68428 137884 68434 137896
rect 69658 137884 69664 137896
rect 68428 137856 69664 137884
rect 68428 137844 68434 137856
rect 69658 137844 69664 137856
rect 69716 137844 69722 137896
rect 154850 137708 154856 137760
rect 154908 137748 154914 137760
rect 164694 137748 164700 137760
rect 154908 137720 164700 137748
rect 154908 137708 154914 137720
rect 164694 137708 164700 137720
rect 164752 137708 164758 137760
rect 144454 137640 144460 137692
rect 144512 137680 144518 137692
rect 156874 137680 156880 137692
rect 144512 137652 156880 137680
rect 144512 137640 144518 137652
rect 156874 137640 156880 137652
rect 156932 137640 156938 137692
rect 163498 137640 163504 137692
rect 163556 137680 163562 137692
rect 174078 137680 174084 137692
rect 163556 137652 174084 137680
rect 163556 137640 163562 137652
rect 174078 137640 174084 137652
rect 174136 137640 174142 137692
rect 114094 137572 114100 137624
rect 114152 137612 114158 137624
rect 396902 137612 396908 137624
rect 114152 137584 396908 137612
rect 114152 137572 114158 137584
rect 396902 137572 396908 137584
rect 396960 137572 396966 137624
rect 114186 137504 114192 137556
rect 114244 137544 114250 137556
rect 397086 137544 397092 137556
rect 114244 137516 397092 137544
rect 114244 137504 114250 137516
rect 397086 137504 397092 137516
rect 397144 137504 397150 137556
rect 114278 137436 114284 137488
rect 114336 137476 114342 137488
rect 397178 137476 397184 137488
rect 114336 137448 397184 137476
rect 114336 137436 114342 137448
rect 397178 137436 397184 137448
rect 397236 137436 397242 137488
rect 113818 137368 113824 137420
rect 113876 137408 113882 137420
rect 412634 137408 412640 137420
rect 113876 137380 412640 137408
rect 113876 137368 113882 137380
rect 412634 137368 412640 137380
rect 412692 137368 412698 137420
rect 115106 137300 115112 137352
rect 115164 137340 115170 137352
rect 477494 137340 477500 137352
rect 115164 137312 477500 137340
rect 115164 137300 115170 137312
rect 477494 137300 477500 137312
rect 477552 137300 477558 137352
rect 115382 137232 115388 137284
rect 115440 137272 115446 137284
rect 580626 137272 580632 137284
rect 115440 137244 580632 137272
rect 115440 137232 115446 137244
rect 580626 137232 580632 137244
rect 580684 137232 580690 137284
rect 152458 137164 152464 137216
rect 152516 137204 152522 137216
rect 153746 137204 153752 137216
rect 152516 137176 153752 137204
rect 152516 137164 152522 137176
rect 153746 137164 153752 137176
rect 153804 137164 153810 137216
rect 163590 136756 163596 136808
rect 163648 136796 163654 136808
rect 170950 136796 170956 136808
rect 163648 136768 170956 136796
rect 163648 136756 163654 136768
rect 170950 136756 170956 136768
rect 171008 136756 171014 136808
rect 138106 136688 138112 136740
rect 138164 136728 138170 136740
rect 142522 136728 142528 136740
rect 138164 136700 142528 136728
rect 138164 136688 138170 136700
rect 142522 136688 142528 136700
rect 142580 136688 142586 136740
rect 153470 136688 153476 136740
rect 153528 136728 153534 136740
rect 155310 136728 155316 136740
rect 153528 136700 155316 136728
rect 153528 136688 153534 136700
rect 155310 136688 155316 136700
rect 155368 136688 155374 136740
rect 3418 136620 3424 136672
rect 3476 136660 3482 136672
rect 115198 136660 115204 136672
rect 3476 136632 115204 136660
rect 3476 136620 3482 136632
rect 115198 136620 115204 136632
rect 115256 136620 115262 136672
rect 174354 136552 174360 136604
rect 174412 136592 174418 136604
rect 176010 136592 176016 136604
rect 174412 136564 176016 136592
rect 174412 136552 174418 136564
rect 176010 136552 176016 136564
rect 176068 136552 176074 136604
rect 162118 136484 162124 136536
rect 162176 136524 162182 136536
rect 175918 136524 175924 136536
rect 162176 136496 175924 136524
rect 162176 136484 162182 136496
rect 175918 136484 175924 136496
rect 175976 136484 175982 136536
rect 40034 136416 40040 136468
rect 40092 136456 40098 136468
rect 176838 136456 176844 136468
rect 40092 136428 176844 136456
rect 40092 136416 40098 136428
rect 176838 136416 176844 136428
rect 176896 136416 176902 136468
rect 3970 136348 3976 136400
rect 4028 136388 4034 136400
rect 178126 136388 178132 136400
rect 4028 136360 178132 136388
rect 4028 136348 4034 136360
rect 178126 136348 178132 136360
rect 178184 136348 178190 136400
rect 3786 136280 3792 136332
rect 3844 136320 3850 136332
rect 178586 136320 178592 136332
rect 3844 136292 178592 136320
rect 3844 136280 3850 136292
rect 178586 136280 178592 136292
rect 178644 136280 178650 136332
rect 3878 136212 3884 136264
rect 3936 136252 3942 136264
rect 178402 136252 178408 136264
rect 3936 136224 178408 136252
rect 3936 136212 3942 136224
rect 178402 136212 178408 136224
rect 178460 136212 178466 136264
rect 3694 136144 3700 136196
rect 3752 136184 3758 136196
rect 178770 136184 178776 136196
rect 3752 136156 178776 136184
rect 3752 136144 3758 136156
rect 178770 136144 178776 136156
rect 178828 136144 178834 136196
rect 3234 136076 3240 136128
rect 3292 136116 3298 136128
rect 178034 136116 178040 136128
rect 3292 136088 178040 136116
rect 3292 136076 3298 136088
rect 178034 136076 178040 136088
rect 178092 136076 178098 136128
rect 3326 136008 3332 136060
rect 3384 136048 3390 136060
rect 178494 136048 178500 136060
rect 3384 136020 178500 136048
rect 3384 136008 3390 136020
rect 178494 136008 178500 136020
rect 178552 136008 178558 136060
rect 295334 136008 295340 136060
rect 295392 136048 295398 136060
rect 300854 136048 300860 136060
rect 295392 136020 300860 136048
rect 295392 136008 295398 136020
rect 300854 136008 300860 136020
rect 300912 136008 300918 136060
rect 115474 135940 115480 135992
rect 115532 135980 115538 135992
rect 580810 135980 580816 135992
rect 115532 135952 580816 135980
rect 115532 135940 115538 135952
rect 580810 135940 580816 135952
rect 580868 135940 580874 135992
rect 94038 135872 94044 135924
rect 94096 135912 94102 135924
rect 105538 135912 105544 135924
rect 94096 135884 105544 135912
rect 94096 135872 94102 135884
rect 105538 135872 105544 135884
rect 105596 135872 105602 135924
rect 113910 135872 113916 135924
rect 113968 135912 113974 135924
rect 580074 135912 580080 135924
rect 113968 135884 580080 135912
rect 113968 135872 113974 135884
rect 580074 135872 580080 135884
rect 580132 135872 580138 135924
rect 71130 135192 71136 135244
rect 71188 135232 71194 135244
rect 72418 135232 72424 135244
rect 71188 135204 72424 135232
rect 71188 135192 71194 135204
rect 72418 135192 72424 135204
rect 72476 135192 72482 135244
rect 115566 134784 115572 134836
rect 115624 134824 115630 134836
rect 127618 134824 127624 134836
rect 115624 134796 127624 134824
rect 115624 134784 115630 134796
rect 127618 134784 127624 134796
rect 127676 134784 127682 134836
rect 87598 134716 87604 134768
rect 87656 134756 87662 134768
rect 177298 134756 177304 134768
rect 87656 134728 177304 134756
rect 87656 134716 87662 134728
rect 177298 134716 177304 134728
rect 177356 134716 177362 134768
rect 3602 134648 3608 134700
rect 3660 134688 3666 134700
rect 178310 134688 178316 134700
rect 3660 134660 178316 134688
rect 3660 134648 3666 134660
rect 178310 134648 178316 134660
rect 178368 134648 178374 134700
rect 4062 134580 4068 134632
rect 4120 134620 4126 134632
rect 178678 134620 178684 134632
rect 4120 134592 178684 134620
rect 4120 134580 4126 134592
rect 178678 134580 178684 134592
rect 178736 134580 178742 134632
rect 113726 134512 113732 134564
rect 113784 134552 113790 134564
rect 295334 134552 295340 134564
rect 113784 134524 295340 134552
rect 113784 134512 113790 134524
rect 295334 134512 295340 134524
rect 295392 134512 295398 134564
rect 3786 133900 3792 133952
rect 3844 133940 3850 133952
rect 175366 133940 175372 133952
rect 3844 133912 175372 133940
rect 3844 133900 3850 133912
rect 175366 133900 175372 133912
rect 175424 133900 175430 133952
rect 94682 133832 94688 133884
rect 94740 133872 94746 133884
rect 95602 133872 95608 133884
rect 94740 133844 95608 133872
rect 94740 133832 94746 133844
rect 95602 133832 95608 133844
rect 95660 133832 95666 133884
rect 76650 133152 76656 133204
rect 76708 133192 76714 133204
rect 86218 133192 86224 133204
rect 76708 133164 86224 133192
rect 76708 133152 76714 133164
rect 86218 133152 86224 133164
rect 86276 133152 86282 133204
rect 115106 132676 115112 132728
rect 115164 132716 115170 132728
rect 115290 132716 115296 132728
rect 115164 132688 115296 132716
rect 115164 132676 115170 132688
rect 115290 132676 115296 132688
rect 115348 132676 115354 132728
rect 95602 131724 95608 131776
rect 95660 131764 95666 131776
rect 97534 131764 97540 131776
rect 95660 131736 97540 131764
rect 95660 131724 95666 131736
rect 97534 131724 97540 131736
rect 97592 131724 97598 131776
rect 97258 131588 97264 131640
rect 97316 131628 97322 131640
rect 99282 131628 99288 131640
rect 97316 131600 99288 131628
rect 97316 131588 97322 131600
rect 99282 131588 99288 131600
rect 99340 131588 99346 131640
rect 3418 131112 3424 131164
rect 3476 131152 3482 131164
rect 113634 131152 113640 131164
rect 3476 131124 113640 131152
rect 3476 131112 3482 131124
rect 113634 131112 113640 131124
rect 113692 131112 113698 131164
rect 3602 128324 3608 128376
rect 3660 128364 3666 128376
rect 113542 128364 113548 128376
rect 3660 128336 113548 128364
rect 3660 128324 3666 128336
rect 113542 128324 113548 128336
rect 113600 128324 113606 128376
rect 93118 128256 93124 128308
rect 93176 128296 93182 128308
rect 95878 128296 95884 128308
rect 93176 128268 95884 128296
rect 93176 128256 93182 128268
rect 95878 128256 95884 128268
rect 95936 128256 95942 128308
rect 76558 127576 76564 127628
rect 76616 127616 76622 127628
rect 79318 127616 79324 127628
rect 76616 127588 79324 127616
rect 76616 127576 76622 127588
rect 79318 127576 79324 127588
rect 79376 127576 79382 127628
rect 105538 127576 105544 127628
rect 105596 127616 105602 127628
rect 111058 127616 111064 127628
rect 105596 127588 111064 127616
rect 105596 127576 105602 127588
rect 111058 127576 111064 127588
rect 111116 127576 111122 127628
rect 3694 126964 3700 127016
rect 3752 127004 3758 127016
rect 113542 127004 113548 127016
rect 3752 126976 113548 127004
rect 3752 126964 3758 126976
rect 113542 126964 113548 126976
rect 113600 126964 113606 127016
rect 25498 126896 25504 126948
rect 25556 126936 25562 126948
rect 113634 126936 113640 126948
rect 25556 126908 113640 126936
rect 25556 126896 25562 126908
rect 113634 126896 113640 126908
rect 113692 126896 113698 126948
rect 99374 126828 99380 126880
rect 99432 126868 99438 126880
rect 101490 126868 101496 126880
rect 99432 126840 101496 126868
rect 99432 126828 99438 126840
rect 101490 126828 101496 126840
rect 101548 126828 101554 126880
rect 184198 125604 184204 125656
rect 184256 125644 184262 125656
rect 580074 125644 580080 125656
rect 184256 125616 580080 125644
rect 184256 125604 184262 125616
rect 580074 125604 580080 125616
rect 580132 125604 580138 125656
rect 22830 125536 22836 125588
rect 22888 125576 22894 125588
rect 113634 125576 113640 125588
rect 22888 125548 113640 125576
rect 22888 125536 22894 125548
rect 113634 125536 113640 125548
rect 113692 125536 113698 125588
rect 350718 124176 350724 124228
rect 350776 124216 350782 124228
rect 356698 124216 356704 124228
rect 350776 124188 356704 124216
rect 350776 124176 350782 124188
rect 356698 124176 356704 124188
rect 356756 124176 356762 124228
rect 22738 124108 22744 124160
rect 22796 124148 22802 124160
rect 113634 124148 113640 124160
rect 22796 124120 113640 124148
rect 22796 124108 22802 124120
rect 113634 124108 113640 124120
rect 113692 124108 113698 124160
rect 97534 124040 97540 124092
rect 97592 124080 97598 124092
rect 99282 124080 99288 124092
rect 97592 124052 99288 124080
rect 97592 124040 97598 124052
rect 99282 124040 99288 124052
rect 99340 124040 99346 124092
rect 24118 122748 24124 122800
rect 24176 122788 24182 122800
rect 113634 122788 113640 122800
rect 24176 122760 113640 122788
rect 24176 122748 24182 122760
rect 113634 122748 113640 122760
rect 113692 122748 113698 122800
rect 72418 121456 72424 121508
rect 72476 121496 72482 121508
rect 73798 121496 73804 121508
rect 72476 121468 73804 121496
rect 72476 121456 72482 121468
rect 73798 121456 73804 121468
rect 73856 121456 73862 121508
rect 86218 121456 86224 121508
rect 86276 121496 86282 121508
rect 88978 121496 88984 121508
rect 86276 121468 88984 121496
rect 86276 121456 86282 121468
rect 88978 121456 88984 121468
rect 89036 121456 89042 121508
rect 345750 121456 345756 121508
rect 345808 121496 345814 121508
rect 347038 121496 347044 121508
rect 345808 121468 347044 121496
rect 345808 121456 345814 121468
rect 347038 121456 347044 121468
rect 347096 121456 347102 121508
rect 347866 121456 347872 121508
rect 347924 121496 347930 121508
rect 350718 121496 350724 121508
rect 347924 121468 350724 121496
rect 347924 121456 347930 121468
rect 350718 121456 350724 121468
rect 350776 121456 350782 121508
rect 10318 121388 10324 121440
rect 10376 121428 10382 121440
rect 113634 121428 113640 121440
rect 10376 121400 113640 121428
rect 10376 121388 10382 121400
rect 113634 121388 113640 121400
rect 113692 121388 113698 121440
rect 101490 121320 101496 121372
rect 101548 121360 101554 121372
rect 104894 121360 104900 121372
rect 101548 121332 104900 121360
rect 101548 121320 101554 121332
rect 104894 121320 104900 121332
rect 104952 121320 104958 121372
rect 99374 121252 99380 121304
rect 99432 121292 99438 121304
rect 102042 121292 102048 121304
rect 99432 121264 102048 121292
rect 99432 121252 99438 121264
rect 102042 121252 102048 121264
rect 102100 121252 102106 121304
rect 8938 120028 8944 120080
rect 8996 120068 9002 120080
rect 113634 120068 113640 120080
rect 8996 120040 113640 120068
rect 8996 120028 9002 120040
rect 113634 120028 113640 120040
rect 113692 120028 113698 120080
rect 69658 119960 69664 120012
rect 69716 120000 69722 120012
rect 70486 120000 70492 120012
rect 69716 119972 70492 120000
rect 69716 119960 69722 119972
rect 70486 119960 70492 119972
rect 70544 119960 70550 120012
rect 104894 119620 104900 119672
rect 104952 119660 104958 119672
rect 106918 119660 106924 119672
rect 104952 119632 106924 119660
rect 104952 119620 104958 119632
rect 106918 119620 106924 119632
rect 106976 119620 106982 119672
rect 5074 118600 5080 118652
rect 5132 118640 5138 118652
rect 113634 118640 113640 118652
rect 5132 118612 113640 118640
rect 5132 118600 5138 118612
rect 113634 118600 113640 118612
rect 113692 118600 113698 118652
rect 70486 118532 70492 118584
rect 70544 118572 70550 118584
rect 76282 118572 76288 118584
rect 70544 118544 76288 118572
rect 70544 118532 70550 118544
rect 76282 118532 76288 118544
rect 76340 118532 76346 118584
rect 177298 118532 177304 118584
rect 177356 118572 177362 118584
rect 178218 118572 178224 118584
rect 177356 118544 178224 118572
rect 177356 118532 177362 118544
rect 178218 118532 178224 118544
rect 178276 118532 178282 118584
rect 79318 118260 79324 118312
rect 79376 118300 79382 118312
rect 81158 118300 81164 118312
rect 79376 118272 81164 118300
rect 79376 118260 79382 118272
rect 81158 118260 81164 118272
rect 81216 118260 81222 118312
rect 342254 118192 342260 118244
rect 342312 118232 342318 118244
rect 345750 118232 345756 118244
rect 342312 118204 345756 118232
rect 342312 118192 342318 118204
rect 345750 118192 345756 118204
rect 345808 118192 345814 118244
rect 343634 117920 343640 117972
rect 343692 117960 343698 117972
rect 347866 117960 347872 117972
rect 343692 117932 347872 117960
rect 343692 117920 343698 117932
rect 347866 117920 347872 117932
rect 347924 117920 347930 117972
rect 33778 117240 33784 117292
rect 33836 117280 33842 117292
rect 113634 117280 113640 117292
rect 33836 117252 113640 117280
rect 33836 117240 33842 117252
rect 113634 117240 113640 117252
rect 113692 117240 113698 117292
rect 176010 117240 176016 117292
rect 176068 117280 176074 117292
rect 176654 117280 176660 117292
rect 176068 117252 176660 117280
rect 176068 117240 176074 117252
rect 176654 117240 176660 117252
rect 176712 117240 176718 117292
rect 76282 116016 76288 116068
rect 76340 116056 76346 116068
rect 77938 116056 77944 116068
rect 76340 116028 77944 116056
rect 76340 116016 76346 116028
rect 77938 116016 77944 116028
rect 77996 116016 78002 116068
rect 29638 115880 29644 115932
rect 29696 115920 29702 115932
rect 113542 115920 113548 115932
rect 29696 115892 113548 115920
rect 29696 115880 29702 115892
rect 113542 115880 113548 115892
rect 113600 115880 113606 115932
rect 342254 114560 342260 114572
rect 340892 114532 342260 114560
rect 81158 114452 81164 114504
rect 81216 114492 81222 114504
rect 82814 114492 82820 114504
rect 81216 114464 82820 114492
rect 81216 114452 81222 114464
rect 82814 114452 82820 114464
rect 82872 114452 82878 114504
rect 340414 114452 340420 114504
rect 340472 114492 340478 114504
rect 340892 114492 340920 114532
rect 342254 114520 342260 114532
rect 342312 114520 342318 114572
rect 340472 114464 340920 114492
rect 340472 114452 340478 114464
rect 341518 113704 341524 113756
rect 341576 113744 341582 113756
rect 343634 113744 343640 113756
rect 341576 113716 343640 113744
rect 341576 113704 341582 113716
rect 343634 113704 343640 113716
rect 343692 113704 343698 113756
rect 37918 113092 37924 113144
rect 37976 113132 37982 113144
rect 113634 113132 113640 113144
rect 37976 113104 113640 113132
rect 37976 113092 37982 113104
rect 113634 113092 113640 113104
rect 113692 113092 113698 113144
rect 95878 112412 95884 112464
rect 95936 112452 95942 112464
rect 108298 112452 108304 112464
rect 95936 112424 108304 112452
rect 95936 112412 95942 112424
rect 108298 112412 108304 112424
rect 108356 112412 108362 112464
rect 333974 112412 333980 112464
rect 334032 112452 334038 112464
rect 340414 112452 340420 112464
rect 334032 112424 340420 112452
rect 334032 112412 334038 112424
rect 340414 112412 340420 112424
rect 340472 112412 340478 112464
rect 77938 112276 77944 112328
rect 77996 112316 78002 112328
rect 79962 112316 79968 112328
rect 77996 112288 79968 112316
rect 77996 112276 78002 112288
rect 79962 112276 79968 112288
rect 80020 112276 80026 112328
rect 15838 111732 15844 111784
rect 15896 111772 15902 111784
rect 113634 111772 113640 111784
rect 15896 111744 113640 111772
rect 15896 111732 15902 111744
rect 113634 111732 113640 111744
rect 113692 111732 113698 111784
rect 82814 111052 82820 111104
rect 82872 111092 82878 111104
rect 88242 111092 88248 111104
rect 82872 111064 88248 111092
rect 82872 111052 82878 111064
rect 88242 111052 88248 111064
rect 88300 111052 88306 111104
rect 324314 111052 324320 111104
rect 324372 111092 324378 111104
rect 333974 111092 333980 111104
rect 324372 111064 333980 111092
rect 324372 111052 324378 111064
rect 333974 111052 333980 111064
rect 334032 111052 334038 111104
rect 23474 110372 23480 110424
rect 23532 110412 23538 110424
rect 113634 110412 113640 110424
rect 23532 110384 113640 110412
rect 23532 110372 23538 110384
rect 113634 110372 113640 110384
rect 113692 110372 113698 110424
rect 108298 108944 108304 108996
rect 108356 108984 108362 108996
rect 113634 108984 113640 108996
rect 108356 108956 113640 108984
rect 108356 108944 108362 108956
rect 113634 108944 113640 108956
rect 113692 108944 113698 108996
rect 80054 107584 80060 107636
rect 80112 107624 80118 107636
rect 113634 107624 113640 107636
rect 80112 107596 113640 107624
rect 80112 107584 80118 107596
rect 113634 107584 113640 107596
rect 113692 107584 113698 107636
rect 102134 107516 102140 107568
rect 102192 107556 102198 107568
rect 106182 107556 106188 107568
rect 102192 107528 106188 107556
rect 102192 107516 102198 107528
rect 106182 107516 106188 107528
rect 106240 107516 106246 107568
rect 106182 106224 106188 106276
rect 106240 106264 106246 106276
rect 113542 106264 113548 106276
rect 106240 106236 113548 106264
rect 106240 106224 106246 106236
rect 113542 106224 113548 106236
rect 113600 106224 113606 106276
rect 178034 106224 178040 106276
rect 178092 106264 178098 106276
rect 341518 106264 341524 106276
rect 178092 106236 341524 106264
rect 178092 106224 178098 106236
rect 341518 106224 341524 106236
rect 341576 106224 341582 106276
rect 88242 104864 88248 104916
rect 88300 104904 88306 104916
rect 88300 104876 93854 104904
rect 88300 104864 88306 104876
rect 93826 104836 93854 104876
rect 113634 104836 113640 104848
rect 93826 104808 113640 104836
rect 113634 104796 113640 104808
rect 113692 104796 113698 104848
rect 178034 104796 178040 104848
rect 178092 104836 178098 104848
rect 324222 104836 324228 104848
rect 178092 104808 324228 104836
rect 178092 104796 178098 104808
rect 324222 104796 324228 104808
rect 324280 104796 324286 104848
rect 106918 104728 106924 104780
rect 106976 104768 106982 104780
rect 108390 104768 108396 104780
rect 106976 104740 108396 104768
rect 106976 104728 106982 104740
rect 108390 104728 108396 104740
rect 108448 104728 108454 104780
rect 88978 103844 88984 103896
rect 89036 103884 89042 103896
rect 95234 103884 95240 103896
rect 89036 103856 95240 103884
rect 89036 103844 89042 103856
rect 95234 103844 95240 103856
rect 95292 103844 95298 103896
rect 178034 103436 178040 103488
rect 178092 103476 178098 103488
rect 410518 103476 410524 103488
rect 178092 103448 410524 103476
rect 178092 103436 178098 103448
rect 410518 103436 410524 103448
rect 410576 103436 410582 103488
rect 178034 102076 178040 102128
rect 178092 102116 178098 102128
rect 409138 102116 409144 102128
rect 178092 102088 409144 102116
rect 178092 102076 178098 102088
rect 409138 102076 409144 102088
rect 409196 102076 409202 102128
rect 178034 100648 178040 100700
rect 178092 100688 178098 100700
rect 407758 100688 407764 100700
rect 178092 100660 407764 100688
rect 178092 100648 178098 100660
rect 407758 100648 407764 100660
rect 407816 100648 407822 100700
rect 175918 99356 175924 99408
rect 175976 99396 175982 99408
rect 580074 99396 580080 99408
rect 175976 99368 580080 99396
rect 175976 99356 175982 99368
rect 580074 99356 580080 99368
rect 580132 99356 580138 99408
rect 178034 99288 178040 99340
rect 178092 99328 178098 99340
rect 566458 99328 566464 99340
rect 178092 99300 566464 99328
rect 178092 99288 178098 99300
rect 566458 99288 566464 99300
rect 566516 99288 566522 99340
rect 95234 98676 95240 98728
rect 95292 98716 95298 98728
rect 98638 98716 98644 98728
rect 95292 98688 98644 98716
rect 95292 98676 95298 98688
rect 98638 98676 98644 98688
rect 98696 98676 98702 98728
rect 73798 98608 73804 98660
rect 73856 98648 73862 98660
rect 77938 98648 77944 98660
rect 73856 98620 77944 98648
rect 73856 98608 73862 98620
rect 77938 98608 77944 98620
rect 77996 98608 78002 98660
rect 178034 97928 178040 97980
rect 178092 97968 178098 97980
rect 406378 97968 406384 97980
rect 178092 97940 406384 97968
rect 178092 97928 178098 97940
rect 406378 97928 406384 97940
rect 406436 97928 406442 97980
rect 108390 96636 108396 96688
rect 108448 96676 108454 96688
rect 108448 96648 109080 96676
rect 108448 96636 108454 96648
rect 109052 96608 109080 96648
rect 110966 96608 110972 96620
rect 109052 96580 110972 96608
rect 110966 96568 110972 96580
rect 111024 96568 111030 96620
rect 178034 95140 178040 95192
rect 178092 95180 178098 95192
rect 404998 95180 405004 95192
rect 178092 95152 405004 95180
rect 178092 95140 178098 95152
rect 404998 95140 405004 95152
rect 405056 95140 405062 95192
rect 178034 93780 178040 93832
rect 178092 93820 178098 93832
rect 403618 93820 403624 93832
rect 178092 93792 403624 93820
rect 178092 93780 178098 93792
rect 403618 93780 403624 93792
rect 403676 93780 403682 93832
rect 178034 92420 178040 92472
rect 178092 92460 178098 92472
rect 400858 92460 400864 92472
rect 178092 92432 400864 92460
rect 178092 92420 178098 92432
rect 400858 92420 400864 92432
rect 400916 92420 400922 92472
rect 320818 91740 320824 91792
rect 320876 91780 320882 91792
rect 338758 91780 338764 91792
rect 320876 91752 338764 91780
rect 320876 91740 320882 91752
rect 338758 91740 338764 91752
rect 338816 91740 338822 91792
rect 178034 90992 178040 91044
rect 178092 91032 178098 91044
rect 417418 91032 417424 91044
rect 178092 91004 417424 91032
rect 178092 90992 178098 91004
rect 417418 90992 417424 91004
rect 417476 90992 417482 91044
rect 178034 89632 178040 89684
rect 178092 89672 178098 89684
rect 414658 89672 414664 89684
rect 178092 89644 414664 89672
rect 178092 89632 178098 89644
rect 414658 89632 414664 89644
rect 414716 89632 414722 89684
rect 110966 88272 110972 88324
rect 111024 88312 111030 88324
rect 113818 88312 113824 88324
rect 111024 88284 113824 88312
rect 111024 88272 111030 88284
rect 113818 88272 113824 88284
rect 113876 88272 113882 88324
rect 178034 88272 178040 88324
rect 178092 88312 178098 88324
rect 552658 88312 552664 88324
rect 178092 88284 552664 88312
rect 178092 88272 178098 88284
rect 552658 88272 552664 88284
rect 552716 88272 552722 88324
rect 77938 86980 77944 87032
rect 77996 87020 78002 87032
rect 77996 86992 81480 87020
rect 77996 86980 78002 86992
rect 81452 86952 81480 86992
rect 83550 86952 83556 86964
rect 81452 86924 83556 86952
rect 83550 86912 83556 86924
rect 83608 86912 83614 86964
rect 178034 86912 178040 86964
rect 178092 86952 178098 86964
rect 413278 86952 413284 86964
rect 178092 86924 413284 86952
rect 178092 86912 178098 86924
rect 413278 86912 413284 86924
rect 413336 86912 413342 86964
rect 179230 85552 179236 85604
rect 179288 85592 179294 85604
rect 580074 85592 580080 85604
rect 179288 85564 580080 85592
rect 179288 85552 179294 85564
rect 580074 85552 580080 85564
rect 580132 85552 580138 85604
rect 178034 85484 178040 85536
rect 178092 85524 178098 85536
rect 188338 85524 188344 85536
rect 178092 85496 188344 85524
rect 178092 85484 178098 85496
rect 188338 85484 188344 85496
rect 188396 85484 188402 85536
rect 307754 84804 307760 84856
rect 307812 84844 307818 84856
rect 320818 84844 320824 84856
rect 307812 84816 320824 84844
rect 307812 84804 307818 84816
rect 320818 84804 320824 84816
rect 320876 84804 320882 84856
rect 3326 84192 3332 84244
rect 3384 84232 3390 84244
rect 116578 84232 116584 84244
rect 3384 84204 116584 84232
rect 3384 84192 3390 84204
rect 116578 84192 116584 84204
rect 116636 84192 116642 84244
rect 178034 84124 178040 84176
rect 178092 84164 178098 84176
rect 185578 84164 185584 84176
rect 178092 84136 185584 84164
rect 178092 84124 178098 84136
rect 185578 84124 185584 84136
rect 185636 84124 185642 84176
rect 98638 82832 98644 82884
rect 98696 82872 98702 82884
rect 104158 82872 104164 82884
rect 98696 82844 104164 82872
rect 98696 82832 98702 82844
rect 104158 82832 104164 82844
rect 104216 82832 104222 82884
rect 178034 82764 178040 82816
rect 178092 82804 178098 82816
rect 184198 82804 184204 82816
rect 178092 82776 184204 82804
rect 178092 82764 178098 82776
rect 184198 82764 184204 82776
rect 184256 82764 184262 82816
rect 113818 81608 113824 81660
rect 113876 81648 113882 81660
rect 114554 81648 114560 81660
rect 113876 81620 114560 81648
rect 113876 81608 113882 81620
rect 114554 81608 114560 81620
rect 114612 81608 114618 81660
rect 83550 79976 83556 80028
rect 83608 80016 83614 80028
rect 84838 80016 84844 80028
rect 83608 79988 84844 80016
rect 83608 79976 83614 79988
rect 84838 79976 84844 79988
rect 84896 79976 84902 80028
rect 299382 77936 299388 77988
rect 299440 77976 299446 77988
rect 307754 77976 307760 77988
rect 299440 77948 307760 77976
rect 299440 77936 299446 77948
rect 307754 77936 307760 77948
rect 307812 77936 307818 77988
rect 178034 75896 178040 75948
rect 178092 75936 178098 75948
rect 562318 75936 562324 75948
rect 178092 75908 562324 75936
rect 178092 75896 178098 75908
rect 562318 75896 562324 75908
rect 562376 75896 562382 75948
rect 114462 75692 114468 75744
rect 114520 75732 114526 75744
rect 175918 75732 175924 75744
rect 114520 75704 175924 75732
rect 114520 75692 114526 75704
rect 175918 75692 175924 75704
rect 175976 75692 175982 75744
rect 114554 75624 114560 75676
rect 114612 75664 114618 75676
rect 118602 75664 118608 75676
rect 114612 75636 118608 75664
rect 114612 75624 114618 75636
rect 118602 75624 118608 75636
rect 118660 75624 118666 75676
rect 170674 75664 170680 75676
rect 157306 75636 170680 75664
rect 157306 75460 157334 75636
rect 170674 75624 170680 75636
rect 170732 75624 170738 75676
rect 147646 75432 157334 75460
rect 159376 75568 164234 75596
rect 29730 75216 29736 75268
rect 29788 75256 29794 75268
rect 147646 75256 147674 75432
rect 159376 75392 159404 75568
rect 150406 75364 159404 75392
rect 164206 75392 164234 75568
rect 164206 75364 172376 75392
rect 150406 75324 150434 75364
rect 172238 75324 172244 75336
rect 29788 75228 147674 75256
rect 149716 75296 150434 75324
rect 164206 75296 172244 75324
rect 29788 75216 29794 75228
rect 149716 75120 149744 75296
rect 164206 75256 164234 75296
rect 172238 75284 172244 75296
rect 172296 75284 172302 75336
rect 170398 75256 170404 75268
rect 142126 75092 149744 75120
rect 150636 75228 164234 75256
rect 164528 75228 170404 75256
rect 141786 74876 141792 74928
rect 141844 74916 141850 74928
rect 142126 74916 142154 75092
rect 150636 74928 150664 75228
rect 164528 75188 164556 75228
rect 170398 75216 170404 75228
rect 170456 75216 170462 75268
rect 170490 75188 170496 75200
rect 162826 75160 164556 75188
rect 164988 75160 170496 75188
rect 141844 74888 142154 74916
rect 141844 74876 141850 74888
rect 150618 74876 150624 74928
rect 150676 74876 150682 74928
rect 162826 74916 162854 75160
rect 157306 74888 162854 74916
rect 145098 74808 145104 74860
rect 145156 74848 145162 74860
rect 157306 74848 157334 74888
rect 164418 74876 164424 74928
rect 164476 74916 164482 74928
rect 164988 74916 165016 75160
rect 170490 75148 170496 75160
rect 170548 75148 170554 75200
rect 170582 75120 170588 75132
rect 165080 75092 170588 75120
rect 165080 74928 165108 75092
rect 170582 75080 170588 75092
rect 170640 75080 170646 75132
rect 172348 75120 172376 75364
rect 175366 75148 175372 75200
rect 175424 75188 175430 75200
rect 299382 75188 299388 75200
rect 175424 75160 299388 75188
rect 175424 75148 175430 75160
rect 299382 75148 299388 75160
rect 299440 75148 299446 75200
rect 259454 75120 259460 75132
rect 172348 75092 259460 75120
rect 259454 75080 259460 75092
rect 259512 75080 259518 75132
rect 170858 75012 170864 75064
rect 170916 75052 170922 75064
rect 195974 75052 195980 75064
rect 170916 75024 195980 75052
rect 170916 75012 170922 75024
rect 195974 75012 195980 75024
rect 196032 75012 196038 75064
rect 170398 74944 170404 74996
rect 170456 74984 170462 74996
rect 302234 74984 302240 74996
rect 170456 74956 302240 74984
rect 170456 74944 170462 74956
rect 302234 74944 302240 74956
rect 302292 74944 302298 74996
rect 164476 74888 165016 74916
rect 164476 74876 164482 74888
rect 165062 74876 165068 74928
rect 165120 74876 165126 74928
rect 165356 74888 169616 74916
rect 145156 74820 157334 74848
rect 162826 74820 164234 74848
rect 145156 74808 145162 74820
rect 157306 74752 161474 74780
rect 146754 74672 146760 74724
rect 146812 74712 146818 74724
rect 157306 74712 157334 74752
rect 161446 74712 161474 74752
rect 162826 74712 162854 74820
rect 164206 74780 164234 74820
rect 165356 74780 165384 74888
rect 164206 74752 165384 74780
rect 168098 74740 168104 74792
rect 168156 74740 168162 74792
rect 146812 74684 157334 74712
rect 160388 74684 160600 74712
rect 161446 74684 162854 74712
rect 168116 74712 168144 74740
rect 168116 74684 169432 74712
rect 146812 74672 146818 74684
rect 153378 74400 153384 74452
rect 153436 74440 153442 74452
rect 160388 74440 160416 74684
rect 160572 74576 160600 74684
rect 169404 74656 169432 74684
rect 168098 74644 168104 74656
rect 164206 74616 168104 74644
rect 164206 74576 164234 74616
rect 168098 74604 168104 74616
rect 168156 74604 168162 74656
rect 169386 74604 169392 74656
rect 169444 74604 169450 74656
rect 169588 74644 169616 74888
rect 169754 74876 169760 74928
rect 169812 74916 169818 74928
rect 169812 74888 169984 74916
rect 169812 74876 169818 74888
rect 169956 74848 169984 74888
rect 170766 74876 170772 74928
rect 170824 74916 170830 74928
rect 324314 74916 324320 74928
rect 170824 74888 324320 74916
rect 170824 74876 170830 74888
rect 324314 74876 324320 74888
rect 324372 74876 324378 74928
rect 170674 74848 170680 74860
rect 169956 74820 170680 74848
rect 170674 74808 170680 74820
rect 170732 74808 170738 74860
rect 172238 74808 172244 74860
rect 172296 74848 172302 74860
rect 373994 74848 374000 74860
rect 172296 74820 374000 74848
rect 172296 74808 172302 74820
rect 373994 74808 374000 74820
rect 374052 74808 374058 74860
rect 172146 74740 172152 74792
rect 172204 74780 172210 74792
rect 396718 74780 396724 74792
rect 172204 74752 396724 74780
rect 172204 74740 172210 74752
rect 396718 74740 396724 74752
rect 396776 74740 396782 74792
rect 170398 74672 170404 74724
rect 170456 74712 170462 74724
rect 170456 74684 170812 74712
rect 170456 74672 170462 74684
rect 170674 74644 170680 74656
rect 169588 74616 170680 74644
rect 170674 74604 170680 74616
rect 170732 74604 170738 74656
rect 170784 74644 170812 74684
rect 172054 74672 172060 74724
rect 172112 74712 172118 74724
rect 396810 74712 396816 74724
rect 172112 74684 396816 74712
rect 172112 74672 172118 74684
rect 396810 74672 396816 74684
rect 396868 74672 396874 74724
rect 462406 74644 462412 74656
rect 170784 74616 462412 74644
rect 462406 74604 462412 74616
rect 462464 74604 462470 74656
rect 160572 74548 164234 74576
rect 164418 74536 164424 74588
rect 164476 74576 164482 74588
rect 170398 74576 170404 74588
rect 164476 74548 170404 74576
rect 164476 74536 164482 74548
rect 170398 74536 170404 74548
rect 170456 74536 170462 74588
rect 170490 74536 170496 74588
rect 170548 74576 170554 74588
rect 550634 74576 550640 74588
rect 170548 74548 550640 74576
rect 170548 74536 170554 74548
rect 550634 74536 550640 74548
rect 550692 74536 550698 74588
rect 161658 74468 161664 74520
rect 161716 74508 161722 74520
rect 167638 74508 167644 74520
rect 161716 74480 167644 74508
rect 161716 74468 161722 74480
rect 167638 74468 167644 74480
rect 167696 74468 167702 74520
rect 168558 74468 168564 74520
rect 168616 74508 168622 74520
rect 175366 74508 175372 74520
rect 168616 74480 175372 74508
rect 168616 74468 168622 74480
rect 175366 74468 175372 74480
rect 175424 74468 175430 74520
rect 580534 74508 580540 74520
rect 175476 74480 580540 74508
rect 153436 74412 160416 74440
rect 153436 74400 153442 74412
rect 167086 74400 167092 74452
rect 167144 74440 167150 74452
rect 175476 74440 175504 74480
rect 580534 74468 580540 74480
rect 580592 74468 580598 74520
rect 580442 74440 580448 74452
rect 167144 74412 175504 74440
rect 176626 74412 580448 74440
rect 167144 74400 167150 74412
rect 111058 74332 111064 74384
rect 111116 74372 111122 74384
rect 113910 74372 113916 74384
rect 111116 74344 113916 74372
rect 111116 74332 111122 74344
rect 113910 74332 113916 74344
rect 113968 74332 113974 74384
rect 157518 74332 157524 74384
rect 157576 74372 157582 74384
rect 164418 74372 164424 74384
rect 157576 74344 164424 74372
rect 157576 74332 157582 74344
rect 164418 74332 164424 74344
rect 164476 74332 164482 74384
rect 167178 74332 167184 74384
rect 167236 74372 167242 74384
rect 176626 74372 176654 74412
rect 580442 74400 580448 74412
rect 580500 74400 580506 74452
rect 167236 74344 176654 74372
rect 167236 74332 167242 74344
rect 115198 74264 115204 74316
rect 115256 74304 115262 74316
rect 170030 74304 170036 74316
rect 115256 74276 170036 74304
rect 115256 74264 115262 74276
rect 170030 74264 170036 74276
rect 170088 74264 170094 74316
rect 140958 74196 140964 74248
rect 141016 74236 141022 74248
rect 249794 74236 249800 74248
rect 141016 74208 249800 74236
rect 141016 74196 141022 74208
rect 249794 74196 249800 74208
rect 249852 74196 249858 74248
rect 143718 74128 143724 74180
rect 143776 74168 143782 74180
rect 284294 74168 284300 74180
rect 143776 74140 284300 74168
rect 143776 74128 143782 74140
rect 284294 74128 284300 74140
rect 284352 74128 284358 74180
rect 146478 74060 146484 74112
rect 146536 74100 146542 74112
rect 320174 74100 320180 74112
rect 146536 74072 320180 74100
rect 146536 74060 146542 74072
rect 320174 74060 320180 74072
rect 320232 74060 320238 74112
rect 147858 73992 147864 74044
rect 147916 74032 147922 74044
rect 338114 74032 338120 74044
rect 147916 74004 338120 74032
rect 147916 73992 147922 74004
rect 338114 73992 338120 74004
rect 338172 73992 338178 74044
rect 151998 73924 152004 73976
rect 152056 73964 152062 73976
rect 390554 73964 390560 73976
rect 152056 73936 390560 73964
rect 152056 73924 152062 73936
rect 390554 73924 390560 73936
rect 390612 73924 390618 73976
rect 116578 73856 116584 73908
rect 116636 73896 116642 73908
rect 116636 73868 162072 73896
rect 116636 73856 116642 73868
rect 157794 73788 157800 73840
rect 157852 73828 157858 73840
rect 161658 73828 161664 73840
rect 157852 73800 161664 73828
rect 157852 73788 157858 73800
rect 161658 73788 161664 73800
rect 161716 73788 161722 73840
rect 112438 73720 112444 73772
rect 112496 73760 112502 73772
rect 162044 73760 162072 73868
rect 168374 73856 168380 73908
rect 168432 73896 168438 73908
rect 462314 73896 462320 73908
rect 168432 73868 462320 73896
rect 168432 73856 168438 73868
rect 462314 73856 462320 73868
rect 462372 73856 462378 73908
rect 164418 73788 164424 73840
rect 164476 73828 164482 73840
rect 465166 73828 465172 73840
rect 164476 73800 465172 73828
rect 164476 73788 164482 73800
rect 465166 73788 465172 73800
rect 465224 73788 465230 73840
rect 170122 73760 170128 73772
rect 112496 73732 161980 73760
rect 162044 73732 170128 73760
rect 112496 73720 112502 73732
rect 5258 73652 5264 73704
rect 5316 73692 5322 73704
rect 161952 73692 161980 73732
rect 170122 73720 170128 73732
rect 170180 73720 170186 73772
rect 169938 73692 169944 73704
rect 5316 73664 160094 73692
rect 161952 73664 169944 73692
rect 5316 73652 5322 73664
rect 44818 73584 44824 73636
rect 44876 73624 44882 73636
rect 44876 73596 157334 73624
rect 44876 73584 44882 73596
rect 157306 73420 157334 73596
rect 160066 73488 160094 73664
rect 169938 73652 169944 73664
rect 169996 73652 170002 73704
rect 167730 73584 167736 73636
rect 167788 73624 167794 73636
rect 172146 73624 172152 73636
rect 167788 73596 172152 73624
rect 167788 73584 167794 73596
rect 172146 73584 172152 73596
rect 172204 73584 172210 73636
rect 161658 73516 161664 73568
rect 161716 73556 161722 73568
rect 167454 73556 167460 73568
rect 161716 73528 167460 73556
rect 161716 73516 161722 73528
rect 167454 73516 167460 73528
rect 167512 73516 167518 73568
rect 167546 73516 167552 73568
rect 167604 73556 167610 73568
rect 172054 73556 172060 73568
rect 167604 73528 172060 73556
rect 167604 73516 167610 73528
rect 172054 73516 172060 73528
rect 172112 73516 172118 73568
rect 169662 73488 169668 73500
rect 160066 73460 169668 73488
rect 169662 73448 169668 73460
rect 169720 73448 169726 73500
rect 169846 73420 169852 73432
rect 157306 73392 169852 73420
rect 169846 73380 169852 73392
rect 169904 73380 169910 73432
rect 151998 73312 152004 73364
rect 152056 73352 152062 73364
rect 152182 73352 152188 73364
rect 152056 73324 152188 73352
rect 152056 73312 152062 73324
rect 152182 73312 152188 73324
rect 152240 73312 152246 73364
rect 162320 73324 169754 73352
rect 84838 73176 84844 73228
rect 84896 73216 84902 73228
rect 84896 73188 85620 73216
rect 84896 73176 84902 73188
rect 85592 73148 85620 73188
rect 152182 73176 152188 73228
rect 152240 73216 152246 73228
rect 152734 73216 152740 73228
rect 152240 73188 152740 73216
rect 152240 73176 152246 73188
rect 152734 73176 152740 73188
rect 152792 73176 152798 73228
rect 162320 73216 162348 73324
rect 162394 73244 162400 73296
rect 162452 73284 162458 73296
rect 162452 73256 162900 73284
rect 162452 73244 162458 73256
rect 162320 73188 162716 73216
rect 92474 73148 92480 73160
rect 85592 73120 92480 73148
rect 92474 73108 92480 73120
rect 92532 73108 92538 73160
rect 118602 73108 118608 73160
rect 118660 73148 118666 73160
rect 120074 73148 120080 73160
rect 118660 73120 120080 73148
rect 118660 73108 118666 73120
rect 120074 73108 120080 73120
rect 120132 73108 120138 73160
rect 120902 73108 120908 73160
rect 120960 73148 120966 73160
rect 127894 73148 127900 73160
rect 120960 73120 127900 73148
rect 120960 73108 120966 73120
rect 127894 73108 127900 73120
rect 127952 73108 127958 73160
rect 136818 73108 136824 73160
rect 136876 73148 136882 73160
rect 161658 73148 161664 73160
rect 136876 73120 161664 73148
rect 136876 73108 136882 73120
rect 161658 73108 161664 73120
rect 161716 73108 161722 73160
rect 137646 73040 137652 73092
rect 137704 73080 137710 73092
rect 162688 73080 162716 73188
rect 162872 73154 162900 73256
rect 169726 73216 169754 73324
rect 207014 73216 207020 73228
rect 169726 73188 207020 73216
rect 207014 73176 207020 73188
rect 207072 73176 207078 73228
rect 162780 73148 162900 73154
rect 164418 73148 164424 73160
rect 162780 73120 164424 73148
rect 164418 73108 164424 73120
rect 164476 73108 164482 73160
rect 166718 73108 166724 73160
rect 166776 73148 166782 73160
rect 172882 73148 172888 73160
rect 166776 73120 172888 73148
rect 166776 73108 166782 73120
rect 172882 73108 172888 73120
rect 172940 73108 172946 73160
rect 137704 73052 162716 73080
rect 137704 73040 137710 73052
rect 165062 73040 165068 73092
rect 165120 73080 165126 73092
rect 167730 73080 167736 73092
rect 165120 73052 167736 73080
rect 165120 73040 165126 73052
rect 167730 73040 167736 73052
rect 167788 73040 167794 73092
rect 167822 73040 167828 73092
rect 167880 73080 167886 73092
rect 580718 73080 580724 73092
rect 167880 73052 580724 73080
rect 167880 73040 167886 73052
rect 580718 73040 580724 73052
rect 580776 73040 580782 73092
rect 120718 72972 120724 73024
rect 120776 73012 120782 73024
rect 128170 73012 128176 73024
rect 120776 72984 128176 73012
rect 120776 72972 120782 72984
rect 128170 72972 128176 72984
rect 128228 72972 128234 73024
rect 136266 72972 136272 73024
rect 136324 73012 136330 73024
rect 168098 73012 168104 73024
rect 136324 72984 168104 73012
rect 136324 72972 136330 72984
rect 168098 72972 168104 72984
rect 168156 72972 168162 73024
rect 168466 72972 168472 73024
rect 168524 73012 168530 73024
rect 397454 73012 397460 73024
rect 168524 72984 397460 73012
rect 168524 72972 168530 72984
rect 397454 72972 397460 72984
rect 397512 72972 397518 73024
rect 120810 72904 120816 72956
rect 120868 72944 120874 72956
rect 129274 72944 129280 72956
rect 120868 72916 129280 72944
rect 120868 72904 120874 72916
rect 129274 72904 129280 72916
rect 129332 72904 129338 72956
rect 141602 72904 141608 72956
rect 141660 72944 141666 72956
rect 146754 72944 146760 72956
rect 141660 72916 146760 72944
rect 141660 72904 141666 72916
rect 146754 72904 146760 72916
rect 146812 72904 146818 72956
rect 154390 72904 154396 72956
rect 154448 72944 154454 72956
rect 422294 72944 422300 72956
rect 154448 72916 422300 72944
rect 154448 72904 154454 72916
rect 422294 72904 422300 72916
rect 422352 72904 422358 72956
rect 121086 72836 121092 72888
rect 121144 72876 121150 72888
rect 130378 72876 130384 72888
rect 121144 72848 130384 72876
rect 121144 72836 121150 72848
rect 130378 72836 130384 72848
rect 130436 72836 130442 72888
rect 142154 72836 142160 72888
rect 142212 72876 142218 72888
rect 152734 72876 152740 72888
rect 142212 72848 152740 72876
rect 142212 72836 142218 72848
rect 152734 72836 152740 72848
rect 152792 72836 152798 72888
rect 156046 72836 156052 72888
rect 156104 72876 156110 72888
rect 442994 72876 443000 72888
rect 156104 72848 443000 72876
rect 156104 72836 156110 72848
rect 442994 72836 443000 72848
rect 443052 72836 443058 72888
rect 149146 72768 149152 72820
rect 149204 72808 149210 72820
rect 154390 72808 154396 72820
rect 149204 72780 154396 72808
rect 149204 72768 149210 72780
rect 154390 72768 154396 72780
rect 154448 72768 154454 72820
rect 156598 72768 156604 72820
rect 156656 72808 156662 72820
rect 449894 72808 449900 72820
rect 156656 72780 449900 72808
rect 156656 72768 156662 72780
rect 449894 72768 449900 72780
rect 449952 72768 449958 72820
rect 120994 72700 121000 72752
rect 121052 72740 121058 72752
rect 129826 72740 129832 72752
rect 121052 72712 129832 72740
rect 121052 72700 121058 72712
rect 129826 72700 129832 72712
rect 129884 72700 129890 72752
rect 140498 72700 140504 72752
rect 140556 72740 140562 72752
rect 151630 72740 151636 72752
rect 140556 72712 151636 72740
rect 140556 72700 140562 72712
rect 151630 72700 151636 72712
rect 151688 72700 151694 72752
rect 151998 72700 152004 72752
rect 152056 72740 152062 72752
rect 152056 72712 157334 72740
rect 152056 72700 152062 72712
rect 121362 72632 121368 72684
rect 121420 72672 121426 72684
rect 132678 72672 132684 72684
rect 121420 72644 132684 72672
rect 121420 72632 121426 72644
rect 132678 72632 132684 72644
rect 132736 72632 132742 72684
rect 138842 72632 138848 72684
rect 138900 72672 138906 72684
rect 146478 72672 146484 72684
rect 138900 72644 146484 72672
rect 138900 72632 138906 72644
rect 146478 72632 146484 72644
rect 146536 72632 146542 72684
rect 150250 72632 150256 72684
rect 150308 72672 150314 72684
rect 150308 72644 154344 72672
rect 150308 72632 150314 72644
rect 132310 72564 132316 72616
rect 132368 72604 132374 72616
rect 137738 72604 137744 72616
rect 132368 72576 137744 72604
rect 132368 72564 132374 72576
rect 137738 72564 137744 72576
rect 137796 72564 137802 72616
rect 139210 72564 139216 72616
rect 139268 72604 139274 72616
rect 139268 72576 150388 72604
rect 139268 72564 139274 72576
rect 60734 72496 60740 72548
rect 60792 72536 60798 72548
rect 126330 72536 126336 72548
rect 60792 72508 126336 72536
rect 60792 72496 60798 72508
rect 126330 72496 126336 72508
rect 126388 72496 126394 72548
rect 134702 72496 134708 72548
rect 134760 72536 134766 72548
rect 149146 72536 149152 72548
rect 134760 72508 149152 72536
rect 134760 72496 134766 72508
rect 149146 72496 149152 72508
rect 149204 72496 149210 72548
rect 150360 72536 150388 72576
rect 151262 72564 151268 72616
rect 151320 72604 151326 72616
rect 154206 72604 154212 72616
rect 151320 72576 154212 72604
rect 151320 72564 151326 72576
rect 154206 72564 154212 72576
rect 154264 72564 154270 72616
rect 153102 72536 153108 72548
rect 150360 72508 153108 72536
rect 153102 72496 153108 72508
rect 153160 72496 153166 72548
rect 154316 72536 154344 72644
rect 157306 72604 157334 72712
rect 157426 72700 157432 72752
rect 157484 72740 157490 72752
rect 158806 72740 158812 72752
rect 157484 72712 158812 72740
rect 157484 72700 157490 72712
rect 158806 72700 158812 72712
rect 158864 72700 158870 72752
rect 158916 72712 162624 72740
rect 158254 72632 158260 72684
rect 158312 72672 158318 72684
rect 158916 72672 158944 72712
rect 158312 72644 158944 72672
rect 162596 72672 162624 72712
rect 164418 72700 164424 72752
rect 164476 72740 164482 72752
rect 166350 72740 166356 72752
rect 164476 72712 166356 72740
rect 164476 72700 164482 72712
rect 166350 72700 166356 72712
rect 166408 72700 166414 72752
rect 167730 72700 167736 72752
rect 167788 72740 167794 72752
rect 460934 72740 460940 72752
rect 167788 72712 460940 72740
rect 167788 72700 167794 72712
rect 460934 72700 460940 72712
rect 460992 72700 460998 72752
rect 471974 72672 471980 72684
rect 162596 72644 471980 72672
rect 158312 72632 158318 72644
rect 471974 72632 471980 72644
rect 472032 72632 472038 72684
rect 157306 72576 158484 72604
rect 158254 72536 158260 72548
rect 154316 72508 158260 72536
rect 158254 72496 158260 72508
rect 158312 72496 158318 72548
rect 25498 72428 25504 72480
rect 25556 72468 25562 72480
rect 123110 72468 123116 72480
rect 25556 72440 123116 72468
rect 25556 72428 25562 72440
rect 123110 72428 123116 72440
rect 123168 72428 123174 72480
rect 135714 72428 135720 72480
rect 135772 72468 135778 72480
rect 157518 72468 157524 72480
rect 135772 72440 145604 72468
rect 135772 72428 135778 72440
rect 116578 72360 116584 72412
rect 116636 72400 116642 72412
rect 124858 72400 124864 72412
rect 116636 72372 124864 72400
rect 116636 72360 116642 72372
rect 124858 72360 124864 72372
rect 124916 72360 124922 72412
rect 137646 72360 137652 72412
rect 137704 72400 137710 72412
rect 137704 72372 142154 72400
rect 137704 72360 137710 72372
rect 118142 72292 118148 72344
rect 118200 72332 118206 72344
rect 124306 72332 124312 72344
rect 118200 72304 124312 72332
rect 118200 72292 118206 72304
rect 124306 72292 124312 72304
rect 124364 72292 124370 72344
rect 86218 72224 86224 72276
rect 86276 72264 86282 72276
rect 122374 72264 122380 72276
rect 86276 72236 122380 72264
rect 86276 72224 86282 72236
rect 122374 72224 122380 72236
rect 122432 72224 122438 72276
rect 117958 72156 117964 72208
rect 118016 72196 118022 72208
rect 123754 72196 123760 72208
rect 118016 72168 123760 72196
rect 118016 72156 118022 72168
rect 123754 72156 123760 72168
rect 123812 72156 123818 72208
rect 118050 72088 118056 72140
rect 118108 72128 118114 72140
rect 123018 72128 123024 72140
rect 118108 72100 123024 72128
rect 118108 72088 118114 72100
rect 123018 72088 123024 72100
rect 123076 72088 123082 72140
rect 142126 72060 142154 72372
rect 145576 72332 145604 72440
rect 147140 72440 157524 72468
rect 147140 72332 147168 72440
rect 157518 72428 157524 72440
rect 157576 72428 157582 72480
rect 150802 72360 150808 72412
rect 150860 72400 150866 72412
rect 152918 72400 152924 72412
rect 150860 72372 152924 72400
rect 150860 72360 150866 72372
rect 152918 72360 152924 72372
rect 152976 72360 152982 72412
rect 158456 72400 158484 72576
rect 162486 72564 162492 72616
rect 162544 72604 162550 72616
rect 514754 72604 514760 72616
rect 162544 72576 514760 72604
rect 162544 72564 162550 72576
rect 514754 72564 514760 72576
rect 514812 72564 514818 72616
rect 158806 72496 158812 72548
rect 158864 72536 158870 72548
rect 165062 72536 165068 72548
rect 158864 72508 165068 72536
rect 158864 72496 158870 72508
rect 165062 72496 165068 72508
rect 165120 72496 165126 72548
rect 170582 72496 170588 72548
rect 170640 72536 170646 72548
rect 558914 72536 558920 72548
rect 170640 72508 558920 72536
rect 170640 72496 170646 72508
rect 558914 72496 558920 72508
rect 558972 72496 558978 72548
rect 166626 72428 166632 72480
rect 166684 72468 166690 72480
rect 580994 72468 581000 72480
rect 166684 72440 581000 72468
rect 166684 72428 166690 72440
rect 580994 72428 581000 72440
rect 581052 72428 581058 72480
rect 167362 72400 167368 72412
rect 158456 72372 167368 72400
rect 167362 72360 167368 72372
rect 167420 72360 167426 72412
rect 167914 72360 167920 72412
rect 167972 72400 167978 72412
rect 217318 72400 217324 72412
rect 167972 72372 217324 72400
rect 167972 72360 167978 72372
rect 217318 72360 217324 72372
rect 217376 72360 217382 72412
rect 145576 72304 147168 72332
rect 152182 72292 152188 72344
rect 152240 72332 152246 72344
rect 167454 72332 167460 72344
rect 152240 72304 167460 72332
rect 152240 72292 152246 72304
rect 167454 72292 167460 72304
rect 167512 72292 167518 72344
rect 145466 72224 145472 72276
rect 145524 72264 145530 72276
rect 145524 72236 151032 72264
rect 145524 72224 145530 72236
rect 146478 72156 146484 72208
rect 146536 72196 146542 72208
rect 150158 72196 150164 72208
rect 146536 72168 150164 72196
rect 146536 72156 146542 72168
rect 150158 72156 150164 72168
rect 150216 72156 150222 72208
rect 151004 72196 151032 72236
rect 153838 72224 153844 72276
rect 153896 72264 153902 72276
rect 168282 72264 168288 72276
rect 153896 72236 168288 72264
rect 153896 72224 153902 72236
rect 168282 72224 168288 72236
rect 168340 72224 168346 72276
rect 154390 72196 154396 72208
rect 151004 72168 154396 72196
rect 154390 72156 154396 72168
rect 154448 72156 154454 72208
rect 167730 72196 167736 72208
rect 157306 72168 167736 72196
rect 142706 72088 142712 72140
rect 142764 72128 142770 72140
rect 142764 72100 146248 72128
rect 142764 72088 142770 72100
rect 146018 72060 146024 72072
rect 142126 72032 146024 72060
rect 146018 72020 146024 72032
rect 146076 72020 146082 72072
rect 146220 72060 146248 72100
rect 154942 72088 154948 72140
rect 155000 72128 155006 72140
rect 157306 72128 157334 72168
rect 167730 72156 167736 72168
rect 167788 72156 167794 72208
rect 167546 72128 167552 72140
rect 155000 72100 157334 72128
rect 162136 72100 167552 72128
rect 155000 72088 155006 72100
rect 153010 72060 153016 72072
rect 146220 72032 153016 72060
rect 153010 72020 153016 72032
rect 153068 72020 153074 72072
rect 153286 72020 153292 72072
rect 153344 72060 153350 72072
rect 162136 72060 162164 72100
rect 167546 72088 167552 72100
rect 167604 72088 167610 72140
rect 178862 72060 178868 72072
rect 153344 72032 162164 72060
rect 166966 72032 178868 72060
rect 153344 72020 153350 72032
rect 151906 71952 151912 72004
rect 151964 71992 151970 72004
rect 155770 71992 155776 72004
rect 151964 71964 155776 71992
rect 151964 71952 151970 71964
rect 155770 71952 155776 71964
rect 155828 71952 155834 72004
rect 146754 71884 146760 71936
rect 146812 71924 146818 71936
rect 151538 71924 151544 71936
rect 146812 71896 151544 71924
rect 146812 71884 146818 71896
rect 151538 71884 151544 71896
rect 151596 71884 151602 71936
rect 151814 71884 151820 71936
rect 151872 71924 151878 71936
rect 157150 71924 157156 71936
rect 151872 71896 157156 71924
rect 151872 71884 151878 71896
rect 157150 71884 157156 71896
rect 157208 71884 157214 71936
rect 157518 71884 157524 71936
rect 157576 71924 157582 71936
rect 165246 71924 165252 71936
rect 157576 71896 165252 71924
rect 157576 71884 157582 71896
rect 165246 71884 165252 71896
rect 165304 71884 165310 71936
rect 119338 71816 119344 71868
rect 119396 71856 119402 71868
rect 122742 71856 122748 71868
rect 119396 71828 122748 71856
rect 119396 71816 119402 71828
rect 122742 71816 122748 71828
rect 122800 71816 122806 71868
rect 132494 71816 132500 71868
rect 132552 71856 132558 71868
rect 136266 71856 136272 71868
rect 132552 71828 136272 71856
rect 132552 71816 132558 71828
rect 136266 71816 136272 71828
rect 136324 71816 136330 71868
rect 136634 71816 136640 71868
rect 136692 71856 136698 71868
rect 136692 71828 142154 71856
rect 136692 71816 136698 71828
rect 122374 71748 122380 71800
rect 122432 71788 122438 71800
rect 127342 71788 127348 71800
rect 122432 71760 127348 71788
rect 122432 71748 122438 71760
rect 127342 71748 127348 71760
rect 127400 71748 127406 71800
rect 133966 71748 133972 71800
rect 134024 71788 134030 71800
rect 137646 71788 137652 71800
rect 134024 71760 137652 71788
rect 134024 71748 134030 71760
rect 137646 71748 137652 71760
rect 137704 71748 137710 71800
rect 142126 71788 142154 71828
rect 151354 71816 151360 71868
rect 151412 71856 151418 71868
rect 158438 71856 158444 71868
rect 151412 71828 158444 71856
rect 151412 71816 151418 71828
rect 158438 71816 158444 71828
rect 158496 71816 158502 71868
rect 143166 71788 143172 71800
rect 142126 71760 143172 71788
rect 143166 71748 143172 71760
rect 143224 71748 143230 71800
rect 145834 71748 145840 71800
rect 145892 71788 145898 71800
rect 147306 71788 147312 71800
rect 145892 71760 147312 71788
rect 145892 71748 145898 71760
rect 147306 71748 147312 71760
rect 147364 71748 147370 71800
rect 149698 71748 149704 71800
rect 149756 71788 149762 71800
rect 156966 71788 156972 71800
rect 149756 71760 156972 71788
rect 149756 71748 149762 71760
rect 156966 71748 156972 71760
rect 157024 71748 157030 71800
rect 3510 71680 3516 71732
rect 3568 71720 3574 71732
rect 166966 71720 166994 72032
rect 178862 72020 178868 72032
rect 178920 72020 178926 72072
rect 167086 71952 167092 72004
rect 167144 71992 167150 72004
rect 580166 71992 580172 72004
rect 167144 71964 580172 71992
rect 167144 71952 167150 71964
rect 580166 71952 580172 71964
rect 580224 71952 580230 72004
rect 3568 71692 166994 71720
rect 3568 71680 3574 71692
rect 6914 71612 6920 71664
rect 6972 71652 6978 71664
rect 169018 71652 169024 71664
rect 6972 71624 169024 71652
rect 6972 71612 6978 71624
rect 169018 71612 169024 71624
rect 169076 71612 169082 71664
rect 92474 71544 92480 71596
rect 92532 71584 92538 71596
rect 168650 71584 168656 71596
rect 92532 71556 168656 71584
rect 92532 71544 92538 71556
rect 168650 71544 168656 71556
rect 168708 71544 168714 71596
rect 104158 71476 104164 71528
rect 104216 71516 104222 71528
rect 168926 71516 168932 71528
rect 104216 71488 168932 71516
rect 104216 71476 104222 71488
rect 168926 71476 168932 71488
rect 168984 71476 168990 71528
rect 113910 71408 113916 71460
rect 113968 71448 113974 71460
rect 168742 71448 168748 71460
rect 113968 71420 168748 71448
rect 113968 71408 113974 71420
rect 168742 71408 168748 71420
rect 168800 71408 168806 71460
rect 120074 71340 120080 71392
rect 120132 71380 120138 71392
rect 168834 71380 168840 71392
rect 120132 71352 168840 71380
rect 120132 71340 120138 71352
rect 168834 71340 168840 71352
rect 168892 71340 168898 71392
rect 166902 71000 166908 71052
rect 166960 71040 166966 71052
rect 580258 71040 580264 71052
rect 166960 71012 580264 71040
rect 166960 71000 166966 71012
rect 580258 71000 580264 71012
rect 580316 71000 580322 71052
rect 122926 70048 122932 70100
rect 122984 70088 122990 70100
rect 124122 70088 124128 70100
rect 122984 70060 124128 70088
rect 122984 70048 122990 70060
rect 124122 70048 124128 70060
rect 124180 70048 124186 70100
rect 131206 70048 131212 70100
rect 131264 70088 131270 70100
rect 131574 70088 131580 70100
rect 131264 70060 131580 70088
rect 131264 70048 131270 70060
rect 131574 70048 131580 70060
rect 131632 70048 131638 70100
rect 121546 69980 121552 70032
rect 121604 70020 121610 70032
rect 122558 70020 122564 70032
rect 121604 69992 122564 70020
rect 121604 69980 121610 69992
rect 122558 69980 122564 69992
rect 122616 69980 122622 70032
rect 123018 69980 123024 70032
rect 123076 70020 123082 70032
rect 123846 70020 123852 70032
rect 123076 69992 123852 70020
rect 123076 69980 123082 69992
rect 123846 69980 123852 69992
rect 123904 69980 123910 70032
rect 124306 69980 124312 70032
rect 124364 70020 124370 70032
rect 125226 70020 125232 70032
rect 124364 69992 125232 70020
rect 124364 69980 124370 69992
rect 125226 69980 125232 69992
rect 125284 69980 125290 70032
rect 128538 69980 128544 70032
rect 128596 70020 128602 70032
rect 129366 70020 129372 70032
rect 128596 69992 129372 70020
rect 128596 69980 128602 69992
rect 129366 69980 129372 69992
rect 129424 69980 129430 70032
rect 123202 69912 123208 69964
rect 123260 69952 123266 69964
rect 123662 69952 123668 69964
rect 123260 69924 123668 69952
rect 123260 69912 123266 69924
rect 123662 69912 123668 69924
rect 123720 69912 123726 69964
rect 129182 69912 129188 69964
rect 129240 69912 129246 69964
rect 130102 69912 130108 69964
rect 130160 69952 130166 69964
rect 130378 69952 130384 69964
rect 130160 69924 130384 69952
rect 130160 69912 130166 69924
rect 130378 69912 130384 69924
rect 130436 69912 130442 69964
rect 121454 69844 121460 69896
rect 121512 69884 121518 69896
rect 122006 69884 122012 69896
rect 121512 69856 122012 69884
rect 121512 69844 121518 69856
rect 122006 69844 122012 69856
rect 122064 69844 122070 69896
rect 122098 69844 122104 69896
rect 122156 69884 122162 69896
rect 122558 69884 122564 69896
rect 122156 69856 122564 69884
rect 122156 69844 122162 69856
rect 122558 69844 122564 69856
rect 122616 69844 122622 69896
rect 123570 69844 123576 69896
rect 123628 69884 123634 69896
rect 124122 69884 124128 69896
rect 123628 69856 124128 69884
rect 123628 69844 123634 69856
rect 124122 69844 124128 69856
rect 124180 69844 124186 69896
rect 124582 69844 124588 69896
rect 124640 69884 124646 69896
rect 125226 69884 125232 69896
rect 124640 69856 125232 69884
rect 124640 69844 124646 69856
rect 125226 69844 125232 69856
rect 125284 69844 125290 69896
rect 121730 69776 121736 69828
rect 121788 69816 121794 69828
rect 122190 69816 122196 69828
rect 121788 69788 122196 69816
rect 121788 69776 121794 69788
rect 122190 69776 122196 69788
rect 122248 69776 122254 69828
rect 123938 69816 123944 69828
rect 123496 69788 123944 69816
rect 123496 69624 123524 69788
rect 123938 69776 123944 69788
rect 123996 69776 124002 69828
rect 124490 69776 124496 69828
rect 124548 69816 124554 69828
rect 124950 69816 124956 69828
rect 124548 69788 124956 69816
rect 124548 69776 124554 69788
rect 124950 69776 124956 69788
rect 125008 69776 125014 69828
rect 127066 69776 127072 69828
rect 127124 69816 127130 69828
rect 127710 69816 127716 69828
rect 127124 69788 127716 69816
rect 127124 69776 127130 69788
rect 127710 69776 127716 69788
rect 127768 69776 127774 69828
rect 125686 69708 125692 69760
rect 125744 69748 125750 69760
rect 126606 69748 126612 69760
rect 125744 69720 126612 69748
rect 125744 69708 125750 69720
rect 126606 69708 126612 69720
rect 126664 69708 126670 69760
rect 129200 69692 129228 69912
rect 130470 69816 130476 69828
rect 130028 69788 130476 69816
rect 130028 69760 130056 69788
rect 130470 69776 130476 69788
rect 130528 69776 130534 69828
rect 138106 69776 138112 69828
rect 138164 69816 138170 69828
rect 138842 69816 138848 69828
rect 138164 69788 138848 69816
rect 138164 69776 138170 69788
rect 138842 69776 138848 69788
rect 138900 69776 138906 69828
rect 130010 69708 130016 69760
rect 130068 69708 130074 69760
rect 125778 69640 125784 69692
rect 125836 69680 125842 69692
rect 126422 69680 126428 69692
rect 125836 69652 126428 69680
rect 125836 69640 125842 69652
rect 126422 69640 126428 69652
rect 126480 69640 126486 69692
rect 129182 69640 129188 69692
rect 129240 69640 129246 69692
rect 130470 69640 130476 69692
rect 130528 69680 130534 69692
rect 130930 69680 130936 69692
rect 130528 69652 130936 69680
rect 130528 69640 130534 69652
rect 130930 69640 130936 69652
rect 130988 69640 130994 69692
rect 131114 69640 131120 69692
rect 131172 69680 131178 69692
rect 131758 69680 131764 69692
rect 131172 69652 131764 69680
rect 131172 69640 131178 69652
rect 131758 69640 131764 69652
rect 131816 69640 131822 69692
rect 122098 69572 122104 69624
rect 122156 69612 122162 69624
rect 122650 69612 122656 69624
rect 122156 69584 122656 69612
rect 122156 69572 122162 69584
rect 122650 69572 122656 69584
rect 122708 69572 122714 69624
rect 123478 69572 123484 69624
rect 123536 69572 123542 69624
rect 127158 69572 127164 69624
rect 127216 69612 127222 69624
rect 127434 69612 127440 69624
rect 127216 69584 127440 69612
rect 127216 69572 127222 69584
rect 127434 69572 127440 69584
rect 127492 69572 127498 69624
rect 128814 69572 128820 69624
rect 128872 69612 128878 69624
rect 129274 69612 129280 69624
rect 128872 69584 129280 69612
rect 128872 69572 128878 69584
rect 129274 69572 129280 69584
rect 129332 69572 129338 69624
rect 130194 69572 130200 69624
rect 130252 69612 130258 69624
rect 130562 69612 130568 69624
rect 130252 69584 130568 69612
rect 130252 69572 130258 69584
rect 130562 69572 130568 69584
rect 130620 69572 130626 69624
rect 123110 69504 123116 69556
rect 123168 69544 123174 69556
rect 123754 69544 123760 69556
rect 123168 69516 123760 69544
rect 123168 69504 123174 69516
rect 123754 69504 123760 69516
rect 123812 69504 123818 69556
rect 127342 69504 127348 69556
rect 127400 69544 127406 69556
rect 127618 69544 127624 69556
rect 127400 69516 127624 69544
rect 127400 69504 127406 69516
rect 127618 69504 127624 69516
rect 127676 69504 127682 69556
rect 130102 69504 130108 69556
rect 130160 69544 130166 69556
rect 130838 69544 130844 69556
rect 130160 69516 130844 69544
rect 130160 69504 130166 69516
rect 130838 69504 130844 69516
rect 130896 69504 130902 69556
rect 131298 69504 131304 69556
rect 131356 69544 131362 69556
rect 131356 69516 131436 69544
rect 131356 69504 131362 69516
rect 124858 69436 124864 69488
rect 124916 69476 124922 69488
rect 125410 69476 125416 69488
rect 124916 69448 125416 69476
rect 124916 69436 124922 69448
rect 125410 69436 125416 69448
rect 125468 69436 125474 69488
rect 131408 69352 131436 69516
rect 131574 69368 131580 69420
rect 131632 69368 131638 69420
rect 126422 69300 126428 69352
rect 126480 69340 126486 69352
rect 126790 69340 126796 69352
rect 126480 69312 126796 69340
rect 126480 69300 126486 69312
rect 126790 69300 126796 69312
rect 126848 69300 126854 69352
rect 127434 69300 127440 69352
rect 127492 69340 127498 69352
rect 127894 69340 127900 69352
rect 127492 69312 127900 69340
rect 127492 69300 127498 69312
rect 127894 69300 127900 69312
rect 127952 69300 127958 69352
rect 131390 69300 131396 69352
rect 131448 69300 131454 69352
rect 127342 69232 127348 69284
rect 127400 69272 127406 69284
rect 128262 69272 128268 69284
rect 127400 69244 128268 69272
rect 127400 69232 127406 69244
rect 128262 69232 128268 69244
rect 128320 69232 128326 69284
rect 131592 69216 131620 69368
rect 126054 69164 126060 69216
rect 126112 69204 126118 69216
rect 126514 69204 126520 69216
rect 126112 69176 126520 69204
rect 126112 69164 126118 69176
rect 126514 69164 126520 69176
rect 126572 69164 126578 69216
rect 131574 69164 131580 69216
rect 131632 69164 131638 69216
rect 127710 69096 127716 69148
rect 127768 69136 127774 69148
rect 128078 69136 128084 69148
rect 127768 69108 128084 69136
rect 127768 69096 127774 69108
rect 128078 69096 128084 69108
rect 128136 69096 128142 69148
rect 121638 68212 121644 68264
rect 121696 68252 121702 68264
rect 122282 68252 122288 68264
rect 121696 68224 122288 68252
rect 121696 68212 121702 68224
rect 122282 68212 122288 68224
rect 122340 68212 122346 68264
rect 125962 67804 125968 67856
rect 126020 67844 126026 67856
rect 126238 67844 126244 67856
rect 126020 67816 126244 67844
rect 126020 67804 126026 67816
rect 126238 67804 126244 67816
rect 126296 67804 126302 67856
rect 129918 67600 129924 67652
rect 129976 67640 129982 67652
rect 130746 67640 130752 67652
rect 129976 67612 130752 67640
rect 129976 67600 129982 67612
rect 130746 67600 130752 67612
rect 130804 67600 130810 67652
rect 125778 67532 125784 67584
rect 125836 67572 125842 67584
rect 125962 67572 125968 67584
rect 125836 67544 125968 67572
rect 125836 67532 125842 67544
rect 125962 67532 125968 67544
rect 126020 67532 126026 67584
rect 126054 67532 126060 67584
rect 126112 67572 126118 67584
rect 126698 67572 126704 67584
rect 126112 67544 126704 67572
rect 126112 67532 126118 67544
rect 126698 67532 126704 67544
rect 126756 67532 126762 67584
rect 124674 67328 124680 67380
rect 124732 67368 124738 67380
rect 125318 67368 125324 67380
rect 124732 67340 125324 67368
rect 124732 67328 124738 67340
rect 125318 67328 125324 67340
rect 125376 67328 125382 67380
rect 5534 66852 5540 66904
rect 5592 66892 5598 66904
rect 121454 66892 121460 66904
rect 5592 66864 121460 66892
rect 5592 66852 5598 66864
rect 121454 66852 121460 66864
rect 121512 66852 121518 66904
rect 124766 65900 124772 65952
rect 124824 65940 124830 65952
rect 125042 65940 125048 65952
rect 124824 65912 125048 65940
rect 124824 65900 124830 65912
rect 125042 65900 125048 65912
rect 125100 65900 125106 65952
rect 128814 65628 128820 65680
rect 128872 65668 128878 65680
rect 129458 65668 129464 65680
rect 128872 65640 129464 65668
rect 128872 65628 128878 65640
rect 129458 65628 129464 65640
rect 129516 65628 129522 65680
rect 128906 65560 128912 65612
rect 128964 65600 128970 65612
rect 129182 65600 129188 65612
rect 128964 65572 129188 65600
rect 128964 65560 128970 65572
rect 129182 65560 129188 65572
rect 129240 65560 129246 65612
rect 129090 65492 129096 65544
rect 129148 65532 129154 65544
rect 129550 65532 129556 65544
rect 129148 65504 129556 65532
rect 129148 65492 129154 65504
rect 129550 65492 129556 65504
rect 129608 65492 129614 65544
rect 128630 65424 128636 65476
rect 128688 65464 128694 65476
rect 129182 65464 129188 65476
rect 128688 65436 129188 65464
rect 128688 65424 128694 65436
rect 129182 65424 129188 65436
rect 129240 65424 129246 65476
rect 128630 65288 128636 65340
rect 128688 65328 128694 65340
rect 129642 65328 129648 65340
rect 128688 65300 129648 65328
rect 128688 65288 128694 65300
rect 129642 65288 129648 65300
rect 129700 65288 129706 65340
rect 114370 60664 114376 60716
rect 114428 60704 114434 60716
rect 580166 60704 580172 60716
rect 114428 60676 580172 60704
rect 114428 60664 114434 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 163498 58624 163504 58676
rect 163556 58664 163562 58676
rect 326338 58664 326344 58676
rect 163556 58636 326344 58664
rect 163556 58624 163562 58636
rect 326338 58624 326344 58636
rect 326396 58624 326402 58676
rect 15194 54476 15200 54528
rect 15252 54516 15258 54528
rect 119338 54516 119344 54528
rect 15252 54488 119344 54516
rect 15252 54476 15258 54488
rect 119338 54476 119344 54488
rect 119396 54476 119402 54528
rect 113174 51076 113180 51128
rect 113232 51116 113238 51128
rect 121086 51116 121092 51128
rect 113232 51088 121092 51116
rect 113232 51076 113238 51088
rect 121086 51076 121092 51088
rect 121144 51076 121150 51128
rect 178678 46860 178684 46912
rect 178736 46900 178742 46912
rect 580166 46900 580172 46912
rect 178736 46872 580172 46900
rect 178736 46860 178742 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 170214 45540 170220 45552
rect 3568 45512 170220 45540
rect 3568 45500 3574 45512
rect 170214 45500 170220 45512
rect 170272 45500 170278 45552
rect 106274 43392 106280 43444
rect 106332 43432 106338 43444
rect 120994 43432 121000 43444
rect 106332 43404 121000 43432
rect 106332 43392 106338 43404
rect 120994 43392 121000 43404
rect 121052 43392 121058 43444
rect 153102 40672 153108 40724
rect 153160 40712 153166 40724
rect 226334 40712 226340 40724
rect 153160 40684 226340 40712
rect 153160 40672 153166 40684
rect 226334 40672 226340 40684
rect 226392 40672 226398 40724
rect 158438 36660 158444 36712
rect 158496 36700 158502 36712
rect 382274 36700 382280 36712
rect 158496 36672 382280 36700
rect 158496 36660 158502 36672
rect 382274 36660 382280 36672
rect 382332 36660 382338 36712
rect 155770 36592 155776 36644
rect 155828 36632 155834 36644
rect 390646 36632 390652 36644
rect 155828 36604 390652 36632
rect 155828 36592 155834 36604
rect 390646 36592 390652 36604
rect 390704 36592 390710 36644
rect 152458 36524 152464 36576
rect 152516 36564 152522 36576
rect 397454 36564 397460 36576
rect 152516 36536 397460 36564
rect 152516 36524 152522 36536
rect 397454 36524 397460 36536
rect 397512 36524 397518 36576
rect 145558 35844 145564 35896
rect 145616 35884 145622 35896
rect 307754 35884 307760 35896
rect 145616 35856 307760 35884
rect 145616 35844 145622 35856
rect 307754 35844 307760 35856
rect 307812 35844 307818 35896
rect 147306 35776 147312 35828
rect 147364 35816 147370 35828
rect 311894 35816 311900 35828
rect 147364 35788 311900 35816
rect 147364 35776 147370 35788
rect 311894 35776 311900 35788
rect 311952 35776 311958 35828
rect 146386 35708 146392 35760
rect 146444 35748 146450 35760
rect 318794 35748 318800 35760
rect 146444 35720 318800 35748
rect 146444 35708 146450 35720
rect 318794 35708 318800 35720
rect 318852 35708 318858 35760
rect 146662 35640 146668 35692
rect 146720 35680 146726 35692
rect 322934 35680 322940 35692
rect 146720 35652 322940 35680
rect 146720 35640 146726 35652
rect 322934 35640 322940 35652
rect 322992 35640 322998 35692
rect 146938 35572 146944 35624
rect 146996 35612 147002 35624
rect 325694 35612 325700 35624
rect 146996 35584 325700 35612
rect 146996 35572 147002 35584
rect 325694 35572 325700 35584
rect 325752 35572 325758 35624
rect 147766 35504 147772 35556
rect 147824 35544 147830 35556
rect 336734 35544 336740 35556
rect 147824 35516 336740 35544
rect 147824 35504 147830 35516
rect 336734 35504 336740 35516
rect 336792 35504 336798 35556
rect 148594 35436 148600 35488
rect 148652 35476 148658 35488
rect 347774 35476 347780 35488
rect 148652 35448 347780 35476
rect 148652 35436 148658 35448
rect 347774 35436 347780 35448
rect 347832 35436 347838 35488
rect 154482 35368 154488 35420
rect 154540 35408 154546 35420
rect 354674 35408 354680 35420
rect 154540 35380 354680 35408
rect 154540 35368 154546 35380
rect 354674 35368 354680 35380
rect 354732 35368 354738 35420
rect 149422 35300 149428 35352
rect 149480 35340 149486 35352
rect 357434 35340 357440 35352
rect 149480 35312 357440 35340
rect 149480 35300 149486 35312
rect 357434 35300 357440 35312
rect 357492 35300 357498 35352
rect 158346 35232 158352 35284
rect 158404 35272 158410 35284
rect 368474 35272 368480 35284
rect 158404 35244 368480 35272
rect 158404 35232 158410 35244
rect 368474 35232 368480 35244
rect 368532 35232 368538 35284
rect 157794 35164 157800 35216
rect 157852 35204 157858 35216
rect 456794 35204 456800 35216
rect 157852 35176 456800 35204
rect 157852 35164 157858 35176
rect 456794 35164 456800 35176
rect 456852 35164 456858 35216
rect 145282 35096 145288 35148
rect 145340 35136 145346 35148
rect 304994 35136 305000 35148
rect 145340 35108 305000 35136
rect 145340 35096 145346 35108
rect 304994 35096 305000 35108
rect 305052 35096 305058 35148
rect 138842 34416 138848 34468
rect 138900 34456 138906 34468
rect 212534 34456 212540 34468
rect 138900 34428 212540 34456
rect 138900 34416 138906 34428
rect 212534 34416 212540 34428
rect 212592 34416 212598 34468
rect 138382 34348 138388 34400
rect 138440 34388 138446 34400
rect 216674 34388 216680 34400
rect 138440 34360 216680 34388
rect 138440 34348 138446 34360
rect 216674 34348 216680 34360
rect 216732 34348 216738 34400
rect 138658 34280 138664 34332
rect 138716 34320 138722 34332
rect 219434 34320 219440 34332
rect 138716 34292 219440 34320
rect 138716 34280 138722 34292
rect 219434 34280 219440 34292
rect 219492 34280 219498 34332
rect 139762 34212 139768 34264
rect 139820 34252 139826 34264
rect 234614 34252 234620 34264
rect 139820 34224 234620 34252
rect 139820 34212 139826 34224
rect 234614 34212 234620 34224
rect 234672 34212 234678 34264
rect 140866 34144 140872 34196
rect 140924 34184 140930 34196
rect 248414 34184 248420 34196
rect 140924 34156 248420 34184
rect 140924 34144 140930 34156
rect 248414 34144 248420 34156
rect 248472 34144 248478 34196
rect 141418 34076 141424 34128
rect 141476 34116 141482 34128
rect 255314 34116 255320 34128
rect 141476 34088 255320 34116
rect 141476 34076 141482 34088
rect 255314 34076 255320 34088
rect 255372 34076 255378 34128
rect 142522 34008 142528 34060
rect 142580 34048 142586 34060
rect 269114 34048 269120 34060
rect 142580 34020 269120 34048
rect 142580 34008 142586 34020
rect 269114 34008 269120 34020
rect 269172 34008 269178 34060
rect 143074 33940 143080 33992
rect 143132 33980 143138 33992
rect 276014 33980 276020 33992
rect 143132 33952 276020 33980
rect 143132 33940 143138 33952
rect 276014 33940 276020 33952
rect 276072 33940 276078 33992
rect 143626 33872 143632 33924
rect 143684 33912 143690 33924
rect 284386 33912 284392 33924
rect 143684 33884 284392 33912
rect 143684 33872 143690 33884
rect 284386 33872 284392 33884
rect 284444 33872 284450 33924
rect 144178 33804 144184 33856
rect 144236 33844 144242 33856
rect 291194 33844 291200 33856
rect 144236 33816 291200 33844
rect 144236 33804 144242 33816
rect 291194 33804 291200 33816
rect 291252 33804 291258 33856
rect 145006 33736 145012 33788
rect 145064 33776 145070 33788
rect 300854 33776 300860 33788
rect 145064 33748 300860 33776
rect 145064 33736 145070 33748
rect 300854 33736 300860 33748
rect 300912 33736 300918 33788
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 175274 33096 175280 33108
rect 2924 33068 175280 33096
rect 2924 33056 2930 33068
rect 175274 33056 175280 33068
rect 175332 33056 175338 33108
rect 135346 32920 135352 32972
rect 135404 32960 135410 32972
rect 176654 32960 176660 32972
rect 135404 32932 176660 32960
rect 135404 32920 135410 32932
rect 176654 32920 176660 32932
rect 176712 32920 176718 32972
rect 135622 32852 135628 32904
rect 135680 32892 135686 32904
rect 180794 32892 180800 32904
rect 135680 32864 180800 32892
rect 135680 32852 135686 32864
rect 180794 32852 180800 32864
rect 180852 32852 180858 32904
rect 135898 32784 135904 32836
rect 135956 32824 135962 32836
rect 184934 32824 184940 32836
rect 135956 32796 184940 32824
rect 135956 32784 135962 32796
rect 184934 32784 184940 32796
rect 184992 32784 184998 32836
rect 136726 32716 136732 32768
rect 136784 32756 136790 32768
rect 194594 32756 194600 32768
rect 136784 32728 194600 32756
rect 136784 32716 136790 32728
rect 194594 32716 194600 32728
rect 194652 32716 194658 32768
rect 137002 32648 137008 32700
rect 137060 32688 137066 32700
rect 198734 32688 198740 32700
rect 137060 32660 198740 32688
rect 137060 32648 137066 32660
rect 198734 32648 198740 32660
rect 198792 32648 198798 32700
rect 137554 32580 137560 32632
rect 137612 32620 137618 32632
rect 205634 32620 205640 32632
rect 137612 32592 205640 32620
rect 137612 32580 137618 32592
rect 205634 32580 205640 32592
rect 205692 32580 205698 32632
rect 142246 32512 142252 32564
rect 142304 32552 142310 32564
rect 266354 32552 266360 32564
rect 142304 32524 266360 32552
rect 142304 32512 142310 32524
rect 266354 32512 266360 32524
rect 266412 32512 266418 32564
rect 164326 32444 164332 32496
rect 164384 32484 164390 32496
rect 549254 32484 549260 32496
rect 164384 32456 549260 32484
rect 164384 32444 164390 32456
rect 549254 32444 549260 32456
rect 549312 32444 549318 32496
rect 166258 32376 166264 32428
rect 166316 32416 166322 32428
rect 574094 32416 574100 32428
rect 166316 32388 574100 32416
rect 166316 32376 166322 32388
rect 574094 32376 574100 32388
rect 574152 32376 574158 32428
rect 157610 31696 157616 31748
rect 157668 31736 157674 31748
rect 463694 31736 463700 31748
rect 157668 31708 463700 31736
rect 157668 31696 157674 31708
rect 463694 31696 463700 31708
rect 463752 31696 463758 31748
rect 158162 31628 158168 31680
rect 158220 31668 158226 31680
rect 470594 31668 470600 31680
rect 158220 31640 470600 31668
rect 158220 31628 158226 31640
rect 470594 31628 470600 31640
rect 470652 31628 470658 31680
rect 158714 31560 158720 31612
rect 158772 31600 158778 31612
rect 477494 31600 477500 31612
rect 158772 31572 477500 31600
rect 158772 31560 158778 31572
rect 477494 31560 477500 31572
rect 477552 31560 477558 31612
rect 159082 31492 159088 31544
rect 159140 31532 159146 31544
rect 481634 31532 481640 31544
rect 159140 31504 481640 31532
rect 159140 31492 159146 31504
rect 481634 31492 481640 31504
rect 481692 31492 481698 31544
rect 161106 31424 161112 31476
rect 161164 31464 161170 31476
rect 490006 31464 490012 31476
rect 161164 31436 490012 31464
rect 161164 31424 161170 31436
rect 490006 31424 490012 31436
rect 490064 31424 490070 31476
rect 160186 31356 160192 31408
rect 160244 31396 160250 31408
rect 496814 31396 496820 31408
rect 160244 31368 496820 31396
rect 160244 31356 160250 31368
rect 496814 31356 496820 31368
rect 496872 31356 496878 31408
rect 160738 31288 160744 31340
rect 160796 31328 160802 31340
rect 503714 31328 503720 31340
rect 160796 31300 503720 31328
rect 160796 31288 160802 31300
rect 503714 31288 503720 31300
rect 503772 31288 503778 31340
rect 162578 31220 162584 31272
rect 162636 31260 162642 31272
rect 510614 31260 510620 31272
rect 162636 31232 510620 31260
rect 162636 31220 162642 31232
rect 510614 31220 510620 31232
rect 510672 31220 510678 31272
rect 161842 31152 161848 31204
rect 161900 31192 161906 31204
rect 517514 31192 517520 31204
rect 161900 31164 517520 31192
rect 161900 31152 161906 31164
rect 517514 31152 517520 31164
rect 517572 31152 517578 31204
rect 166350 31084 166356 31136
rect 166408 31124 166414 31136
rect 524414 31124 524420 31136
rect 166408 31096 524420 31124
rect 166408 31084 166414 31096
rect 524414 31084 524420 31096
rect 524472 31084 524478 31136
rect 162118 31016 162124 31068
rect 162176 31056 162182 31068
rect 521654 31056 521660 31068
rect 162176 31028 521660 31056
rect 162176 31016 162182 31028
rect 521654 31016 521660 31028
rect 521712 31016 521718 31068
rect 154298 30268 154304 30320
rect 154356 30308 154362 30320
rect 307846 30308 307852 30320
rect 154356 30280 307852 30308
rect 154356 30268 154362 30280
rect 307846 30268 307852 30280
rect 307904 30268 307910 30320
rect 144914 30200 144920 30252
rect 144972 30240 144978 30252
rect 299474 30240 299480 30252
rect 144972 30212 299480 30240
rect 144972 30200 144978 30212
rect 299474 30200 299480 30212
rect 299532 30200 299538 30252
rect 145190 30132 145196 30184
rect 145248 30172 145254 30184
rect 303614 30172 303620 30184
rect 145248 30144 303620 30172
rect 145248 30132 145254 30144
rect 303614 30132 303620 30144
rect 303672 30132 303678 30184
rect 150710 30064 150716 30116
rect 150768 30104 150774 30116
rect 374086 30104 374092 30116
rect 150768 30076 374092 30104
rect 150768 30064 150774 30076
rect 374086 30064 374092 30076
rect 374144 30064 374150 30116
rect 154206 29996 154212 30048
rect 154264 30036 154270 30048
rect 382366 30036 382372 30048
rect 154264 30008 382372 30036
rect 154264 29996 154270 30008
rect 382366 29996 382372 30008
rect 382424 29996 382430 30048
rect 157242 29928 157248 29980
rect 157300 29968 157306 29980
rect 389174 29968 389180 29980
rect 157300 29940 389180 29968
rect 157300 29928 157306 29940
rect 389174 29928 389180 29940
rect 389232 29928 389238 29980
rect 155126 29860 155132 29912
rect 155184 29900 155190 29912
rect 431954 29900 431960 29912
rect 155184 29872 431960 29900
rect 155184 29860 155190 29872
rect 431954 29860 431960 29872
rect 432012 29860 432018 29912
rect 157058 29792 157064 29844
rect 157116 29832 157122 29844
rect 438854 29832 438860 29844
rect 157116 29804 438860 29832
rect 157116 29792 157122 29804
rect 438854 29792 438860 29804
rect 438912 29792 438918 29844
rect 155954 29724 155960 29776
rect 156012 29764 156018 29776
rect 441614 29764 441620 29776
rect 156012 29736 441620 29764
rect 156012 29724 156018 29736
rect 441614 29724 441620 29736
rect 441672 29724 441678 29776
rect 156230 29656 156236 29708
rect 156288 29696 156294 29708
rect 445754 29696 445760 29708
rect 156288 29668 445760 29696
rect 156288 29656 156294 29668
rect 445754 29656 445760 29668
rect 445812 29656 445818 29708
rect 156782 29588 156788 29640
rect 156840 29628 156846 29640
rect 452654 29628 452660 29640
rect 156840 29600 452660 29628
rect 156840 29588 156846 29600
rect 452654 29588 452660 29600
rect 452712 29588 452718 29640
rect 139394 28908 139400 28960
rect 139452 28948 139458 28960
rect 229094 28948 229100 28960
rect 139452 28920 229100 28948
rect 139452 28908 139458 28920
rect 229094 28908 229100 28920
rect 229152 28908 229158 28960
rect 151630 28840 151636 28892
rect 151688 28880 151694 28892
rect 242894 28880 242900 28892
rect 151688 28852 242900 28880
rect 151688 28840 151694 28852
rect 242894 28840 242900 28852
rect 242952 28840 242958 28892
rect 140222 28772 140228 28824
rect 140280 28812 140286 28824
rect 240134 28812 240140 28824
rect 140280 28784 240140 28812
rect 140280 28772 140286 28784
rect 240134 28772 240140 28784
rect 240192 28772 240198 28824
rect 140774 28704 140780 28756
rect 140832 28744 140838 28756
rect 247034 28744 247040 28756
rect 140832 28716 247040 28744
rect 140832 28704 140838 28716
rect 247034 28704 247040 28716
rect 247092 28704 247098 28756
rect 151538 28636 151544 28688
rect 151596 28676 151602 28688
rect 258074 28676 258080 28688
rect 151596 28648 258080 28676
rect 151596 28636 151602 28648
rect 258074 28636 258080 28648
rect 258132 28636 258138 28688
rect 141050 28568 141056 28620
rect 141108 28608 141114 28620
rect 251174 28608 251180 28620
rect 141108 28580 251180 28608
rect 141108 28568 141114 28580
rect 251174 28568 251180 28580
rect 251232 28568 251238 28620
rect 152826 28500 152832 28552
rect 152884 28540 152890 28552
rect 264974 28540 264980 28552
rect 152884 28512 264980 28540
rect 152884 28500 152890 28512
rect 264974 28500 264980 28512
rect 265032 28500 265038 28552
rect 153010 28432 153016 28484
rect 153068 28472 153074 28484
rect 271874 28472 271880 28484
rect 153068 28444 271880 28472
rect 153068 28432 153074 28444
rect 271874 28432 271880 28444
rect 271932 28432 271938 28484
rect 150434 28364 150440 28416
rect 150492 28404 150498 28416
rect 371234 28404 371240 28416
rect 150492 28376 371240 28404
rect 150492 28364 150498 28376
rect 371234 28364 371240 28376
rect 371292 28364 371298 28416
rect 152918 28296 152924 28348
rect 152976 28336 152982 28348
rect 375374 28336 375380 28348
rect 152976 28308 375380 28336
rect 152976 28296 152982 28308
rect 375374 28296 375380 28308
rect 375432 28296 375438 28348
rect 165982 28228 165988 28280
rect 166040 28268 166046 28280
rect 571334 28268 571340 28280
rect 166040 28240 571340 28268
rect 166040 28228 166046 28240
rect 571334 28228 571340 28240
rect 571392 28228 571398 28280
rect 138290 28160 138296 28212
rect 138348 28200 138354 28212
rect 215294 28200 215300 28212
rect 138348 28172 215300 28200
rect 138348 28160 138354 28172
rect 215294 28160 215300 28172
rect 215352 28160 215358 28212
rect 138106 28092 138112 28144
rect 138164 28132 138170 28144
rect 211154 28132 211160 28144
rect 138164 28104 211160 28132
rect 138164 28092 138170 28104
rect 211154 28092 211160 28104
rect 211212 28092 211218 28144
rect 150158 28024 150164 28076
rect 150216 28064 150222 28076
rect 222194 28064 222200 28076
rect 150216 28036 222200 28064
rect 150216 28024 150222 28036
rect 222194 28024 222200 28036
rect 222252 28024 222258 28076
rect 143166 27548 143172 27600
rect 143224 27588 143230 27600
rect 193214 27588 193220 27600
rect 143224 27560 193220 27588
rect 143224 27548 143230 27560
rect 193214 27548 193220 27560
rect 193272 27548 193278 27600
rect 136082 27480 136088 27532
rect 136140 27520 136146 27532
rect 186314 27520 186320 27532
rect 136140 27492 186320 27520
rect 136140 27480 136146 27492
rect 186314 27480 186320 27492
rect 186372 27480 186378 27532
rect 136910 27412 136916 27464
rect 136968 27452 136974 27464
rect 197354 27452 197360 27464
rect 136968 27424 197360 27452
rect 136968 27412 136974 27424
rect 197354 27412 197360 27424
rect 197412 27412 197418 27464
rect 146018 27344 146024 27396
rect 146076 27384 146082 27396
rect 208394 27384 208400 27396
rect 146076 27356 208400 27384
rect 146076 27344 146082 27356
rect 208394 27344 208400 27356
rect 208452 27344 208458 27396
rect 137186 27276 137192 27328
rect 137244 27316 137250 27328
rect 201494 27316 201500 27328
rect 137244 27288 201500 27316
rect 137244 27276 137250 27288
rect 201494 27276 201500 27288
rect 201552 27276 201558 27328
rect 137462 27208 137468 27260
rect 137520 27248 137526 27260
rect 204254 27248 204260 27260
rect 137520 27220 204260 27248
rect 137520 27208 137526 27220
rect 204254 27208 204260 27220
rect 204312 27208 204318 27260
rect 138566 27140 138572 27192
rect 138624 27180 138630 27192
rect 218054 27180 218060 27192
rect 138624 27152 218060 27180
rect 138624 27140 138630 27152
rect 218054 27140 218060 27152
rect 218112 27140 218118 27192
rect 139670 27072 139676 27124
rect 139728 27112 139734 27124
rect 233234 27112 233240 27124
rect 139728 27084 233240 27112
rect 139728 27072 139734 27084
rect 233234 27072 233240 27084
rect 233292 27072 233298 27124
rect 148318 27004 148324 27056
rect 148376 27044 148382 27056
rect 343634 27044 343640 27056
rect 148376 27016 343640 27044
rect 148376 27004 148382 27016
rect 343634 27004 343640 27016
rect 343692 27004 343698 27056
rect 154574 26936 154580 26988
rect 154632 26976 154638 26988
rect 423674 26976 423680 26988
rect 154632 26948 423680 26976
rect 154632 26936 154638 26948
rect 423674 26936 423680 26948
rect 423732 26936 423738 26988
rect 157978 26868 157984 26920
rect 158036 26908 158042 26920
rect 467834 26908 467840 26920
rect 158036 26880 467840 26908
rect 158036 26868 158042 26880
rect 467834 26868 467840 26880
rect 467892 26868 467898 26920
rect 135530 26188 135536 26240
rect 135588 26228 135594 26240
rect 179414 26228 179420 26240
rect 135588 26200 179420 26228
rect 135588 26188 135594 26200
rect 179414 26188 179420 26200
rect 179472 26188 179478 26240
rect 135806 26120 135812 26172
rect 135864 26160 135870 26172
rect 183554 26160 183560 26172
rect 135864 26132 183560 26160
rect 135864 26120 135870 26132
rect 183554 26120 183560 26132
rect 183612 26120 183618 26172
rect 139946 26052 139952 26104
rect 140004 26092 140010 26104
rect 235994 26092 236000 26104
rect 140004 26064 236000 26092
rect 140004 26052 140010 26064
rect 235994 26052 236000 26064
rect 236052 26052 236058 26104
rect 141878 25984 141884 26036
rect 141936 26024 141942 26036
rect 260834 26024 260840 26036
rect 141936 25996 260840 26024
rect 141936 25984 141942 25996
rect 260834 25984 260840 25996
rect 260892 25984 260898 26036
rect 144362 25916 144368 25968
rect 144420 25956 144426 25968
rect 292574 25956 292580 25968
rect 144420 25928 292580 25956
rect 144420 25916 144426 25928
rect 292574 25916 292580 25928
rect 292632 25916 292638 25968
rect 149330 25848 149336 25900
rect 149388 25888 149394 25900
rect 357526 25888 357532 25900
rect 149388 25860 357532 25888
rect 149388 25848 149394 25860
rect 357526 25848 357532 25860
rect 357584 25848 357590 25900
rect 150526 25780 150532 25832
rect 150584 25820 150590 25832
rect 372614 25820 372620 25832
rect 150584 25792 372620 25820
rect 150584 25780 150590 25792
rect 372614 25780 372620 25792
rect 372672 25780 372678 25832
rect 153746 25712 153752 25764
rect 153804 25752 153810 25764
rect 414014 25752 414020 25764
rect 153804 25724 414020 25752
rect 153804 25712 153810 25724
rect 414014 25712 414020 25724
rect 414072 25712 414078 25764
rect 164786 25644 164792 25696
rect 164844 25684 164850 25696
rect 556154 25684 556160 25696
rect 164844 25656 556160 25684
rect 164844 25644 164850 25656
rect 556154 25644 556160 25656
rect 556212 25644 556218 25696
rect 165614 25576 165620 25628
rect 165672 25616 165678 25628
rect 565814 25616 565820 25628
rect 165672 25588 565820 25616
rect 165672 25576 165678 25588
rect 565814 25576 565820 25588
rect 565872 25576 565878 25628
rect 81434 25508 81440 25560
rect 81492 25548 81498 25560
rect 120902 25548 120908 25560
rect 81492 25520 120908 25548
rect 81492 25508 81498 25520
rect 120902 25508 120908 25520
rect 120960 25508 120966 25560
rect 166166 25508 166172 25560
rect 166224 25548 166230 25560
rect 572714 25548 572720 25560
rect 166224 25520 572720 25548
rect 166224 25508 166230 25520
rect 572714 25508 572720 25520
rect 572772 25508 572778 25560
rect 135254 25440 135260 25492
rect 135312 25480 135318 25492
rect 176746 25480 176752 25492
rect 135312 25452 176752 25480
rect 135312 25440 135318 25452
rect 176746 25440 176752 25452
rect 176804 25440 176810 25492
rect 141326 24760 141332 24812
rect 141384 24800 141390 24812
rect 253934 24800 253940 24812
rect 141384 24772 253940 24800
rect 141384 24760 141390 24772
rect 253934 24760 253940 24772
rect 253992 24760 253998 24812
rect 143534 24692 143540 24744
rect 143592 24732 143598 24744
rect 282914 24732 282920 24744
rect 143592 24704 282920 24732
rect 143592 24692 143598 24704
rect 282914 24692 282920 24704
rect 282972 24692 282978 24744
rect 153194 24624 153200 24676
rect 153252 24664 153258 24676
rect 407206 24664 407212 24676
rect 153252 24636 407212 24664
rect 153252 24624 153258 24636
rect 407206 24624 407212 24636
rect 407264 24624 407270 24676
rect 162854 24556 162860 24608
rect 162912 24596 162918 24608
rect 531314 24596 531320 24608
rect 162912 24568 531320 24596
rect 162912 24556 162918 24568
rect 531314 24556 531320 24568
rect 531372 24556 531378 24608
rect 163130 24488 163136 24540
rect 163188 24528 163194 24540
rect 534074 24528 534080 24540
rect 163188 24500 534080 24528
rect 163188 24488 163194 24500
rect 534074 24488 534080 24500
rect 534132 24488 534138 24540
rect 163406 24420 163412 24472
rect 163464 24460 163470 24472
rect 538214 24460 538220 24472
rect 163464 24432 538220 24460
rect 163464 24420 163470 24432
rect 538214 24420 538220 24432
rect 538272 24420 538278 24472
rect 163682 24352 163688 24404
rect 163740 24392 163746 24404
rect 540974 24392 540980 24404
rect 163740 24364 540980 24392
rect 163740 24352 163746 24364
rect 540974 24352 540980 24364
rect 541032 24352 541038 24404
rect 164234 24284 164240 24336
rect 164292 24324 164298 24336
rect 547874 24324 547880 24336
rect 164292 24296 547880 24324
rect 164292 24284 164298 24296
rect 547874 24284 547880 24296
rect 547932 24284 547938 24336
rect 164510 24216 164516 24268
rect 164568 24256 164574 24268
rect 552014 24256 552020 24268
rect 164568 24228 552020 24256
rect 164568 24216 164574 24228
rect 552014 24216 552020 24228
rect 552072 24216 552078 24268
rect 165706 24148 165712 24200
rect 165764 24188 165770 24200
rect 567194 24188 567200 24200
rect 165764 24160 567200 24188
rect 165764 24148 165770 24160
rect 567194 24148 567200 24160
rect 567252 24148 567258 24200
rect 165890 24080 165896 24132
rect 165948 24120 165954 24132
rect 569954 24120 569960 24132
rect 165948 24092 569960 24120
rect 165948 24080 165954 24092
rect 569954 24080 569960 24092
rect 570012 24080 570018 24132
rect 157334 23400 157340 23452
rect 157392 23440 157398 23452
rect 459554 23440 459560 23452
rect 157392 23412 459560 23440
rect 157392 23400 157398 23412
rect 459554 23400 459560 23412
rect 459612 23400 459618 23452
rect 160094 23332 160100 23384
rect 160152 23372 160158 23384
rect 495434 23372 495440 23384
rect 160152 23344 495440 23372
rect 160152 23332 160158 23344
rect 495434 23332 495440 23344
rect 495492 23332 495498 23384
rect 160370 23264 160376 23316
rect 160428 23304 160434 23316
rect 498286 23304 498292 23316
rect 160428 23276 498292 23304
rect 160428 23264 160434 23276
rect 498286 23264 498292 23276
rect 498344 23264 498350 23316
rect 160646 23196 160652 23248
rect 160704 23236 160710 23248
rect 502334 23236 502340 23248
rect 160704 23208 502340 23236
rect 160704 23196 160710 23208
rect 502334 23196 502340 23208
rect 502392 23196 502398 23248
rect 160922 23128 160928 23180
rect 160980 23168 160986 23180
rect 506474 23168 506480 23180
rect 160980 23140 506480 23168
rect 160980 23128 160986 23140
rect 506474 23128 506480 23140
rect 506532 23128 506538 23180
rect 161474 23060 161480 23112
rect 161532 23100 161538 23112
rect 513374 23100 513380 23112
rect 161532 23072 513380 23100
rect 161532 23060 161538 23072
rect 513374 23060 513380 23072
rect 513432 23060 513438 23112
rect 161750 22992 161756 23044
rect 161808 23032 161814 23044
rect 516134 23032 516140 23044
rect 161808 23004 516140 23032
rect 161808 22992 161814 23004
rect 516134 22992 516140 23004
rect 516192 22992 516198 23044
rect 162026 22924 162032 22976
rect 162084 22964 162090 22976
rect 520274 22964 520280 22976
rect 162084 22936 520280 22964
rect 162084 22924 162090 22936
rect 520274 22924 520280 22936
rect 520332 22924 520338 22976
rect 162302 22856 162308 22908
rect 162360 22896 162366 22908
rect 523034 22896 523040 22908
rect 162360 22868 523040 22896
rect 162360 22856 162366 22868
rect 523034 22856 523040 22868
rect 523092 22856 523098 22908
rect 165154 22788 165160 22840
rect 165212 22828 165218 22840
rect 560294 22828 560300 22840
rect 165212 22800 560300 22828
rect 165212 22788 165218 22800
rect 560294 22788 560300 22800
rect 560352 22788 560358 22840
rect 114462 22720 114468 22772
rect 114520 22760 114526 22772
rect 580166 22760 580172 22772
rect 114520 22732 580172 22760
rect 114520 22720 114526 22732
rect 580166 22720 580172 22732
rect 580224 22720 580230 22772
rect 3510 22652 3516 22704
rect 3568 22692 3574 22704
rect 170306 22692 170312 22704
rect 3568 22664 170312 22692
rect 3568 22652 3574 22664
rect 170306 22652 170312 22664
rect 170364 22652 170370 22704
rect 148042 22040 148048 22092
rect 148100 22080 148106 22092
rect 340874 22080 340880 22092
rect 148100 22052 340880 22080
rect 148100 22040 148106 22052
rect 340874 22040 340880 22052
rect 340932 22040 340938 22092
rect 156966 21972 156972 22024
rect 157024 22012 157030 22024
rect 361574 22012 361580 22024
rect 157024 21984 361580 22012
rect 157024 21972 157030 21984
rect 361574 21972 361580 21984
rect 361632 21972 361638 22024
rect 154666 21904 154672 21956
rect 154724 21944 154730 21956
rect 425054 21944 425060 21956
rect 154724 21916 425060 21944
rect 154724 21904 154730 21916
rect 425054 21904 425060 21916
rect 425112 21904 425118 21956
rect 155034 21836 155040 21888
rect 155092 21876 155098 21888
rect 430574 21876 430580 21888
rect 155092 21848 430580 21876
rect 155092 21836 155098 21848
rect 430574 21836 430580 21848
rect 430632 21836 430638 21888
rect 155218 21768 155224 21820
rect 155276 21808 155282 21820
rect 432046 21808 432052 21820
rect 155276 21780 432052 21808
rect 155276 21768 155282 21780
rect 432046 21768 432052 21780
rect 432104 21768 432110 21820
rect 156322 21700 156328 21752
rect 156380 21740 156386 21752
rect 447134 21740 447140 21752
rect 156380 21712 447140 21740
rect 156380 21700 156386 21712
rect 447134 21700 447140 21712
rect 447192 21700 447198 21752
rect 156414 21632 156420 21684
rect 156472 21672 156478 21684
rect 448514 21672 448520 21684
rect 156472 21644 448520 21672
rect 156472 21632 156478 21644
rect 448514 21632 448520 21644
rect 448572 21632 448578 21684
rect 158990 21564 158996 21616
rect 159048 21604 159054 21616
rect 481726 21604 481732 21616
rect 159048 21576 481732 21604
rect 159048 21564 159054 21576
rect 481726 21564 481732 21576
rect 481784 21564 481790 21616
rect 159266 21496 159272 21548
rect 159324 21536 159330 21548
rect 484394 21536 484400 21548
rect 159324 21508 484400 21536
rect 159324 21496 159330 21508
rect 484394 21496 484400 21508
rect 484452 21496 484458 21548
rect 159542 21428 159548 21480
rect 159600 21468 159606 21480
rect 488534 21468 488540 21480
rect 159600 21440 488540 21468
rect 159600 21428 159606 21440
rect 488534 21428 488540 21440
rect 488592 21428 488598 21480
rect 159818 21360 159824 21412
rect 159876 21400 159882 21412
rect 491294 21400 491300 21412
rect 159876 21372 491300 21400
rect 159876 21360 159882 21372
rect 491294 21360 491300 21372
rect 491352 21360 491358 21412
rect 139486 20408 139492 20460
rect 139544 20448 139550 20460
rect 230474 20448 230480 20460
rect 139544 20420 230480 20448
rect 139544 20408 139550 20420
rect 230474 20408 230480 20420
rect 230532 20408 230538 20460
rect 140038 20340 140044 20392
rect 140096 20380 140102 20392
rect 237374 20380 237380 20392
rect 140096 20352 237380 20380
rect 140096 20340 140102 20352
rect 237374 20340 237380 20352
rect 237432 20340 237438 20392
rect 141694 20272 141700 20324
rect 141752 20312 141758 20324
rect 259546 20312 259552 20324
rect 141752 20284 259552 20312
rect 141752 20272 141758 20284
rect 259546 20272 259552 20284
rect 259604 20272 259610 20324
rect 147214 20204 147220 20256
rect 147272 20244 147278 20256
rect 329834 20244 329840 20256
rect 147272 20216 329840 20244
rect 147272 20204 147278 20216
rect 329834 20204 329840 20216
rect 329892 20204 329898 20256
rect 152274 20136 152280 20188
rect 152332 20176 152338 20188
rect 394694 20176 394700 20188
rect 152332 20148 394700 20176
rect 152332 20136 152338 20148
rect 394694 20136 394700 20148
rect 394752 20136 394758 20188
rect 152550 20068 152556 20120
rect 152608 20108 152614 20120
rect 398834 20108 398840 20120
rect 152608 20080 398840 20108
rect 152608 20068 152614 20080
rect 398834 20068 398840 20080
rect 398892 20068 398898 20120
rect 153654 20000 153660 20052
rect 153712 20040 153718 20052
rect 412634 20040 412640 20052
rect 153712 20012 412640 20040
rect 153712 20000 153718 20012
rect 412634 20000 412640 20012
rect 412692 20000 412698 20052
rect 158070 19932 158076 19984
rect 158128 19972 158134 19984
rect 469214 19972 469220 19984
rect 158128 19944 469220 19972
rect 158128 19932 158134 19944
rect 469214 19932 469220 19944
rect 469272 19932 469278 19984
rect 141142 19048 141148 19100
rect 141200 19088 141206 19100
rect 251266 19088 251272 19100
rect 141200 19060 251272 19088
rect 141200 19048 141206 19060
rect 251266 19048 251272 19060
rect 251324 19048 251330 19100
rect 163774 18980 163780 19032
rect 163832 19020 163838 19032
rect 312538 19020 312544 19032
rect 163832 18992 312544 19020
rect 163832 18980 163838 18992
rect 312538 18980 312544 18992
rect 312596 18980 312602 19032
rect 149514 18912 149520 18964
rect 149572 18952 149578 18964
rect 358814 18952 358820 18964
rect 149572 18924 358820 18952
rect 149572 18912 149578 18924
rect 358814 18912 358820 18924
rect 358872 18912 358878 18964
rect 150894 18844 150900 18896
rect 150952 18884 150958 18896
rect 376754 18884 376760 18896
rect 150952 18856 376760 18884
rect 150952 18844 150958 18856
rect 376754 18844 376760 18856
rect 376812 18844 376818 18896
rect 151170 18776 151176 18828
rect 151228 18816 151234 18828
rect 380894 18816 380900 18828
rect 151228 18788 380900 18816
rect 151228 18776 151234 18788
rect 380894 18776 380900 18788
rect 380952 18776 380958 18828
rect 156690 18708 156696 18760
rect 156748 18748 156754 18760
rect 451274 18748 451280 18760
rect 156748 18720 451280 18748
rect 156748 18708 156754 18720
rect 451274 18708 451280 18720
rect 451332 18708 451338 18760
rect 163222 18640 163228 18692
rect 163280 18680 163286 18692
rect 535454 18680 535460 18692
rect 163280 18652 535460 18680
rect 163280 18640 163286 18652
rect 535454 18640 535460 18652
rect 535512 18640 535518 18692
rect 35894 18572 35900 18624
rect 35952 18612 35958 18624
rect 118142 18612 118148 18624
rect 35952 18584 118148 18612
rect 35952 18572 35958 18584
rect 118142 18572 118148 18584
rect 118200 18572 118206 18624
rect 164602 18572 164608 18624
rect 164660 18612 164666 18624
rect 553394 18612 553400 18624
rect 164660 18584 553400 18612
rect 164660 18572 164666 18584
rect 553394 18572 553400 18584
rect 553452 18572 553458 18624
rect 142798 17620 142804 17672
rect 142856 17660 142862 17672
rect 273254 17660 273260 17672
rect 142856 17632 273260 17660
rect 142856 17620 142862 17632
rect 273254 17620 273260 17632
rect 273312 17620 273318 17672
rect 147030 17552 147036 17604
rect 147088 17592 147094 17604
rect 327074 17592 327080 17604
rect 147088 17564 327080 17592
rect 147088 17552 147094 17564
rect 327074 17552 327080 17564
rect 327132 17552 327138 17604
rect 154850 17484 154856 17536
rect 154908 17524 154914 17536
rect 427814 17524 427820 17536
rect 154908 17496 427820 17524
rect 154908 17484 154914 17496
rect 427814 17484 427820 17496
rect 427872 17484 427878 17536
rect 155310 17416 155316 17468
rect 155368 17456 155374 17468
rect 433334 17456 433340 17468
rect 155368 17428 433340 17456
rect 155368 17416 155374 17428
rect 433334 17416 433340 17428
rect 433392 17416 433398 17468
rect 155402 17348 155408 17400
rect 155460 17388 155466 17400
rect 434714 17388 434720 17400
rect 155460 17360 434720 17388
rect 155460 17348 155466 17360
rect 434714 17348 434720 17360
rect 434772 17348 434778 17400
rect 155586 17280 155592 17332
rect 155644 17320 155650 17332
rect 437474 17320 437480 17332
rect 155644 17292 437480 17320
rect 155644 17280 155650 17292
rect 437474 17280 437480 17292
rect 437532 17280 437538 17332
rect 164878 17212 164884 17264
rect 164936 17252 164942 17264
rect 556246 17252 556252 17264
rect 164936 17224 556252 17252
rect 164936 17212 164942 17224
rect 556246 17212 556252 17224
rect 556304 17212 556310 17264
rect 142890 16328 142896 16380
rect 142948 16368 142954 16380
rect 274818 16368 274824 16380
rect 142948 16340 274824 16368
rect 142948 16328 142954 16340
rect 274818 16328 274824 16340
rect 274876 16328 274882 16380
rect 143902 16260 143908 16312
rect 143960 16300 143966 16312
rect 287330 16300 287336 16312
rect 143960 16272 287336 16300
rect 143960 16260 143966 16272
rect 287330 16260 287336 16272
rect 287388 16260 287394 16312
rect 143994 16192 144000 16244
rect 144052 16232 144058 16244
rect 288986 16232 288992 16244
rect 144052 16204 288992 16232
rect 144052 16192 144058 16204
rect 288986 16192 288992 16204
rect 289044 16192 289050 16244
rect 144270 16124 144276 16176
rect 144328 16164 144334 16176
rect 292666 16164 292672 16176
rect 144328 16136 292672 16164
rect 144328 16124 144334 16136
rect 292666 16124 292672 16136
rect 292724 16124 292730 16176
rect 148502 16056 148508 16108
rect 148560 16096 148566 16108
rect 346946 16096 346952 16108
rect 148560 16068 346952 16096
rect 148560 16056 148566 16068
rect 346946 16056 346952 16068
rect 347004 16056 347010 16108
rect 149054 15988 149060 16040
rect 149112 16028 149118 16040
rect 353570 16028 353576 16040
rect 149112 16000 353576 16028
rect 149112 15988 149118 16000
rect 353570 15988 353576 16000
rect 353628 15988 353634 16040
rect 153930 15920 153936 15972
rect 153988 15960 153994 15972
rect 415486 15960 415492 15972
rect 153988 15932 415492 15960
rect 153988 15920 153994 15932
rect 415486 15920 415492 15932
rect 415544 15920 415550 15972
rect 162946 15852 162952 15904
rect 163004 15892 163010 15904
rect 532050 15892 532056 15904
rect 163004 15864 532056 15892
rect 163004 15852 163010 15864
rect 532050 15852 532056 15864
rect 532108 15852 532114 15904
rect 141234 14832 141240 14884
rect 141292 14872 141298 14884
rect 253474 14872 253480 14884
rect 141292 14844 253480 14872
rect 141292 14832 141298 14844
rect 253474 14832 253480 14844
rect 253532 14832 253538 14884
rect 141510 14764 141516 14816
rect 141568 14804 141574 14816
rect 256694 14804 256700 14816
rect 141568 14776 256700 14804
rect 141568 14764 141574 14776
rect 256694 14764 256700 14776
rect 256752 14764 256758 14816
rect 142338 14696 142344 14748
rect 142396 14736 142402 14748
rect 267734 14736 267740 14748
rect 142396 14708 267740 14736
rect 142396 14696 142402 14708
rect 267734 14696 267740 14708
rect 267792 14696 267798 14748
rect 142614 14628 142620 14680
rect 142672 14668 142678 14680
rect 270770 14668 270776 14680
rect 142672 14640 270776 14668
rect 142672 14628 142678 14640
rect 270770 14628 270776 14640
rect 270828 14628 270834 14680
rect 149606 14560 149612 14612
rect 149664 14600 149670 14612
rect 361114 14600 361120 14612
rect 149664 14572 361120 14600
rect 149664 14560 149670 14572
rect 361114 14560 361120 14572
rect 361172 14560 361178 14612
rect 151446 14492 151452 14544
rect 151504 14532 151510 14544
rect 384298 14532 384304 14544
rect 151504 14504 384304 14532
rect 151504 14492 151510 14504
rect 384298 14492 384304 14504
rect 384356 14492 384362 14544
rect 157886 14424 157892 14476
rect 157944 14464 157950 14476
rect 467466 14464 467472 14476
rect 157944 14436 467472 14464
rect 157944 14424 157950 14436
rect 467466 14424 467472 14436
rect 467524 14424 467530 14476
rect 139578 13404 139584 13456
rect 139636 13444 139642 13456
rect 231854 13444 231860 13456
rect 139636 13416 231860 13444
rect 139636 13404 139642 13416
rect 231854 13404 231860 13416
rect 231912 13404 231918 13456
rect 140130 13336 140136 13388
rect 140188 13376 140194 13388
rect 239306 13376 239312 13388
rect 140188 13348 239312 13376
rect 140188 13336 140194 13348
rect 239306 13336 239312 13348
rect 239364 13336 239370 13388
rect 146846 13268 146852 13320
rect 146904 13308 146910 13320
rect 324406 13308 324412 13320
rect 146904 13280 324412 13308
rect 146904 13268 146910 13280
rect 324406 13268 324412 13280
rect 324464 13268 324470 13320
rect 147122 13200 147128 13252
rect 147180 13240 147186 13252
rect 328730 13240 328736 13252
rect 147180 13212 328736 13240
rect 147180 13200 147186 13212
rect 328730 13200 328736 13212
rect 328788 13200 328794 13252
rect 149790 13132 149796 13184
rect 149848 13172 149854 13184
rect 363506 13172 363512 13184
rect 149848 13144 363512 13172
rect 149848 13132 149854 13144
rect 363506 13132 363512 13144
rect 363564 13132 363570 13184
rect 14274 13064 14280 13116
rect 14332 13104 14338 13116
rect 122098 13104 122104 13116
rect 14332 13076 122104 13104
rect 14332 13064 14338 13076
rect 122098 13064 122104 13076
rect 122156 13064 122162 13116
rect 150986 13064 150992 13116
rect 151044 13104 151050 13116
rect 378410 13104 378416 13116
rect 151044 13076 378416 13104
rect 151044 13064 151050 13076
rect 378410 13064 378416 13076
rect 378468 13064 378474 13116
rect 157702 12248 157708 12300
rect 157760 12288 157766 12300
rect 169018 12288 169024 12300
rect 157760 12260 169024 12288
rect 157760 12248 157766 12260
rect 169018 12248 169024 12260
rect 169076 12248 169082 12300
rect 138198 12180 138204 12232
rect 138256 12220 138262 12232
rect 214466 12220 214472 12232
rect 138256 12192 214472 12220
rect 138256 12180 138262 12192
rect 214466 12180 214472 12192
rect 214524 12180 214530 12232
rect 138474 12112 138480 12164
rect 138532 12152 138538 12164
rect 218146 12152 218152 12164
rect 138532 12124 218152 12152
rect 138532 12112 138538 12124
rect 218146 12112 218152 12124
rect 218204 12112 218210 12164
rect 138750 12044 138756 12096
rect 138808 12084 138814 12096
rect 221090 12084 221096 12096
rect 138808 12056 221096 12084
rect 138808 12044 138814 12056
rect 221090 12044 221096 12056
rect 221148 12044 221154 12096
rect 146570 11976 146576 12028
rect 146628 12016 146634 12028
rect 322106 12016 322112 12028
rect 146628 11988 322112 12016
rect 146628 11976 146634 11988
rect 322106 11976 322112 11988
rect 322164 11976 322170 12028
rect 148226 11908 148232 11960
rect 148284 11948 148290 11960
rect 342898 11948 342904 11960
rect 148284 11920 342904 11948
rect 148284 11908 148290 11920
rect 342898 11908 342904 11920
rect 342956 11908 342962 11960
rect 131390 11840 131396 11892
rect 131448 11840 131454 11892
rect 148410 11840 148416 11892
rect 148468 11880 148474 11892
rect 345290 11880 345296 11892
rect 148468 11852 345296 11880
rect 148468 11840 148474 11852
rect 345290 11840 345296 11852
rect 345348 11840 345354 11892
rect 131114 11636 131120 11688
rect 131172 11676 131178 11688
rect 131298 11676 131304 11688
rect 131172 11648 131304 11676
rect 131172 11636 131178 11648
rect 131298 11636 131304 11648
rect 131356 11636 131362 11688
rect 131114 11500 131120 11552
rect 131172 11540 131178 11552
rect 131408 11540 131436 11840
rect 149238 11772 149244 11824
rect 149296 11812 149302 11824
rect 356330 11812 356336 11824
rect 149296 11784 356336 11812
rect 149296 11772 149302 11784
rect 356330 11772 356336 11784
rect 356388 11772 356394 11824
rect 159358 11704 159364 11756
rect 159416 11744 159422 11756
rect 486418 11744 486424 11756
rect 159416 11716 486424 11744
rect 159416 11704 159422 11716
rect 486418 11704 486424 11716
rect 486476 11704 486482 11756
rect 176654 11636 176660 11688
rect 176712 11676 176718 11688
rect 177850 11676 177856 11688
rect 176712 11648 177856 11676
rect 176712 11636 176718 11648
rect 177850 11636 177856 11648
rect 177908 11636 177914 11688
rect 218054 11636 218060 11688
rect 218112 11676 218118 11688
rect 219250 11676 219256 11688
rect 218112 11648 219256 11676
rect 218112 11636 218118 11648
rect 219250 11636 219256 11648
rect 219308 11636 219314 11688
rect 242894 11636 242900 11688
rect 242952 11676 242958 11688
rect 244090 11676 244096 11688
rect 242952 11648 244096 11676
rect 242952 11636 242958 11648
rect 244090 11636 244096 11648
rect 244148 11636 244154 11688
rect 259454 11636 259460 11688
rect 259512 11676 259518 11688
rect 260650 11676 260656 11688
rect 259512 11648 260656 11676
rect 259512 11636 259518 11648
rect 260650 11636 260656 11648
rect 260708 11636 260714 11688
rect 131172 11512 131436 11540
rect 131172 11500 131178 11512
rect 110506 10956 110512 11008
rect 110564 10996 110570 11008
rect 130378 10996 130384 11008
rect 110564 10968 130384 10996
rect 110564 10956 110570 10968
rect 130378 10956 130384 10968
rect 130436 10956 130442 11008
rect 102134 10888 102140 10940
rect 102192 10928 102198 10940
rect 129090 10928 129096 10940
rect 102192 10900 129096 10928
rect 102192 10888 102198 10900
rect 129090 10888 129096 10900
rect 129148 10888 129154 10940
rect 95786 10820 95792 10872
rect 95844 10860 95850 10872
rect 128998 10860 129004 10872
rect 95844 10832 129004 10860
rect 95844 10820 95850 10832
rect 128998 10820 129004 10832
rect 129056 10820 129062 10872
rect 134794 10820 134800 10872
rect 134852 10860 134858 10872
rect 170306 10860 170312 10872
rect 134852 10832 170312 10860
rect 134852 10820 134858 10832
rect 170306 10820 170312 10832
rect 170364 10820 170370 10872
rect 92474 10752 92480 10804
rect 92532 10792 92538 10804
rect 129182 10792 129188 10804
rect 92532 10764 129188 10792
rect 92532 10752 92538 10764
rect 129182 10752 129188 10764
rect 129240 10752 129246 10804
rect 137094 10752 137100 10804
rect 137152 10792 137158 10804
rect 200298 10792 200304 10804
rect 137152 10764 200304 10792
rect 137152 10752 137158 10764
rect 200298 10752 200304 10764
rect 200356 10752 200362 10804
rect 74994 10684 75000 10736
rect 75052 10724 75058 10736
rect 122190 10724 122196 10736
rect 75052 10696 122196 10724
rect 75052 10684 75058 10696
rect 122190 10684 122196 10696
rect 122248 10684 122254 10736
rect 137370 10684 137376 10736
rect 137428 10724 137434 10736
rect 203426 10724 203432 10736
rect 137428 10696 203432 10724
rect 137428 10684 137434 10696
rect 203426 10684 203432 10696
rect 203484 10684 203490 10736
rect 78122 10616 78128 10668
rect 78180 10656 78186 10668
rect 127802 10656 127808 10668
rect 78180 10628 127808 10656
rect 78180 10616 78186 10628
rect 127802 10616 127808 10628
rect 127860 10616 127866 10668
rect 142982 10616 142988 10668
rect 143040 10656 143046 10668
rect 276106 10656 276112 10668
rect 143040 10628 276112 10656
rect 143040 10616 143046 10628
rect 276106 10616 276112 10628
rect 276164 10616 276170 10668
rect 67634 10548 67640 10600
rect 67692 10588 67698 10600
rect 126422 10588 126428 10600
rect 67692 10560 126428 10588
rect 67692 10548 67698 10560
rect 126422 10548 126428 10560
rect 126480 10548 126486 10600
rect 144454 10548 144460 10600
rect 144512 10588 144518 10600
rect 294874 10588 294880 10600
rect 144512 10560 294880 10588
rect 144512 10548 144518 10560
rect 294874 10548 294880 10560
rect 294932 10548 294938 10600
rect 64322 10480 64328 10532
rect 64380 10520 64386 10532
rect 126330 10520 126336 10532
rect 64380 10492 126336 10520
rect 64380 10480 64386 10492
rect 126330 10480 126336 10492
rect 126388 10480 126394 10532
rect 145926 10480 145932 10532
rect 145984 10520 145990 10532
rect 313826 10520 313832 10532
rect 145984 10492 313832 10520
rect 145984 10480 145990 10492
rect 313826 10480 313832 10492
rect 313884 10480 313890 10532
rect 46658 10412 46664 10464
rect 46716 10452 46722 10464
rect 125042 10452 125048 10464
rect 46716 10424 125048 10452
rect 46716 10412 46722 10424
rect 125042 10412 125048 10424
rect 125100 10412 125106 10464
rect 146294 10412 146300 10464
rect 146352 10452 146358 10464
rect 318058 10452 318064 10464
rect 146352 10424 318064 10452
rect 146352 10412 146358 10424
rect 318058 10412 318064 10424
rect 318116 10412 318122 10464
rect 31938 10344 31944 10396
rect 31996 10384 32002 10396
rect 123662 10384 123668 10396
rect 31996 10356 123668 10384
rect 31996 10344 32002 10356
rect 123662 10344 123668 10356
rect 123720 10344 123726 10396
rect 152642 10344 152648 10396
rect 152700 10384 152706 10396
rect 398926 10384 398932 10396
rect 152700 10356 398932 10384
rect 152700 10344 152706 10356
rect 398926 10344 398932 10356
rect 398984 10344 398990 10396
rect 25314 10276 25320 10328
rect 25372 10316 25378 10328
rect 123570 10316 123576 10328
rect 25372 10288 123576 10316
rect 25372 10276 25378 10288
rect 123570 10276 123576 10288
rect 123628 10276 123634 10328
rect 156506 10276 156512 10328
rect 156564 10316 156570 10328
rect 448606 10316 448612 10328
rect 156564 10288 448612 10316
rect 156564 10276 156570 10288
rect 448606 10276 448612 10288
rect 448664 10276 448670 10328
rect 117314 10208 117320 10260
rect 117372 10248 117378 10260
rect 130562 10248 130568 10260
rect 117372 10220 130568 10248
rect 117372 10208 117378 10220
rect 130562 10208 130568 10220
rect 130620 10208 130626 10260
rect 120626 10140 120632 10192
rect 120684 10180 120690 10192
rect 130470 10180 130476 10192
rect 120684 10152 130476 10180
rect 120684 10140 120690 10152
rect 130470 10140 130476 10152
rect 130528 10140 130534 10192
rect 116394 9596 116400 9648
rect 116452 9636 116458 9648
rect 130194 9636 130200 9648
rect 116452 9608 130200 9636
rect 116452 9596 116458 9608
rect 130194 9596 130200 9608
rect 130252 9596 130258 9648
rect 134886 9596 134892 9648
rect 134944 9636 134950 9648
rect 171962 9636 171968 9648
rect 134944 9608 171968 9636
rect 134944 9596 134950 9608
rect 171962 9596 171968 9608
rect 172020 9596 172026 9648
rect 112806 9528 112812 9580
rect 112864 9568 112870 9580
rect 130286 9568 130292 9580
rect 112864 9540 130292 9568
rect 112864 9528 112870 9540
rect 130286 9528 130292 9540
rect 130344 9528 130350 9580
rect 135438 9528 135444 9580
rect 135496 9568 135502 9580
rect 179046 9568 179052 9580
rect 135496 9540 179052 9568
rect 135496 9528 135502 9540
rect 179046 9528 179052 9540
rect 179104 9528 179110 9580
rect 60826 9460 60832 9512
rect 60884 9500 60890 9512
rect 126146 9500 126152 9512
rect 60884 9472 126152 9500
rect 60884 9460 60890 9472
rect 126146 9460 126152 9472
rect 126204 9460 126210 9512
rect 135990 9460 135996 9512
rect 136048 9500 136054 9512
rect 186130 9500 186136 9512
rect 136048 9472 186136 9500
rect 136048 9460 136054 9472
rect 186130 9460 186136 9472
rect 186188 9460 186194 9512
rect 57238 9392 57244 9444
rect 57296 9432 57302 9444
rect 126238 9432 126244 9444
rect 57296 9404 126244 9432
rect 57296 9392 57302 9404
rect 126238 9392 126244 9404
rect 126296 9392 126302 9444
rect 145374 9392 145380 9444
rect 145432 9432 145438 9444
rect 306742 9432 306748 9444
rect 145432 9404 306748 9432
rect 145432 9392 145438 9404
rect 306742 9392 306748 9404
rect 306800 9392 306806 9444
rect 43070 9324 43076 9376
rect 43128 9364 43134 9376
rect 116578 9364 116584 9376
rect 43128 9336 116584 9364
rect 43128 9324 43134 9336
rect 116578 9324 116584 9336
rect 116636 9324 116642 9376
rect 145650 9324 145656 9376
rect 145708 9364 145714 9376
rect 310238 9364 310244 9376
rect 145708 9336 310244 9364
rect 145708 9324 145714 9336
rect 310238 9324 310244 9336
rect 310296 9324 310302 9376
rect 50154 9256 50160 9308
rect 50212 9296 50218 9308
rect 124858 9296 124864 9308
rect 50212 9268 124864 9296
rect 50212 9256 50218 9268
rect 124858 9256 124864 9268
rect 124916 9256 124922 9308
rect 145742 9256 145748 9308
rect 145800 9296 145806 9308
rect 311434 9296 311440 9308
rect 145800 9268 311440 9296
rect 145800 9256 145806 9268
rect 311434 9256 311440 9268
rect 311492 9256 311498 9308
rect 45462 9188 45468 9240
rect 45520 9228 45526 9240
rect 124766 9228 124772 9240
rect 45520 9200 124772 9228
rect 45520 9188 45526 9200
rect 124766 9188 124772 9200
rect 124824 9188 124830 9240
rect 147950 9188 147956 9240
rect 148008 9228 148014 9240
rect 339862 9228 339868 9240
rect 148008 9200 339868 9228
rect 148008 9188 148014 9200
rect 339862 9188 339868 9200
rect 339920 9188 339926 9240
rect 41874 9120 41880 9172
rect 41932 9160 41938 9172
rect 124950 9160 124956 9172
rect 41932 9132 124956 9160
rect 41932 9120 41938 9132
rect 124950 9120 124956 9132
rect 125008 9120 125014 9172
rect 148134 9120 148140 9172
rect 148192 9160 148198 9172
rect 342162 9160 342168 9172
rect 148192 9132 342168 9160
rect 148192 9120 148198 9132
rect 342162 9120 342168 9132
rect 342220 9120 342226 9172
rect 31294 9052 31300 9104
rect 31352 9092 31358 9104
rect 123478 9092 123484 9104
rect 31352 9064 123484 9092
rect 31352 9052 31358 9064
rect 123478 9052 123484 9064
rect 123536 9052 123542 9104
rect 152090 9052 152096 9104
rect 152148 9092 152154 9104
rect 393038 9092 393044 9104
rect 152148 9064 393044 9092
rect 152148 9052 152154 9064
rect 393038 9052 393044 9064
rect 393096 9052 393102 9104
rect 24210 8984 24216 9036
rect 24268 9024 24274 9036
rect 123386 9024 123392 9036
rect 24268 8996 123392 9024
rect 24268 8984 24274 8996
rect 123386 8984 123392 8996
rect 123444 8984 123450 9036
rect 153470 8984 153476 9036
rect 153528 9024 153534 9036
rect 410794 9024 410800 9036
rect 153528 8996 410800 9024
rect 153528 8984 153534 8996
rect 410794 8984 410800 8996
rect 410852 8984 410858 9036
rect 9950 8916 9956 8968
rect 10008 8956 10014 8968
rect 122006 8956 122012 8968
rect 10008 8928 122012 8956
rect 10008 8916 10014 8928
rect 122006 8916 122012 8928
rect 122064 8916 122070 8968
rect 153562 8916 153568 8968
rect 153620 8956 153626 8968
rect 411898 8956 411904 8968
rect 153620 8928 411904 8956
rect 153620 8916 153626 8928
rect 411898 8916 411904 8928
rect 411956 8916 411962 8968
rect 98638 8236 98644 8288
rect 98696 8276 98702 8288
rect 128906 8276 128912 8288
rect 98696 8248 128912 8276
rect 98696 8236 98702 8248
rect 128906 8236 128912 8248
rect 128964 8236 128970 8288
rect 481634 8236 481640 8288
rect 481692 8276 481698 8288
rect 482462 8276 482468 8288
rect 481692 8248 482468 8276
rect 481692 8236 481698 8248
rect 482462 8236 482468 8248
rect 482520 8236 482526 8288
rect 95142 8168 95148 8220
rect 95200 8208 95206 8220
rect 128722 8208 128728 8220
rect 95200 8180 128728 8208
rect 95200 8168 95206 8180
rect 128722 8168 128728 8180
rect 128780 8168 128786 8220
rect 84470 8100 84476 8152
rect 84528 8140 84534 8152
rect 127710 8140 127716 8152
rect 84528 8112 127716 8140
rect 84528 8100 84534 8112
rect 127710 8100 127716 8112
rect 127768 8100 127774 8152
rect 80882 8032 80888 8084
rect 80940 8072 80946 8084
rect 127434 8072 127440 8084
rect 80940 8044 127440 8072
rect 80940 8032 80946 8044
rect 127434 8032 127440 8044
rect 127492 8032 127498 8084
rect 77386 7964 77392 8016
rect 77444 8004 77450 8016
rect 127526 8004 127532 8016
rect 77444 7976 127532 8004
rect 77444 7964 77450 7976
rect 127526 7964 127532 7976
rect 127584 7964 127590 8016
rect 73798 7896 73804 7948
rect 73856 7936 73862 7948
rect 127618 7936 127624 7948
rect 73856 7908 127624 7936
rect 73856 7896 73862 7908
rect 127618 7896 127624 7908
rect 127676 7896 127682 7948
rect 142430 7896 142436 7948
rect 142488 7936 142494 7948
rect 268838 7936 268844 7948
rect 142488 7908 268844 7936
rect 142488 7896 142494 7908
rect 268838 7896 268844 7908
rect 268896 7896 268902 7948
rect 66714 7828 66720 7880
rect 66772 7868 66778 7880
rect 126054 7868 126060 7880
rect 66772 7840 126060 7868
rect 66772 7828 66778 7840
rect 126054 7828 126060 7840
rect 126112 7828 126118 7880
rect 144086 7828 144092 7880
rect 144144 7868 144150 7880
rect 290182 7868 290188 7880
rect 144144 7840 290188 7868
rect 144144 7828 144150 7840
rect 290182 7828 290188 7840
rect 290240 7828 290246 7880
rect 63218 7760 63224 7812
rect 63276 7800 63282 7812
rect 125962 7800 125968 7812
rect 63276 7772 125968 7800
rect 63276 7760 63282 7772
rect 125962 7760 125968 7772
rect 126020 7760 126026 7812
rect 147674 7760 147680 7812
rect 147732 7800 147738 7812
rect 336274 7800 336280 7812
rect 147732 7772 336280 7800
rect 147732 7760 147738 7772
rect 336274 7760 336280 7772
rect 336332 7760 336338 7812
rect 27706 7692 27712 7744
rect 27764 7732 27770 7744
rect 123202 7732 123208 7744
rect 27764 7704 123208 7732
rect 27764 7692 27770 7704
rect 123202 7692 123208 7704
rect 123260 7692 123266 7744
rect 154022 7692 154028 7744
rect 154080 7732 154086 7744
rect 417878 7732 417884 7744
rect 154080 7704 417884 7732
rect 154080 7692 154086 7704
rect 417878 7692 417884 7704
rect 417936 7692 417942 7744
rect 19426 7624 19432 7676
rect 19484 7664 19490 7676
rect 118050 7664 118056 7676
rect 19484 7636 118056 7664
rect 19484 7624 19490 7636
rect 118050 7624 118056 7636
rect 118108 7624 118114 7676
rect 119890 7624 119896 7676
rect 119948 7664 119954 7676
rect 130102 7664 130108 7676
rect 119948 7636 130108 7664
rect 119948 7624 119954 7636
rect 130102 7624 130108 7636
rect 130160 7624 130166 7676
rect 164694 7624 164700 7676
rect 164752 7664 164758 7676
rect 554958 7664 554964 7676
rect 164752 7636 554964 7664
rect 164752 7624 164758 7636
rect 554958 7624 554964 7636
rect 555016 7624 555022 7676
rect 23014 7556 23020 7608
rect 23072 7596 23078 7608
rect 123294 7596 123300 7608
rect 23072 7568 123300 7596
rect 23072 7556 23078 7568
rect 123294 7556 123300 7568
rect 123352 7556 123358 7608
rect 164970 7556 164976 7608
rect 165028 7596 165034 7608
rect 558546 7596 558552 7608
rect 165028 7568 558552 7596
rect 165028 7556 165034 7568
rect 558546 7556 558552 7568
rect 558604 7556 558610 7608
rect 102226 7488 102232 7540
rect 102284 7528 102290 7540
rect 128814 7528 128820 7540
rect 102284 7500 128820 7528
rect 102284 7488 102290 7500
rect 128814 7488 128820 7500
rect 128872 7488 128878 7540
rect 115198 6808 115204 6860
rect 115256 6848 115262 6860
rect 130010 6848 130016 6860
rect 115256 6820 130016 6848
rect 115256 6808 115262 6820
rect 130010 6808 130016 6820
rect 130068 6808 130074 6860
rect 562318 6808 562324 6860
rect 562376 6848 562382 6860
rect 580166 6848 580172 6860
rect 562376 6820 580172 6848
rect 562376 6808 562382 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 99834 6740 99840 6792
rect 99892 6780 99898 6792
rect 120810 6780 120816 6792
rect 99892 6752 120816 6780
rect 99892 6740 99898 6752
rect 120810 6740 120816 6752
rect 120868 6740 120874 6792
rect 139854 6740 139860 6792
rect 139912 6780 139918 6792
rect 235810 6780 235816 6792
rect 139912 6752 235816 6780
rect 139912 6740 139918 6752
rect 235810 6740 235816 6752
rect 235868 6740 235874 6792
rect 59630 6672 59636 6724
rect 59688 6712 59694 6724
rect 125870 6712 125876 6724
rect 59688 6684 125876 6712
rect 59688 6672 59694 6684
rect 125870 6672 125876 6684
rect 125928 6672 125934 6724
rect 143810 6672 143816 6724
rect 143868 6712 143874 6724
rect 286594 6712 286600 6724
rect 143868 6684 286600 6712
rect 143868 6672 143874 6684
rect 286594 6672 286600 6684
rect 286652 6672 286658 6724
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 86218 6644 86224 6656
rect 11204 6616 86224 6644
rect 11204 6604 11210 6616
rect 86218 6604 86224 6616
rect 86276 6604 86282 6656
rect 104526 6604 104532 6656
rect 104584 6644 104590 6656
rect 128630 6644 128636 6656
rect 104584 6616 128636 6644
rect 104584 6604 104590 6616
rect 128630 6604 128636 6616
rect 128688 6604 128694 6656
rect 151078 6604 151084 6656
rect 151136 6644 151142 6656
rect 379974 6644 379980 6656
rect 151136 6616 379980 6644
rect 151136 6604 151142 6616
rect 379974 6604 379980 6616
rect 380032 6604 380038 6656
rect 48958 6536 48964 6588
rect 49016 6576 49022 6588
rect 124674 6576 124680 6588
rect 49016 6548 124680 6576
rect 49016 6536 49022 6548
rect 124674 6536 124680 6548
rect 124732 6536 124738 6588
rect 152366 6536 152372 6588
rect 152424 6576 152430 6588
rect 396534 6576 396540 6588
rect 152424 6548 396540 6576
rect 152424 6536 152430 6548
rect 396534 6536 396540 6548
rect 396592 6536 396598 6588
rect 44266 6468 44272 6520
rect 44324 6508 44330 6520
rect 124490 6508 124496 6520
rect 44324 6480 124496 6508
rect 44324 6468 44330 6480
rect 124490 6468 124496 6480
rect 124548 6468 124554 6520
rect 167270 6468 167276 6520
rect 167328 6508 167334 6520
rect 436738 6508 436744 6520
rect 167328 6480 436744 6508
rect 167328 6468 167334 6480
rect 436738 6468 436744 6480
rect 436796 6468 436802 6520
rect 40678 6400 40684 6452
rect 40736 6440 40742 6452
rect 124582 6440 124588 6452
rect 40736 6412 124588 6440
rect 40736 6400 40742 6412
rect 124582 6400 124588 6412
rect 124640 6400 124646 6452
rect 161566 6400 161572 6452
rect 161624 6440 161630 6452
rect 514754 6440 514760 6452
rect 161624 6412 514760 6440
rect 161624 6400 161630 6412
rect 514754 6400 514760 6412
rect 514812 6400 514818 6452
rect 30098 6332 30104 6384
rect 30156 6372 30162 6384
rect 123110 6372 123116 6384
rect 30156 6344 123116 6372
rect 30156 6332 30162 6344
rect 123110 6332 123116 6344
rect 123168 6332 123174 6384
rect 163590 6332 163596 6384
rect 163648 6372 163654 6384
rect 540790 6372 540796 6384
rect 163648 6344 540796 6372
rect 163648 6332 163654 6344
rect 540790 6332 540796 6344
rect 540848 6332 540854 6384
rect 13538 6264 13544 6316
rect 13596 6304 13602 6316
rect 121730 6304 121736 6316
rect 13596 6276 121736 6304
rect 13596 6264 13602 6276
rect 121730 6264 121736 6276
rect 121788 6264 121794 6316
rect 163866 6264 163872 6316
rect 163924 6304 163930 6316
rect 544378 6304 544384 6316
rect 163924 6276 544384 6304
rect 163924 6264 163930 6276
rect 544378 6264 544384 6276
rect 544436 6264 544442 6316
rect 8754 6196 8760 6248
rect 8812 6236 8818 6248
rect 121822 6236 121828 6248
rect 8812 6208 121828 6236
rect 8812 6196 8818 6208
rect 121822 6196 121828 6208
rect 121880 6196 121886 6248
rect 165798 6196 165804 6248
rect 165856 6236 165862 6248
rect 569126 6236 569132 6248
rect 165856 6208 569132 6236
rect 165856 6196 165862 6208
rect 569126 6196 569132 6208
rect 569184 6196 569190 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 121914 6168 121920 6180
rect 4120 6140 121920 6168
rect 4120 6128 4126 6140
rect 121914 6128 121920 6140
rect 121972 6128 121978 6180
rect 166074 6128 166080 6180
rect 166132 6168 166138 6180
rect 572714 6168 572720 6180
rect 166132 6140 572720 6168
rect 166132 6128 166138 6140
rect 572714 6128 572720 6140
rect 572772 6128 572778 6180
rect 97442 5448 97448 5500
rect 97500 5488 97506 5500
rect 129366 5488 129372 5500
rect 97500 5460 129372 5488
rect 97500 5448 97506 5460
rect 129366 5448 129372 5460
rect 129424 5448 129430 5500
rect 93946 5380 93952 5432
rect 94004 5420 94010 5432
rect 129274 5420 129280 5432
rect 94004 5392 129280 5420
rect 94004 5380 94010 5392
rect 129274 5380 129280 5392
rect 129332 5380 129338 5432
rect 132586 5380 132592 5432
rect 132644 5420 132650 5432
rect 142430 5420 142436 5432
rect 132644 5392 142436 5420
rect 132644 5380 132650 5392
rect 142430 5380 142436 5392
rect 142488 5380 142494 5432
rect 85666 5312 85672 5364
rect 85724 5352 85730 5364
rect 120718 5352 120724 5364
rect 85724 5324 120724 5352
rect 85724 5312 85730 5324
rect 120718 5312 120724 5324
rect 120776 5312 120782 5364
rect 132770 5312 132776 5364
rect 132828 5352 132834 5364
rect 144730 5352 144736 5364
rect 132828 5324 144736 5352
rect 132828 5312 132834 5324
rect 144730 5312 144736 5324
rect 144788 5312 144794 5364
rect 86862 5244 86868 5296
rect 86920 5284 86926 5296
rect 127342 5284 127348 5296
rect 86920 5256 127348 5284
rect 86920 5244 86926 5256
rect 127342 5244 127348 5256
rect 127400 5244 127406 5296
rect 134518 5244 134524 5296
rect 134576 5284 134582 5296
rect 167178 5284 167184 5296
rect 134576 5256 167184 5284
rect 134576 5244 134582 5256
rect 167178 5244 167184 5256
rect 167236 5244 167242 5296
rect 76190 5176 76196 5228
rect 76248 5216 76254 5228
rect 127158 5216 127164 5228
rect 76248 5188 127164 5216
rect 76248 5176 76254 5188
rect 127158 5176 127164 5188
rect 127216 5176 127222 5228
rect 137278 5176 137284 5228
rect 137336 5216 137342 5228
rect 202690 5216 202696 5228
rect 137336 5188 202696 5216
rect 137336 5176 137342 5188
rect 202690 5176 202696 5188
rect 202748 5176 202754 5228
rect 72602 5108 72608 5160
rect 72660 5148 72666 5160
rect 127250 5148 127256 5160
rect 72660 5120 127256 5148
rect 72660 5108 72666 5120
rect 127250 5108 127256 5120
rect 127308 5108 127314 5160
rect 133046 5108 133052 5160
rect 133104 5148 133110 5160
rect 148318 5148 148324 5160
rect 133104 5120 148324 5148
rect 133104 5108 133110 5120
rect 148318 5108 148324 5120
rect 148376 5108 148382 5160
rect 149882 5108 149888 5160
rect 149940 5148 149946 5160
rect 364610 5148 364616 5160
rect 149940 5120 364616 5148
rect 149940 5108 149946 5120
rect 364610 5108 364616 5120
rect 364668 5108 364674 5160
rect 65518 5040 65524 5092
rect 65576 5080 65582 5092
rect 125778 5080 125784 5092
rect 65576 5052 125784 5080
rect 65576 5040 65582 5052
rect 125778 5040 125784 5052
rect 125836 5040 125842 5092
rect 133138 5040 133144 5092
rect 133196 5080 133202 5092
rect 149514 5080 149520 5092
rect 133196 5052 149520 5080
rect 133196 5040 133202 5052
rect 149514 5040 149520 5052
rect 149572 5040 149578 5092
rect 160462 5040 160468 5092
rect 160520 5080 160526 5092
rect 500586 5080 500592 5092
rect 160520 5052 500592 5080
rect 160520 5040 160526 5052
rect 500586 5040 500592 5052
rect 500644 5040 500650 5092
rect 33594 4972 33600 5024
rect 33652 5012 33658 5024
rect 123018 5012 123024 5024
rect 33652 4984 123024 5012
rect 33652 4972 33658 4984
rect 123018 4972 123024 4984
rect 123076 4972 123082 5024
rect 133414 4972 133420 5024
rect 133472 5012 133478 5024
rect 153010 5012 153016 5024
rect 133472 4984 153016 5012
rect 133472 4972 133478 4984
rect 153010 4972 153016 4984
rect 153068 4972 153074 5024
rect 160554 4972 160560 5024
rect 160612 5012 160618 5024
rect 501782 5012 501788 5024
rect 160612 4984 501788 5012
rect 160612 4972 160618 4984
rect 501782 4972 501788 4984
rect 501840 4972 501846 5024
rect 28902 4904 28908 4956
rect 28960 4944 28966 4956
rect 117958 4944 117964 4956
rect 28960 4916 117964 4944
rect 28960 4904 28966 4916
rect 117958 4904 117964 4916
rect 118016 4904 118022 4956
rect 118786 4904 118792 4956
rect 118844 4944 118850 4956
rect 129918 4944 129924 4956
rect 118844 4916 129924 4944
rect 118844 4904 118850 4916
rect 129918 4904 129924 4916
rect 129976 4904 129982 4956
rect 133322 4904 133328 4956
rect 133380 4944 133386 4956
rect 151814 4944 151820 4956
rect 133380 4916 151820 4944
rect 133380 4904 133386 4916
rect 151814 4904 151820 4916
rect 151872 4904 151878 4956
rect 161934 4904 161940 4956
rect 161992 4944 161998 4956
rect 519538 4944 519544 4956
rect 161992 4916 519544 4944
rect 161992 4904 161998 4916
rect 519538 4904 519544 4916
rect 519596 4904 519602 4956
rect 5258 4836 5264 4888
rect 5316 4876 5322 4888
rect 22738 4876 22744 4888
rect 5316 4848 22744 4876
rect 5316 4836 5322 4848
rect 22738 4836 22744 4848
rect 22796 4836 22802 4888
rect 26510 4836 26516 4888
rect 26568 4876 26574 4888
rect 124122 4876 124128 4888
rect 26568 4848 124128 4876
rect 26568 4836 26574 4848
rect 124122 4836 124128 4848
rect 124180 4836 124186 4888
rect 133874 4836 133880 4888
rect 133932 4876 133938 4888
rect 158898 4876 158904 4888
rect 133932 4848 158904 4876
rect 133932 4836 133938 4848
rect 158898 4836 158904 4848
rect 158956 4836 158962 4888
rect 162210 4836 162216 4888
rect 162268 4876 162274 4888
rect 523034 4876 523040 4888
rect 162268 4848 523040 4876
rect 162268 4836 162274 4848
rect 523034 4836 523040 4848
rect 523092 4836 523098 4888
rect 21818 4768 21824 4820
rect 21876 4808 21882 4820
rect 123754 4808 123760 4820
rect 21876 4780 123760 4808
rect 21876 4768 21882 4780
rect 123754 4768 123760 4780
rect 123812 4768 123818 4820
rect 134242 4768 134248 4820
rect 134300 4808 134306 4820
rect 163682 4808 163688 4820
rect 134300 4780 163688 4808
rect 134300 4768 134306 4780
rect 163682 4768 163688 4780
rect 163740 4768 163746 4820
rect 166810 4768 166816 4820
rect 166868 4808 166874 4820
rect 577406 4808 577412 4820
rect 166868 4780 577412 4808
rect 166868 4768 166874 4780
rect 577406 4768 577412 4780
rect 577464 4768 577470 4820
rect 111610 4700 111616 4752
rect 111668 4740 111674 4752
rect 129826 4740 129832 4752
rect 111668 4712 129832 4740
rect 111668 4700 111674 4712
rect 129826 4700 129832 4712
rect 129884 4700 129890 4752
rect 117222 4632 117228 4684
rect 117280 4672 117286 4684
rect 128538 4672 128544 4684
rect 117280 4644 128544 4672
rect 117280 4632 117286 4644
rect 128538 4632 128544 4644
rect 128596 4632 128602 4684
rect 101030 4088 101036 4140
rect 101088 4128 101094 4140
rect 117222 4128 117228 4140
rect 101088 4100 117228 4128
rect 101088 4088 101094 4100
rect 117222 4088 117228 4100
rect 117280 4088 117286 4140
rect 121362 4088 121368 4140
rect 121420 4128 121426 4140
rect 143534 4128 143540 4140
rect 121420 4100 143540 4128
rect 121420 4088 121426 4100
rect 143534 4088 143540 4100
rect 143592 4088 143598 4140
rect 168098 4088 168104 4140
rect 168156 4128 168162 4140
rect 189718 4128 189724 4140
rect 168156 4100 189724 4128
rect 168156 4088 168162 4100
rect 189718 4088 189724 4100
rect 189776 4088 189782 4140
rect 276014 4088 276020 4140
rect 276072 4128 276078 4140
rect 276750 4128 276756 4140
rect 276072 4100 276756 4128
rect 276072 4088 276078 4100
rect 276750 4088 276756 4100
rect 276808 4088 276814 4140
rect 284294 4088 284300 4140
rect 284352 4128 284358 4140
rect 285030 4128 285036 4140
rect 284352 4100 285036 4128
rect 284352 4088 284358 4100
rect 285030 4088 285036 4100
rect 285088 4088 285094 4140
rect 292574 4088 292580 4140
rect 292632 4128 292638 4140
rect 293310 4128 293316 4140
rect 292632 4100 293316 4128
rect 292632 4088 292638 4100
rect 293310 4088 293316 4100
rect 293368 4088 293374 4140
rect 312538 4088 312544 4140
rect 312596 4128 312602 4140
rect 543182 4128 543188 4140
rect 312596 4100 543188 4128
rect 312596 4088 312602 4100
rect 543182 4088 543188 4100
rect 543240 4088 543246 4140
rect 83274 4020 83280 4072
rect 83332 4060 83338 4072
rect 127986 4060 127992 4072
rect 83332 4032 127992 4060
rect 83332 4020 83338 4032
rect 127986 4020 127992 4032
rect 128044 4020 128050 4072
rect 131850 4020 131856 4072
rect 131908 4060 131914 4072
rect 132954 4060 132960 4072
rect 131908 4032 132960 4060
rect 131908 4020 131914 4032
rect 132954 4020 132960 4032
rect 133012 4020 133018 4072
rect 133064 4032 135576 4060
rect 79686 3952 79692 4004
rect 79744 3992 79750 4004
rect 127066 3992 127072 4004
rect 79744 3964 127072 3992
rect 79744 3952 79750 3964
rect 127066 3952 127072 3964
rect 127124 3952 127130 4004
rect 132862 3952 132868 4004
rect 132920 3992 132926 4004
rect 133064 3992 133092 4032
rect 132920 3964 133092 3992
rect 132920 3952 132926 3964
rect 134058 3952 134064 4004
rect 134116 3992 134122 4004
rect 135548 3992 135576 4032
rect 146938 4020 146944 4072
rect 146996 4060 147002 4072
rect 160094 4060 160100 4072
rect 146996 4032 160100 4060
rect 146996 4020 147002 4032
rect 160094 4020 160100 4032
rect 160152 4020 160158 4072
rect 167454 4020 167460 4072
rect 167512 4060 167518 4072
rect 401318 4060 401324 4072
rect 167512 4032 401324 4060
rect 167512 4020 167518 4032
rect 401318 4020 401324 4032
rect 401376 4020 401382 4072
rect 145926 3992 145932 4004
rect 134116 3964 135484 3992
rect 135548 3964 145932 3992
rect 134116 3952 134122 3964
rect 69106 3884 69112 3936
rect 69164 3924 69170 3936
rect 126882 3924 126888 3936
rect 69164 3896 126888 3924
rect 69164 3884 69170 3896
rect 126882 3884 126888 3896
rect 126940 3884 126946 3936
rect 132034 3884 132040 3936
rect 132092 3924 132098 3936
rect 135254 3924 135260 3936
rect 132092 3896 135260 3924
rect 132092 3884 132098 3896
rect 135254 3884 135260 3896
rect 135312 3884 135318 3936
rect 135456 3924 135484 3964
rect 145926 3952 145932 3964
rect 145984 3952 145990 4004
rect 167546 3952 167552 4004
rect 167604 3992 167610 4004
rect 408402 3992 408408 4004
rect 167604 3964 408408 3992
rect 167604 3952 167610 3964
rect 408402 3952 408408 3964
rect 408460 3952 408466 4004
rect 161290 3924 161296 3936
rect 135456 3896 161296 3924
rect 161290 3884 161296 3896
rect 161348 3884 161354 3936
rect 168190 3884 168196 3936
rect 168248 3924 168254 3936
rect 409598 3924 409604 3936
rect 168248 3896 409604 3924
rect 168248 3884 168254 3896
rect 409598 3884 409604 3896
rect 409656 3884 409662 3936
rect 58434 3816 58440 3868
rect 58492 3856 58498 3868
rect 126514 3856 126520 3868
rect 58492 3828 126520 3856
rect 58492 3816 58498 3828
rect 126514 3816 126520 3828
rect 126572 3816 126578 3868
rect 134150 3816 134156 3868
rect 134208 3856 134214 3868
rect 162486 3856 162492 3868
rect 134208 3828 162492 3856
rect 134208 3816 134214 3828
rect 162486 3816 162492 3828
rect 162544 3816 162550 3868
rect 168282 3816 168288 3868
rect 168340 3856 168346 3868
rect 415394 3856 415400 3868
rect 168340 3828 415400 3856
rect 168340 3816 168346 3828
rect 415394 3816 415400 3828
rect 415452 3816 415458 3868
rect 51350 3748 51356 3800
rect 51408 3788 51414 3800
rect 125502 3788 125508 3800
rect 51408 3760 125508 3788
rect 51408 3748 51414 3760
rect 125502 3748 125508 3760
rect 125560 3748 125566 3800
rect 134334 3748 134340 3800
rect 134392 3788 134398 3800
rect 164878 3788 164884 3800
rect 134392 3760 164884 3788
rect 134392 3748 134398 3760
rect 164878 3748 164884 3760
rect 164936 3748 164942 3800
rect 167638 3748 167644 3800
rect 167696 3788 167702 3800
rect 427262 3788 427268 3800
rect 167696 3760 427268 3788
rect 167696 3748 167702 3760
rect 427262 3748 427268 3760
rect 427320 3748 427326 3800
rect 47854 3680 47860 3732
rect 47912 3720 47918 3732
rect 124306 3720 124312 3732
rect 47912 3692 124312 3720
rect 47912 3680 47918 3692
rect 124306 3680 124312 3692
rect 124364 3680 124370 3732
rect 134426 3680 134432 3732
rect 134484 3720 134490 3732
rect 166074 3720 166080 3732
rect 134484 3692 166080 3720
rect 134484 3680 134490 3692
rect 166074 3680 166080 3692
rect 166132 3680 166138 3732
rect 167730 3680 167736 3732
rect 167788 3720 167794 3732
rect 429654 3720 429660 3732
rect 167788 3692 429660 3720
rect 167788 3680 167794 3692
rect 429654 3680 429660 3692
rect 429712 3680 429718 3732
rect 445110 3680 445116 3732
rect 445168 3720 445174 3732
rect 546678 3720 546684 3732
rect 445168 3692 546684 3720
rect 445168 3680 445174 3692
rect 546678 3680 546684 3692
rect 546736 3680 546742 3732
rect 39574 3612 39580 3664
rect 39632 3652 39638 3664
rect 125226 3652 125232 3664
rect 39632 3624 125232 3652
rect 39632 3612 39638 3624
rect 125226 3612 125232 3624
rect 125284 3612 125290 3664
rect 134610 3612 134616 3664
rect 134668 3652 134674 3664
rect 168374 3652 168380 3664
rect 134668 3624 168380 3652
rect 134668 3612 134674 3624
rect 168374 3612 168380 3624
rect 168432 3612 168438 3664
rect 169018 3612 169024 3664
rect 169076 3652 169082 3664
rect 465166 3652 465172 3664
rect 169076 3624 465172 3652
rect 169076 3612 169082 3624
rect 465166 3612 465172 3624
rect 465224 3612 465230 3664
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 122466 3584 122472 3596
rect 12400 3556 122472 3584
rect 12400 3544 12406 3556
rect 122466 3544 122472 3556
rect 122524 3544 122530 3596
rect 125870 3544 125876 3596
rect 125928 3584 125934 3596
rect 131114 3584 131120 3596
rect 125928 3556 131120 3584
rect 125928 3544 125934 3556
rect 131114 3544 131120 3556
rect 131172 3544 131178 3596
rect 133046 3544 133052 3596
rect 133104 3584 133110 3596
rect 147122 3584 147128 3596
rect 133104 3556 147128 3584
rect 133104 3544 133110 3556
rect 147122 3544 147128 3556
rect 147180 3544 147186 3596
rect 159174 3544 159180 3596
rect 159232 3584 159238 3596
rect 484026 3584 484032 3596
rect 159232 3556 484032 3584
rect 159232 3544 159238 3556
rect 484026 3544 484032 3556
rect 484084 3544 484090 3596
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 122558 3516 122564 3528
rect 7708 3488 122564 3516
rect 7708 3476 7714 3488
rect 122558 3476 122564 3488
rect 122616 3476 122622 3528
rect 129366 3476 129372 3528
rect 129424 3516 129430 3528
rect 131206 3516 131212 3528
rect 129424 3488 131212 3516
rect 129424 3476 129430 3488
rect 131206 3476 131212 3488
rect 131264 3476 131270 3528
rect 133230 3476 133236 3528
rect 133288 3516 133294 3528
rect 150618 3516 150624 3528
rect 133288 3488 150624 3516
rect 133288 3476 133294 3488
rect 150618 3476 150624 3488
rect 150676 3476 150682 3528
rect 159450 3476 159456 3528
rect 159508 3516 159514 3528
rect 478046 3516 478052 3528
rect 159508 3488 478052 3516
rect 159508 3476 159514 3488
rect 478046 3476 478052 3488
rect 478104 3476 478110 3528
rect 478156 3488 483014 3516
rect 2866 3408 2872 3460
rect 2924 3448 2930 3460
rect 122190 3448 122196 3460
rect 2924 3420 122196 3448
rect 2924 3408 2930 3420
rect 122190 3408 122196 3420
rect 122248 3408 122254 3460
rect 126974 3408 126980 3460
rect 127032 3448 127038 3460
rect 131390 3448 131396 3460
rect 127032 3420 131396 3448
rect 127032 3408 127038 3420
rect 131390 3408 131396 3420
rect 131448 3408 131454 3460
rect 133506 3408 133512 3460
rect 133564 3448 133570 3460
rect 154206 3448 154212 3460
rect 133564 3420 154212 3448
rect 133564 3408 133570 3420
rect 154206 3408 154212 3420
rect 154264 3408 154270 3460
rect 159726 3408 159732 3460
rect 159784 3448 159790 3460
rect 478156 3448 478184 3488
rect 159784 3420 478184 3448
rect 482986 3448 483014 3488
rect 491110 3448 491116 3460
rect 482986 3420 491116 3448
rect 159784 3408 159790 3420
rect 491110 3408 491116 3420
rect 491168 3408 491174 3460
rect 102134 3340 102140 3392
rect 102192 3380 102198 3392
rect 103330 3380 103336 3392
rect 102192 3352 103336 3380
rect 102192 3340 102198 3352
rect 103330 3340 103336 3352
rect 103388 3340 103394 3392
rect 122282 3340 122288 3392
rect 122340 3380 122346 3392
rect 131022 3380 131028 3392
rect 122340 3352 131028 3380
rect 122340 3340 122346 3352
rect 131022 3340 131028 3352
rect 131080 3340 131086 3392
rect 131942 3340 131948 3392
rect 132000 3380 132006 3392
rect 134150 3380 134156 3392
rect 132000 3352 134156 3380
rect 132000 3340 132006 3352
rect 134150 3340 134156 3352
rect 134208 3340 134214 3392
rect 137738 3340 137744 3392
rect 137796 3380 137802 3392
rect 146938 3380 146944 3392
rect 137796 3352 146944 3380
rect 137796 3340 137802 3352
rect 146938 3340 146944 3352
rect 146996 3340 147002 3392
rect 167362 3340 167368 3392
rect 167420 3380 167426 3392
rect 394234 3380 394240 3392
rect 167420 3352 394240 3380
rect 167420 3340 167426 3352
rect 394234 3340 394240 3352
rect 394292 3340 394298 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 415486 3340 415492 3392
rect 415544 3380 415550 3392
rect 416682 3380 416688 3392
rect 415544 3352 416688 3380
rect 415544 3340 415550 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 432046 3340 432052 3392
rect 432104 3380 432110 3392
rect 433242 3380 433248 3392
rect 432104 3352 433248 3380
rect 432104 3340 432110 3352
rect 433242 3340 433248 3352
rect 433300 3340 433306 3392
rect 440326 3340 440332 3392
rect 440384 3380 440390 3392
rect 441522 3380 441528 3392
rect 440384 3352 441528 3380
rect 440384 3340 440390 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 456794 3340 456800 3392
rect 456852 3380 456858 3392
rect 458082 3380 458088 3392
rect 456852 3352 458088 3380
rect 456852 3340 456858 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 473354 3340 473360 3392
rect 473412 3380 473418 3392
rect 474182 3380 474188 3392
rect 473412 3352 474188 3380
rect 473412 3340 473418 3352
rect 474182 3340 474188 3352
rect 474240 3340 474246 3392
rect 478046 3340 478052 3392
rect 478104 3380 478110 3392
rect 487614 3380 487620 3392
rect 478104 3352 487620 3380
rect 478104 3340 478110 3352
rect 487614 3340 487620 3352
rect 487672 3340 487678 3392
rect 130562 3272 130568 3324
rect 130620 3312 130626 3324
rect 131482 3312 131488 3324
rect 130620 3284 131488 3312
rect 130620 3272 130626 3284
rect 131482 3272 131488 3284
rect 131540 3272 131546 3324
rect 132126 3272 132132 3324
rect 132184 3312 132190 3324
rect 136450 3312 136456 3324
rect 132184 3284 136456 3312
rect 132184 3272 132190 3284
rect 136450 3272 136456 3284
rect 136508 3272 136514 3324
rect 149146 3272 149152 3324
rect 149204 3312 149210 3324
rect 169570 3312 169576 3324
rect 149204 3284 169576 3312
rect 149204 3272 149210 3284
rect 169570 3272 169576 3284
rect 169628 3272 169634 3324
rect 169662 3272 169668 3324
rect 169720 3312 169726 3324
rect 175458 3312 175464 3324
rect 169720 3284 175464 3312
rect 169720 3272 169726 3284
rect 175458 3272 175464 3284
rect 175516 3272 175522 3324
rect 193214 3272 193220 3324
rect 193272 3312 193278 3324
rect 194410 3312 194416 3324
rect 193272 3284 194416 3312
rect 193272 3272 193278 3284
rect 194410 3272 194416 3284
rect 194468 3272 194474 3324
rect 226334 3272 226340 3324
rect 226392 3312 226398 3324
rect 227530 3312 227536 3324
rect 226392 3284 227536 3312
rect 226392 3272 226398 3284
rect 227530 3272 227536 3284
rect 227588 3272 227594 3324
rect 299474 3272 299480 3324
rect 299532 3312 299538 3324
rect 300762 3312 300768 3324
rect 299532 3284 300768 3312
rect 299532 3272 299538 3284
rect 300762 3272 300768 3284
rect 300820 3272 300826 3324
rect 307754 3272 307760 3324
rect 307812 3312 307818 3324
rect 309042 3312 309048 3324
rect 307812 3284 309048 3312
rect 307812 3272 307818 3284
rect 309042 3272 309048 3284
rect 309100 3272 309106 3324
rect 316034 3272 316040 3324
rect 316092 3312 316098 3324
rect 317322 3312 317328 3324
rect 316092 3284 317328 3312
rect 316092 3272 316098 3284
rect 317322 3272 317328 3284
rect 317380 3272 317386 3324
rect 324406 3272 324412 3324
rect 324464 3312 324470 3324
rect 325602 3312 325608 3324
rect 324464 3284 325608 3312
rect 324464 3272 324470 3284
rect 325602 3272 325608 3284
rect 325660 3272 325666 3324
rect 332594 3272 332600 3324
rect 332652 3312 332658 3324
rect 333882 3312 333888 3324
rect 332652 3284 333888 3312
rect 332652 3272 332658 3284
rect 333882 3272 333888 3284
rect 333940 3272 333946 3324
rect 539594 3312 539600 3324
rect 335326 3284 539600 3312
rect 20622 3204 20628 3256
rect 20680 3244 20686 3256
rect 25498 3244 25504 3256
rect 20680 3216 25504 3244
rect 20680 3204 20686 3216
rect 25498 3204 25504 3216
rect 25556 3204 25562 3256
rect 165246 3204 165252 3256
rect 165304 3244 165310 3256
rect 182542 3244 182548 3256
rect 165304 3216 182548 3244
rect 165304 3204 165310 3216
rect 182542 3204 182548 3216
rect 182600 3204 182606 3256
rect 326430 3204 326436 3256
rect 326488 3244 326494 3256
rect 335326 3244 335354 3284
rect 539594 3272 539600 3284
rect 539652 3272 539658 3324
rect 326488 3216 335354 3244
rect 326488 3204 326494 3216
rect 349154 3204 349160 3256
rect 349212 3244 349218 3256
rect 350442 3244 350448 3256
rect 349212 3216 350448 3244
rect 349212 3204 349218 3216
rect 350442 3204 350448 3216
rect 350500 3204 350506 3256
rect 357434 3204 357440 3256
rect 357492 3244 357498 3256
rect 358722 3244 358728 3256
rect 357492 3216 358728 3244
rect 357492 3204 357498 3216
rect 358722 3204 358728 3216
rect 358780 3204 358786 3256
rect 365714 3204 365720 3256
rect 365772 3244 365778 3256
rect 367002 3244 367008 3256
rect 365772 3216 367008 3244
rect 365772 3204 365778 3216
rect 367002 3204 367008 3216
rect 367060 3204 367066 3256
rect 374086 3204 374092 3256
rect 374144 3244 374150 3256
rect 375282 3244 375288 3256
rect 374144 3216 375288 3244
rect 374144 3204 374150 3216
rect 375282 3204 375288 3216
rect 375340 3204 375346 3256
rect 382274 3204 382280 3256
rect 382332 3244 382338 3256
rect 383562 3244 383568 3256
rect 382332 3216 383568 3244
rect 382332 3204 382338 3216
rect 383562 3204 383568 3216
rect 383620 3204 383626 3256
rect 390554 3204 390560 3256
rect 390612 3244 390618 3256
rect 391842 3244 391848 3256
rect 390612 3216 391848 3244
rect 390612 3204 390618 3216
rect 391842 3204 391848 3216
rect 391900 3204 391906 3256
rect 128170 3136 128176 3188
rect 128228 3176 128234 3188
rect 131574 3176 131580 3188
rect 128228 3148 131580 3176
rect 128228 3136 128234 3148
rect 131574 3136 131580 3148
rect 131632 3136 131638 3188
rect 136174 2932 136180 2984
rect 136232 2972 136238 2984
rect 141234 2972 141240 2984
rect 136232 2944 141240 2972
rect 136232 2932 136238 2944
rect 141234 2932 141240 2944
rect 141292 2932 141298 2984
rect 423674 1232 423680 1284
rect 423732 1272 423738 1284
rect 424962 1272 424968 1284
rect 423732 1244 424968 1272
rect 423732 1232 423738 1244
rect 424962 1232 424968 1244
rect 425020 1232 425026 1284
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 410524 700408 410576 700460
rect 429844 700408 429896 700460
rect 409144 700340 409196 700392
rect 494796 700340 494848 700392
rect 155224 700272 155276 700324
rect 202788 700272 202840 700324
rect 332508 700272 332560 700324
rect 340144 700272 340196 700324
rect 407764 700272 407816 700324
rect 559656 700272 559708 700324
rect 153016 699660 153068 699712
rect 154120 699660 154172 699712
rect 149704 697688 149756 697740
rect 153016 697688 153068 697740
rect 282184 696328 282236 696380
rect 283840 696328 283892 696380
rect 348792 696192 348844 696244
rect 359464 696192 359516 696244
rect 264244 695104 264296 695156
rect 267648 695104 267700 695156
rect 299480 694764 299532 694816
rect 309784 694764 309836 694816
rect 278688 687148 278740 687200
rect 282184 687216 282236 687268
rect 359464 686468 359516 686520
rect 371884 686468 371936 686520
rect 309784 685108 309836 685160
rect 327724 685108 327776 685160
rect 276664 684496 276716 684548
rect 278688 684496 278740 684548
rect 364340 683748 364392 683800
rect 375380 683748 375432 683800
rect 371884 679600 371936 679652
rect 381544 679600 381596 679652
rect 375380 678240 375432 678292
rect 388444 678240 388496 678292
rect 140780 675452 140832 675504
rect 155224 675452 155276 675504
rect 145564 673412 145616 673464
rect 149704 673480 149756 673532
rect 212540 673412 212592 673464
rect 217968 673480 218020 673532
rect 134524 672052 134576 672104
rect 140780 672052 140832 672104
rect 388444 671100 388496 671152
rect 391940 671100 391992 671152
rect 3516 670692 3568 670744
rect 15844 670692 15896 670744
rect 566464 670692 566516 670744
rect 580172 670692 580224 670744
rect 211068 667836 211120 667888
rect 212540 667904 212592 667956
rect 226984 665796 227036 665848
rect 234620 665796 234672 665848
rect 391940 665184 391992 665236
rect 395344 665184 395396 665236
rect 209044 663756 209096 663808
rect 211068 663756 211120 663808
rect 258724 658180 258776 658232
rect 264244 658180 264296 658232
rect 143172 658112 143224 658164
rect 145564 658112 145616 658164
rect 141424 655528 141476 655580
rect 143172 655528 143224 655580
rect 327724 655460 327776 655512
rect 332692 655460 332744 655512
rect 131764 651856 131816 651908
rect 134524 651856 134576 651908
rect 332692 649952 332744 650004
rect 337384 649952 337436 650004
rect 381544 646484 381596 646536
rect 395528 646484 395580 646536
rect 204904 644376 204956 644428
rect 209044 644444 209096 644496
rect 337384 642132 337436 642184
rect 343640 642132 343692 642184
rect 139400 641724 139452 641776
rect 141424 641724 141476 641776
rect 340144 640976 340196 641028
rect 352564 640976 352616 641028
rect 224224 640296 224276 640348
rect 226984 640296 227036 640348
rect 343640 639548 343692 639600
rect 349160 639548 349212 639600
rect 136548 638868 136600 638920
rect 139400 638936 139452 638988
rect 349160 637508 349212 637560
rect 352656 637508 352708 637560
rect 134524 635536 134576 635588
rect 136548 635536 136600 635588
rect 211804 634040 211856 634092
rect 224224 634040 224276 634092
rect 247040 634040 247092 634092
rect 258724 634040 258776 634092
rect 203524 630640 203576 630692
rect 204904 630640 204956 630692
rect 275376 630640 275428 630692
rect 276664 630640 276716 630692
rect 243544 629620 243596 629672
rect 247040 629620 247092 629672
rect 273904 628736 273956 628788
rect 275376 628736 275428 628788
rect 352656 624384 352708 624436
rect 370504 624384 370556 624436
rect 209044 623772 209096 623824
rect 211804 623772 211856 623824
rect 352564 623024 352616 623076
rect 360200 623024 360252 623076
rect 271144 622412 271196 622464
rect 273904 622412 273956 622464
rect 123484 620984 123536 621036
rect 131764 620984 131816 621036
rect 360200 619556 360252 619608
rect 362960 619556 363012 619608
rect 3516 618264 3568 618316
rect 37924 618264 37976 618316
rect 406384 616836 406436 616888
rect 579988 616836 580040 616888
rect 362960 616088 363012 616140
rect 373264 616088 373316 616140
rect 233148 613368 233200 613420
rect 243544 613368 243596 613420
rect 268384 612756 268436 612808
rect 271144 612756 271196 612808
rect 200764 610512 200816 610564
rect 203524 610512 203576 610564
rect 59268 609220 59320 609272
rect 123484 609220 123536 609272
rect 224224 609220 224276 609272
rect 233148 609220 233200 609272
rect 53104 606432 53156 606484
rect 59268 606432 59320 606484
rect 267004 604460 267056 604512
rect 268384 604460 268436 604512
rect 370504 602352 370556 602404
rect 387064 602352 387116 602404
rect 373264 599564 373316 599616
rect 397552 599564 397604 599616
rect 131764 597524 131816 597576
rect 134524 597524 134576 597576
rect 195244 593308 195296 593360
rect 200764 593308 200816 593360
rect 214564 591268 214616 591320
rect 224224 591268 224276 591320
rect 211804 585148 211856 585200
rect 214564 585148 214616 585200
rect 200764 583720 200816 583772
rect 209044 583720 209096 583772
rect 387064 573996 387116 574048
rect 393964 573996 394016 574048
rect 265716 572704 265768 572756
rect 267004 572704 267056 572756
rect 264244 570664 264296 570716
rect 265716 570664 265768 570716
rect 3332 565836 3384 565888
rect 29644 565836 29696 565888
rect 198004 564952 198056 565004
rect 200764 564952 200816 565004
rect 405004 563048 405056 563100
rect 580172 563048 580224 563100
rect 393964 562640 394016 562692
rect 395436 562640 395488 562692
rect 193956 560260 194008 560312
rect 195244 560260 195296 560312
rect 46204 559716 46256 559768
rect 53104 559716 53156 559768
rect 192484 558560 192536 558612
rect 193956 558560 194008 558612
rect 2780 553800 2832 553852
rect 4804 553800 4856 553852
rect 261484 553392 261536 553444
rect 264244 553392 264296 553444
rect 206284 549244 206336 549296
rect 211804 549244 211856 549296
rect 191104 546456 191156 546508
rect 192484 546456 192536 546508
rect 189724 538840 189776 538892
rect 198004 538840 198056 538892
rect 62672 537480 62724 537532
rect 169760 537480 169812 537532
rect 188344 535100 188396 535152
rect 191104 535100 191156 535152
rect 130384 533332 130436 533384
rect 131764 533332 131816 533384
rect 61384 532992 61436 533044
rect 62672 532992 62724 533044
rect 260104 531224 260156 531276
rect 261484 531224 261536 531276
rect 129004 527144 129056 527196
rect 130384 527144 130436 527196
rect 200764 524424 200816 524476
rect 206284 524424 206336 524476
rect 257344 518916 257396 518968
rect 260104 518916 260156 518968
rect 45100 517488 45152 517540
rect 46204 517488 46256 517540
rect 3332 514768 3384 514820
rect 33784 514768 33836 514820
rect 153200 511232 153252 511284
rect 189724 511232 189776 511284
rect 403624 510620 403676 510672
rect 579804 510620 579856 510672
rect 117964 508512 118016 508564
rect 136640 508512 136692 508564
rect 150440 507832 150492 507884
rect 153200 507832 153252 507884
rect 192484 505724 192536 505776
rect 200764 505724 200816 505776
rect 253940 502256 253992 502308
rect 257344 502324 257396 502376
rect 143540 501712 143592 501764
rect 150440 501712 150492 501764
rect 2780 501032 2832 501084
rect 4896 501032 4948 501084
rect 126980 500896 127032 500948
rect 129004 500896 129056 500948
rect 180064 498788 180116 498840
rect 192484 498788 192536 498840
rect 249524 498108 249576 498160
rect 253940 498176 253992 498228
rect 124864 496748 124916 496800
rect 126980 496816 127032 496868
rect 140044 496680 140096 496732
rect 143540 496680 143592 496732
rect 246304 495456 246356 495508
rect 249524 495456 249576 495508
rect 116584 487160 116636 487212
rect 117964 487160 118016 487212
rect 136456 487160 136508 487212
rect 140044 487160 140096 487212
rect 175924 481992 175976 482044
rect 180064 481992 180116 482044
rect 133144 481448 133196 481500
rect 136456 481448 136508 481500
rect 123484 473968 123536 474020
rect 124864 473968 124916 474020
rect 115204 472948 115256 473000
rect 116584 472948 116636 473000
rect 239404 471928 239456 471980
rect 246304 471996 246356 472048
rect 122104 464992 122156 465044
rect 123484 464992 123536 465044
rect 2780 462544 2832 462596
rect 5080 462544 5132 462596
rect 163504 460164 163556 460216
rect 175924 460164 175976 460216
rect 400864 456764 400916 456816
rect 579988 456764 580040 456816
rect 182824 455336 182876 455388
rect 188344 455404 188396 455456
rect 238024 451256 238076 451308
rect 239404 451256 239456 451308
rect 127624 449896 127676 449948
rect 133144 449896 133196 449948
rect 2780 448808 2832 448860
rect 4988 448808 5040 448860
rect 160744 446972 160796 447024
rect 163504 446972 163556 447024
rect 119436 446156 119488 446208
rect 122104 446156 122156 446208
rect 399484 444388 399536 444440
rect 579988 444388 580040 444440
rect 181444 438880 181496 438932
rect 182824 438880 182876 438932
rect 117964 433236 118016 433288
rect 119436 433236 119488 433288
rect 119344 432556 119396 432608
rect 127624 432556 127676 432608
rect 236644 427796 236696 427848
rect 238024 427796 238076 427848
rect 116584 416712 116636 416764
rect 117964 416712 118016 416764
rect 179328 413992 179380 414044
rect 181444 413992 181496 414044
rect 3148 410048 3200 410100
rect 8944 410048 8996 410100
rect 177304 409844 177356 409896
rect 179328 409844 179380 409896
rect 115296 407192 115348 407244
rect 116584 407192 116636 407244
rect 113916 405424 113968 405476
rect 115296 405424 115348 405476
rect 417424 404336 417476 404388
rect 579988 404336 580040 404388
rect 233884 404268 233936 404320
rect 236644 404268 236696 404320
rect 112444 398488 112496 398540
rect 113916 398488 113968 398540
rect 2780 397468 2832 397520
rect 5172 397468 5224 397520
rect 110420 391960 110472 392012
rect 112444 391960 112496 392012
rect 112444 385636 112496 385688
rect 119344 385636 119396 385688
rect 106924 384616 106976 384668
rect 110420 384616 110472 384668
rect 157984 379516 158036 379568
rect 160744 379516 160796 379568
rect 396724 378156 396776 378208
rect 579988 378156 580040 378208
rect 58624 376592 58676 376644
rect 61384 376592 61436 376644
rect 175280 375300 175332 375352
rect 177304 375300 177356 375352
rect 173164 371152 173216 371204
rect 175280 371220 175332 371272
rect 103520 365644 103572 365696
rect 112444 365644 112496 365696
rect 396908 364352 396960 364404
rect 579988 364352 580040 364404
rect 78588 362176 78640 362228
rect 103520 362176 103572 362228
rect 75184 357756 75236 357808
rect 78588 357756 78640 357808
rect 105268 357552 105320 357604
rect 106924 357552 106976 357604
rect 3332 357416 3384 357468
rect 10324 357416 10376 357468
rect 69664 356668 69716 356720
rect 115204 356668 115256 356720
rect 103520 355784 103572 355836
rect 105268 355784 105320 355836
rect 414664 351908 414716 351960
rect 579988 351908 580040 351960
rect 98644 351840 98696 351892
rect 103520 351840 103572 351892
rect 231124 349460 231176 349512
rect 233884 349460 233936 349512
rect 172152 349120 172204 349172
rect 173164 349120 173216 349172
rect 56876 346332 56928 346384
rect 58624 346332 58676 346384
rect 2780 345176 2832 345228
rect 5264 345176 5316 345228
rect 170404 345040 170456 345092
rect 172152 345040 172204 345092
rect 94504 340892 94556 340944
rect 98644 340892 98696 340944
rect 68284 339668 68336 339720
rect 69664 339668 69716 339720
rect 55864 338240 55916 338292
rect 56876 338240 56928 338292
rect 566556 338104 566608 338156
rect 579988 338104 580040 338156
rect 66260 335996 66312 336048
rect 75184 335996 75236 336048
rect 48964 331848 49016 331900
rect 66260 331848 66312 331900
rect 167644 330352 167696 330404
rect 170404 330352 170456 330404
rect 396816 324300 396868 324352
rect 579804 324300 579856 324352
rect 53104 323348 53156 323400
rect 55864 323348 55916 323400
rect 165620 322940 165672 322992
rect 167644 322940 167696 322992
rect 228364 321512 228416 321564
rect 231124 321580 231176 321632
rect 162124 320424 162176 320476
rect 165620 320424 165672 320476
rect 85580 318112 85632 318164
rect 88340 318112 88392 318164
rect 62764 313896 62816 313948
rect 104900 313896 104952 313948
rect 79324 313352 79376 313404
rect 85580 313352 85632 313404
rect 397092 311856 397144 311908
rect 561956 311856 562008 311908
rect 562232 311856 562284 311908
rect 579988 311856 580040 311908
rect 93124 311516 93176 311568
rect 94504 311516 94556 311568
rect 160100 307776 160152 307828
rect 162124 307776 162176 307828
rect 221464 307708 221516 307760
rect 228364 307776 228416 307828
rect 3240 304988 3292 305040
rect 24124 304988 24176 305040
rect 51724 304988 51776 305040
rect 53104 304988 53156 305040
rect 157340 304988 157392 305040
rect 160100 304988 160152 305040
rect 155960 302268 156012 302320
rect 157340 302268 157392 302320
rect 46204 302200 46256 302252
rect 48964 302200 49016 302252
rect 155224 302200 155276 302252
rect 157984 302200 158036 302252
rect 57244 301452 57296 301504
rect 79324 301452 79376 301504
rect 61384 301044 61436 301096
rect 62764 301044 62816 301096
rect 556068 300840 556120 300892
rect 566556 300840 566608 300892
rect 66904 300160 66956 300212
rect 68284 300160 68336 300212
rect 220084 299412 220136 299464
rect 221464 299412 221516 299464
rect 552664 298732 552716 298784
rect 579988 298732 580040 298784
rect 152004 298528 152056 298580
rect 155868 298528 155920 298580
rect 150440 295944 150492 295996
rect 155224 295944 155276 295996
rect 151084 294040 151136 294092
rect 152004 294040 152056 294092
rect 3240 292544 3292 292596
rect 29736 292544 29788 292596
rect 146944 292544 146996 292596
rect 150440 292544 150492 292596
rect 91836 289756 91888 289808
rect 93124 289756 93176 289808
rect 55864 288328 55916 288380
rect 57244 288328 57296 288380
rect 556160 285608 556212 285660
rect 579988 285608 580040 285660
rect 135904 282140 135956 282192
rect 146944 282140 146996 282192
rect 60004 280780 60056 280832
rect 61384 280780 61436 280832
rect 88984 280100 89036 280152
rect 91836 280168 91888 280220
rect 218060 274728 218112 274780
rect 220084 274728 220136 274780
rect 57980 274660 58032 274712
rect 60004 274660 60056 274712
rect 45376 273164 45428 273216
rect 46204 273164 46256 273216
rect 54484 272892 54536 272944
rect 55864 272892 55916 272944
rect 397000 271872 397052 271924
rect 579988 271872 580040 271924
rect 215944 271056 215996 271108
rect 218060 271056 218112 271108
rect 52368 269084 52420 269136
rect 57888 269084 57940 269136
rect 149060 269016 149112 269068
rect 151084 269016 151136 269068
rect 51080 266364 51132 266416
rect 54484 266364 54536 266416
rect 63500 266364 63552 266416
rect 66904 266364 66956 266416
rect 146944 262896 146996 262948
rect 149060 262896 149112 262948
rect 50344 262828 50396 262880
rect 63500 262828 63552 262880
rect 121460 262828 121512 262880
rect 135904 262828 135956 262880
rect 50896 261196 50948 261248
rect 52368 261196 52420 261248
rect 47584 260448 47636 260500
rect 51080 260448 51132 260500
rect 49240 258952 49292 259004
rect 50896 258952 50948 259004
rect 81716 258680 81768 258732
rect 88984 258680 89036 258732
rect 117228 258680 117280 258732
rect 121460 258680 121512 258732
rect 397184 258068 397236 258120
rect 579988 258068 580040 258120
rect 47492 256708 47544 256760
rect 49240 256708 49292 256760
rect 210424 256640 210476 256692
rect 215944 256708 215996 256760
rect 3148 253920 3200 253972
rect 22744 253920 22796 253972
rect 45836 253920 45888 253972
rect 47492 253920 47544 253972
rect 79324 253920 79376 253972
rect 81716 253920 81768 253972
rect 113824 253920 113876 253972
rect 117228 253920 117280 253972
rect 145564 253920 145616 253972
rect 146944 253920 146996 253972
rect 209044 253920 209096 253972
rect 210424 253920 210476 253972
rect 48688 252560 48740 252612
rect 50344 252560 50396 252612
rect 47676 251812 47728 251864
rect 71780 251812 71832 251864
rect 46940 249432 46992 249484
rect 48688 249432 48740 249484
rect 97264 247664 97316 247716
rect 113824 247664 113876 247716
rect 76196 247052 76248 247104
rect 79324 247052 79376 247104
rect 143172 247052 143224 247104
rect 145564 247052 145616 247104
rect 49700 245624 49752 245676
rect 51724 245624 51776 245676
rect 413284 244264 413336 244316
rect 579988 244264 580040 244316
rect 136088 242836 136140 242888
rect 143172 242904 143224 242956
rect 45192 242224 45244 242276
rect 46940 242224 46992 242276
rect 45836 241408 45888 241460
rect 49608 241408 49660 241460
rect 45560 241340 45612 241392
rect 47676 241340 47728 241392
rect 45652 241272 45704 241324
rect 47584 241272 47636 241324
rect 46848 240864 46900 240916
rect 76196 240864 76248 240916
rect 45376 240796 45428 240848
rect 136088 240796 136140 240848
rect 45008 240728 45060 240780
rect 209044 240728 209096 240780
rect 3056 240116 3108 240168
rect 44824 240116 44876 240168
rect 395436 240048 395488 240100
rect 396540 240048 396592 240100
rect 44732 239708 44784 239760
rect 46848 239708 46900 239760
rect 45468 239368 45520 239420
rect 97264 239368 97316 239420
rect 396540 238824 396592 238876
rect 44916 238756 44968 238808
rect 45744 238756 45796 238808
rect 396540 238688 396592 238740
rect 44916 232908 44968 232960
rect 45836 232840 45888 232892
rect 45008 232772 45060 232824
rect 45744 232772 45796 232824
rect 64144 232364 64196 232416
rect 85764 232364 85816 232416
rect 394700 232092 394752 232144
rect 396540 232092 396592 232144
rect 45284 231888 45336 231940
rect 46848 231888 46900 231940
rect 45376 231820 45428 231872
rect 45468 231820 45520 231872
rect 46664 231820 46716 231872
rect 520924 231820 520976 231872
rect 579804 231820 579856 231872
rect 48320 231752 48372 231804
rect 45192 231072 45244 231124
rect 60740 231072 60792 231124
rect 85764 230664 85816 230716
rect 93768 230664 93820 230716
rect 390836 230460 390888 230512
rect 394700 230460 394752 230512
rect 45744 230392 45796 230444
rect 51908 230392 51960 230444
rect 60740 230120 60792 230172
rect 62764 230120 62816 230172
rect 167644 229712 167696 229764
rect 176660 229712 176712 229764
rect 48320 229100 48372 229152
rect 46664 229032 46716 229084
rect 48228 229032 48280 229084
rect 55864 229032 55916 229084
rect 157984 228420 158036 228472
rect 266544 228420 266596 228472
rect 297364 228420 297416 228472
rect 327080 228420 327132 228472
rect 366364 228420 366416 228472
rect 380164 228420 380216 228472
rect 117228 228352 117280 228404
rect 138664 228352 138716 228404
rect 236644 228352 236696 228404
rect 386512 228352 386564 228404
rect 51908 227740 51960 227792
rect 44732 227672 44784 227724
rect 46204 227672 46256 227724
rect 387064 227740 387116 227792
rect 392584 227740 392636 227792
rect 60004 227672 60056 227724
rect 64144 227060 64196 227112
rect 95884 227060 95936 227112
rect 3976 226992 4028 227044
rect 176660 226992 176712 227044
rect 93860 226448 93912 226500
rect 98000 226448 98052 226500
rect 384948 226244 385000 226296
rect 390836 226312 390888 226364
rect 46940 224340 46992 224392
rect 50344 224340 50396 224392
rect 55864 224136 55916 224188
rect 57244 224136 57296 224188
rect 60004 224136 60056 224188
rect 62120 224136 62172 224188
rect 98000 224136 98052 224188
rect 100024 224136 100076 224188
rect 380900 223524 380952 223576
rect 384948 223592 385000 223644
rect 46204 223252 46256 223304
rect 47676 223252 47728 223304
rect 48228 222096 48280 222148
rect 51448 222096 51500 222148
rect 62764 221416 62816 221468
rect 69020 221416 69072 221468
rect 372620 221416 372672 221468
rect 380900 221416 380952 221468
rect 62120 221212 62172 221264
rect 66260 221212 66312 221264
rect 45100 221076 45152 221128
rect 46940 221076 46992 221128
rect 369860 220396 369912 220448
rect 372620 220396 372672 220448
rect 69020 219444 69072 219496
rect 72424 219376 72476 219428
rect 95884 218696 95936 218748
rect 106188 218696 106240 218748
rect 379520 218696 379572 218748
rect 387064 218696 387116 218748
rect 47676 218016 47728 218068
rect 115848 218016 115900 218068
rect 579804 218016 579856 218068
rect 53840 217948 53892 218000
rect 100024 217948 100076 218000
rect 106004 217948 106056 218000
rect 45652 217268 45704 217320
rect 58256 217268 58308 217320
rect 46940 216656 46992 216708
rect 51724 216656 51776 216708
rect 66260 216656 66312 216708
rect 68284 216656 68336 216708
rect 366456 216588 366508 216640
rect 369860 216656 369912 216708
rect 57244 215772 57296 215824
rect 58716 215772 58768 215824
rect 106004 215296 106056 215348
rect 72424 215228 72476 215280
rect 75184 215228 75236 215280
rect 110420 215228 110472 215280
rect 106188 214616 106240 214668
rect 107844 214616 107896 214668
rect 3148 213936 3200 213988
rect 176752 213936 176804 213988
rect 51448 213868 51500 213920
rect 54484 213868 54536 213920
rect 58716 213868 58768 213920
rect 60004 213868 60056 213920
rect 58256 212440 58308 212492
rect 61936 212440 61988 212492
rect 375288 211896 375340 211948
rect 379428 211896 379480 211948
rect 53840 211148 53892 211200
rect 56692 211080 56744 211132
rect 110420 210468 110472 210520
rect 113180 210468 113232 210520
rect 107844 210400 107896 210452
rect 116584 210400 116636 210452
rect 371148 209788 371200 209840
rect 375288 209788 375340 209840
rect 382924 209040 382976 209092
rect 397552 209040 397604 209092
rect 54484 208156 54536 208208
rect 55864 208156 55916 208208
rect 56692 207748 56744 207800
rect 62028 207748 62080 207800
rect 60004 206932 60056 206984
rect 66168 206932 66220 206984
rect 113180 205980 113232 206032
rect 115112 205980 115164 206032
rect 364984 205708 365036 205760
rect 366456 205708 366508 205760
rect 188344 205640 188396 205692
rect 579988 205640 580040 205692
rect 61936 204892 61988 204944
rect 71044 204892 71096 204944
rect 367744 204756 367796 204808
rect 371148 204756 371200 204808
rect 62120 204212 62172 204264
rect 64144 204212 64196 204264
rect 75184 202852 75236 202904
rect 80704 202784 80756 202836
rect 2964 201492 3016 201544
rect 22836 201492 22888 201544
rect 362960 201492 363012 201544
rect 366364 201492 366416 201544
rect 115112 201424 115164 201476
rect 116860 201424 116912 201476
rect 51724 200744 51776 200796
rect 73160 200744 73212 200796
rect 66444 199384 66496 199436
rect 75460 199384 75512 199436
rect 155960 199384 156012 199436
rect 296720 199384 296772 199436
rect 377404 198704 377456 198756
rect 382924 198704 382976 198756
rect 362224 198024 362276 198076
rect 364984 198024 365036 198076
rect 50344 197956 50396 198008
rect 53840 197956 53892 198008
rect 73160 197956 73212 198008
rect 77944 197956 77996 198008
rect 148968 197956 149020 198008
rect 207020 197956 207072 198008
rect 116860 197820 116912 197872
rect 119988 197820 120040 197872
rect 154488 197412 154540 197464
rect 155960 197412 156012 197464
rect 68284 197344 68336 197396
rect 355324 197344 355376 197396
rect 362960 197344 363012 197396
rect 71780 197276 71832 197328
rect 152740 197276 152792 197328
rect 157984 197276 158036 197328
rect 147956 196732 148008 196784
rect 167644 196732 167696 196784
rect 160836 196664 160888 196716
rect 236644 196664 236696 196716
rect 151176 196596 151228 196648
rect 236000 196596 236052 196648
rect 64144 195916 64196 195968
rect 65524 195916 65576 195968
rect 138664 195916 138716 195968
rect 141424 195916 141476 195968
rect 157524 195916 157576 195968
rect 356060 195916 356112 195968
rect 86960 195848 87012 195900
rect 139400 195848 139452 195900
rect 157432 195848 157484 195900
rect 297364 195848 297416 195900
rect 56600 195780 56652 195832
rect 138112 195780 138164 195832
rect 71780 194488 71832 194540
rect 75184 194488 75236 194540
rect 75460 194488 75512 194540
rect 76564 194488 76616 194540
rect 116584 194488 116636 194540
rect 124864 194488 124916 194540
rect 217324 193808 217376 193860
rect 580172 193808 580224 193860
rect 53840 192448 53892 192500
rect 60372 192448 60424 192500
rect 120080 192448 120132 192500
rect 128360 192448 128412 192500
rect 341524 189728 341576 189780
rect 355324 189728 355376 189780
rect 60372 189048 60424 189100
rect 62764 189048 62816 189100
rect 128360 189048 128412 189100
rect 130384 189048 130436 189100
rect 359464 189048 359516 189100
rect 362224 189048 362276 189100
rect 76564 188572 76616 188624
rect 79968 188572 80020 188624
rect 80704 187892 80756 187944
rect 82176 187892 82228 187944
rect 3148 187688 3200 187740
rect 112444 187688 112496 187740
rect 366364 187688 366416 187740
rect 367744 187688 367796 187740
rect 166172 187620 166224 187672
rect 399484 187620 399536 187672
rect 79968 186328 80020 186380
rect 86224 186260 86276 186312
rect 159548 185852 159600 185904
rect 159916 185512 159968 185564
rect 135260 184152 135312 184204
rect 142436 184220 142488 184272
rect 371884 184152 371936 184204
rect 377404 184152 377456 184204
rect 82176 183472 82228 183524
rect 83556 183472 83608 183524
rect 65524 182112 65576 182164
rect 66904 182112 66956 182164
rect 144644 181500 144696 181552
rect 145196 181500 145248 181552
rect 157248 181160 157300 181212
rect 159916 181160 159968 181212
rect 144736 181092 144788 181144
rect 150900 181024 150952 181076
rect 157248 180616 157300 180668
rect 71044 180072 71096 180124
rect 81440 180072 81492 180124
rect 117320 180072 117372 180124
rect 136364 180072 136416 180124
rect 150900 180072 150952 180124
rect 153936 180072 153988 180124
rect 157248 180072 157300 180124
rect 62764 180004 62816 180056
rect 63776 180004 63828 180056
rect 158628 179596 158680 179648
rect 166540 179596 166592 179648
rect 154396 179528 154448 179580
rect 157800 179528 157852 179580
rect 130384 179392 130436 179444
rect 336556 179392 336608 179444
rect 341524 179392 341576 179444
rect 135168 179324 135220 179376
rect 136732 178780 136784 178832
rect 120724 178644 120776 178696
rect 136456 178644 136508 178696
rect 154396 178508 154448 178560
rect 157248 178508 157300 178560
rect 153108 178440 153160 178492
rect 153936 178440 153988 178492
rect 136364 178372 136416 178424
rect 114468 178032 114520 178084
rect 153936 178032 153988 178084
rect 154396 178032 154448 178084
rect 157800 178032 157852 178084
rect 158628 178032 158680 178084
rect 579988 178032 580040 178084
rect 63776 177964 63828 178016
rect 65524 177964 65576 178016
rect 134708 177760 134760 177812
rect 136640 177760 136692 177812
rect 120080 177284 120132 177336
rect 136456 177284 136508 177336
rect 144460 177216 144512 177268
rect 148048 177216 148100 177268
rect 55864 177148 55916 177200
rect 56876 177148 56928 177200
rect 368480 176672 368532 176724
rect 371884 176672 371936 176724
rect 83556 176604 83608 176656
rect 84936 176604 84988 176656
rect 153108 176400 153160 176452
rect 122840 176060 122892 176112
rect 134708 176060 134760 176112
rect 121460 175924 121512 175976
rect 136364 175924 136416 175976
rect 153108 175380 153160 175432
rect 141608 175312 141660 175364
rect 153936 175312 153988 175364
rect 56876 175244 56928 175296
rect 154396 175244 154448 175296
rect 156512 175244 156564 175296
rect 62120 175176 62172 175228
rect 81440 175176 81492 175228
rect 84844 175176 84896 175228
rect 153108 174836 153160 174888
rect 144092 174700 144144 174752
rect 145472 174700 145524 174752
rect 125600 174496 125652 174548
rect 136456 174496 136508 174548
rect 134524 174428 134576 174480
rect 329104 174632 329156 174684
rect 336556 174632 336608 174684
rect 364984 174632 365036 174684
rect 368480 174632 368532 174684
rect 140504 174360 140556 174412
rect 162492 174496 162544 174548
rect 145472 174428 145524 174480
rect 155500 174428 155552 174480
rect 115756 174292 115808 174344
rect 580448 174292 580500 174344
rect 129740 173884 129792 173936
rect 137376 173884 137428 173936
rect 155500 173884 155552 173936
rect 124864 173816 124916 173868
rect 128268 173816 128320 173868
rect 126980 173204 127032 173256
rect 136548 173204 136600 173256
rect 135168 173136 135220 173188
rect 62120 173000 62172 173052
rect 65248 173000 65300 173052
rect 159456 173000 159508 173052
rect 162860 172932 162912 172984
rect 143448 172864 143500 172916
rect 145656 172864 145708 172916
rect 146484 172864 146536 172916
rect 148600 172864 148652 172916
rect 156512 172864 156564 172916
rect 158444 172864 158496 172916
rect 143540 172796 143592 172848
rect 146668 172796 146720 172848
rect 142436 172728 142488 172780
rect 147588 172728 147640 172780
rect 45560 172456 45612 172508
rect 46940 172456 46992 172508
rect 133880 172116 133932 172168
rect 140780 172116 140832 172168
rect 131120 171844 131172 171896
rect 138664 171844 138716 171896
rect 132500 171504 132552 171556
rect 139676 171504 139728 171556
rect 128360 171096 128412 171148
rect 136732 171096 136784 171148
rect 140780 171096 140832 171148
rect 144920 171096 144972 171148
rect 84936 170076 84988 170128
rect 88248 170076 88300 170128
rect 162860 169668 162912 169720
rect 164976 169668 165028 169720
rect 46940 168988 46992 169040
rect 50988 168988 51040 169040
rect 362224 168512 362276 168564
rect 366364 168512 366416 168564
rect 84844 167628 84896 167680
rect 87696 167628 87748 167680
rect 88248 167016 88300 167068
rect 91100 166948 91152 167000
rect 164976 166268 165028 166320
rect 167644 166268 167696 166320
rect 359372 166268 359424 166320
rect 364984 166268 365036 166320
rect 185584 165588 185636 165640
rect 579804 165588 579856 165640
rect 65248 165520 65300 165572
rect 68284 165520 68336 165572
rect 86224 165520 86276 165572
rect 88984 165520 89036 165572
rect 65524 165452 65576 165504
rect 73804 165452 73856 165504
rect 128268 164840 128320 164892
rect 137284 164840 137336 164892
rect 87696 164160 87748 164212
rect 90364 164160 90416 164212
rect 91100 164160 91152 164212
rect 93124 164160 93176 164212
rect 314660 163480 314712 163532
rect 329104 163480 329156 163532
rect 3148 162868 3200 162920
rect 175372 162868 175424 162920
rect 50988 162120 51040 162172
rect 60556 162120 60608 162172
rect 338764 162120 338816 162172
rect 359372 162120 359424 162172
rect 167644 160080 167696 160132
rect 169024 160080 169076 160132
rect 360200 160080 360252 160132
rect 362224 160080 362276 160132
rect 147496 159264 147548 159316
rect 149704 159264 149756 159316
rect 60556 158992 60608 159044
rect 66996 158992 67048 159044
rect 73804 158652 73856 158704
rect 76748 158652 76800 158704
rect 309784 156544 309836 156596
rect 314660 156544 314712 156596
rect 76748 155932 76800 155984
rect 84844 155864 84896 155916
rect 129832 155864 129884 155916
rect 134524 155864 134576 155916
rect 356704 155864 356756 155916
rect 359464 155932 359516 155984
rect 137284 154504 137336 154556
rect 140688 154504 140740 154556
rect 357992 154164 358044 154216
rect 360200 154164 360252 154216
rect 84844 153212 84896 153264
rect 66996 153144 67048 153196
rect 71044 153144 71096 153196
rect 87604 153144 87656 153196
rect 127624 153144 127676 153196
rect 129832 153212 129884 153264
rect 93124 151784 93176 151836
rect 95240 151716 95292 151768
rect 88984 151512 89036 151564
rect 90456 151512 90508 151564
rect 77944 151036 77996 151088
rect 81440 151036 81492 151088
rect 169024 149676 169076 149728
rect 170128 149676 170180 149728
rect 3148 149064 3200 149116
rect 25504 149064 25556 149116
rect 307668 149064 307720 149116
rect 309784 149064 309836 149116
rect 140688 148316 140740 148368
rect 162124 148316 162176 148368
rect 170128 147568 170180 147620
rect 172428 147568 172480 147620
rect 68284 146208 68336 146260
rect 69664 146208 69716 146260
rect 95240 146208 95292 146260
rect 97264 146208 97316 146260
rect 149704 146208 149756 146260
rect 152648 146208 152700 146260
rect 81440 145528 81492 145580
rect 91744 145528 91796 145580
rect 351920 145528 351972 145580
rect 357992 145528 358044 145580
rect 303620 143556 303672 143608
rect 307668 143556 307720 143608
rect 69664 143488 69716 143540
rect 71136 143488 71188 143540
rect 75184 143488 75236 143540
rect 76564 143488 76616 143540
rect 152648 143488 152700 143540
rect 154856 143488 154908 143540
rect 347044 143488 347096 143540
rect 351920 143556 351972 143608
rect 71044 143012 71096 143064
rect 76656 143012 76708 143064
rect 115664 142808 115716 142860
rect 580540 142808 580592 142860
rect 91744 141516 91796 141568
rect 94044 141516 94096 141568
rect 66904 141244 66956 141296
rect 68376 141244 68428 141296
rect 172520 138388 172572 138440
rect 174360 138388 174412 138440
rect 3424 138320 3476 138372
rect 4068 138320 4120 138372
rect 300860 138048 300912 138100
rect 303620 138048 303672 138100
rect 90364 137980 90416 138032
rect 93124 137980 93176 138032
rect 114376 137980 114428 138032
rect 579988 137980 580040 138032
rect 90456 137912 90508 137964
rect 94688 137912 94740 137964
rect 119344 137912 119396 137964
rect 120724 137912 120776 137964
rect 142436 137912 142488 137964
rect 145932 137912 145984 137964
rect 150532 137912 150584 137964
rect 152188 137912 152240 137964
rect 164516 137912 164568 137964
rect 172520 137912 172572 137964
rect 68376 137844 68428 137896
rect 69664 137844 69716 137896
rect 154856 137708 154908 137760
rect 164700 137708 164752 137760
rect 144460 137640 144512 137692
rect 156880 137640 156932 137692
rect 163504 137640 163556 137692
rect 174084 137640 174136 137692
rect 114100 137572 114152 137624
rect 396908 137572 396960 137624
rect 114192 137504 114244 137556
rect 397092 137504 397144 137556
rect 114284 137436 114336 137488
rect 397184 137436 397236 137488
rect 113824 137368 113876 137420
rect 412640 137368 412692 137420
rect 115112 137300 115164 137352
rect 477500 137300 477552 137352
rect 115388 137232 115440 137284
rect 580632 137232 580684 137284
rect 152464 137164 152516 137216
rect 153752 137164 153804 137216
rect 163596 136756 163648 136808
rect 170956 136756 171008 136808
rect 138112 136688 138164 136740
rect 142528 136688 142580 136740
rect 153476 136688 153528 136740
rect 155316 136688 155368 136740
rect 3424 136620 3476 136672
rect 115204 136620 115256 136672
rect 174360 136552 174412 136604
rect 176016 136552 176068 136604
rect 162124 136484 162176 136536
rect 175924 136484 175976 136536
rect 40040 136416 40092 136468
rect 176844 136416 176896 136468
rect 3976 136348 4028 136400
rect 178132 136348 178184 136400
rect 3792 136280 3844 136332
rect 178592 136280 178644 136332
rect 3884 136212 3936 136264
rect 178408 136212 178460 136264
rect 3700 136144 3752 136196
rect 178776 136144 178828 136196
rect 3240 136076 3292 136128
rect 178040 136076 178092 136128
rect 3332 136008 3384 136060
rect 178500 136008 178552 136060
rect 295340 136008 295392 136060
rect 300860 136008 300912 136060
rect 115480 135940 115532 135992
rect 580816 135940 580868 135992
rect 94044 135872 94096 135924
rect 105544 135872 105596 135924
rect 113916 135872 113968 135924
rect 580080 135872 580132 135924
rect 71136 135192 71188 135244
rect 72424 135192 72476 135244
rect 115572 134784 115624 134836
rect 127624 134784 127676 134836
rect 87604 134716 87656 134768
rect 177304 134716 177356 134768
rect 3608 134648 3660 134700
rect 178316 134648 178368 134700
rect 4068 134580 4120 134632
rect 178684 134580 178736 134632
rect 113732 134512 113784 134564
rect 295340 134512 295392 134564
rect 3792 133900 3844 133952
rect 175372 133900 175424 133952
rect 94688 133832 94740 133884
rect 95608 133832 95660 133884
rect 76656 133152 76708 133204
rect 86224 133152 86276 133204
rect 115112 132676 115164 132728
rect 115296 132676 115348 132728
rect 95608 131724 95660 131776
rect 97540 131724 97592 131776
rect 97264 131588 97316 131640
rect 99288 131588 99340 131640
rect 3424 131112 3476 131164
rect 113640 131112 113692 131164
rect 3608 128324 3660 128376
rect 113548 128324 113600 128376
rect 93124 128256 93176 128308
rect 95884 128256 95936 128308
rect 76564 127576 76616 127628
rect 79324 127576 79376 127628
rect 105544 127576 105596 127628
rect 111064 127576 111116 127628
rect 3700 126964 3752 127016
rect 113548 126964 113600 127016
rect 25504 126896 25556 126948
rect 113640 126896 113692 126948
rect 99380 126828 99432 126880
rect 101496 126828 101548 126880
rect 184204 125604 184256 125656
rect 580080 125604 580132 125656
rect 22836 125536 22888 125588
rect 113640 125536 113692 125588
rect 350724 124176 350776 124228
rect 356704 124176 356756 124228
rect 22744 124108 22796 124160
rect 113640 124108 113692 124160
rect 97540 124040 97592 124092
rect 99288 124040 99340 124092
rect 24124 122748 24176 122800
rect 113640 122748 113692 122800
rect 72424 121456 72476 121508
rect 73804 121456 73856 121508
rect 86224 121456 86276 121508
rect 88984 121456 89036 121508
rect 345756 121456 345808 121508
rect 347044 121456 347096 121508
rect 347872 121456 347924 121508
rect 350724 121456 350776 121508
rect 10324 121388 10376 121440
rect 113640 121388 113692 121440
rect 101496 121320 101548 121372
rect 104900 121320 104952 121372
rect 99380 121252 99432 121304
rect 102048 121252 102100 121304
rect 8944 120028 8996 120080
rect 113640 120028 113692 120080
rect 69664 119960 69716 120012
rect 70492 119960 70544 120012
rect 104900 119620 104952 119672
rect 106924 119620 106976 119672
rect 5080 118600 5132 118652
rect 113640 118600 113692 118652
rect 70492 118532 70544 118584
rect 76288 118532 76340 118584
rect 177304 118532 177356 118584
rect 178224 118532 178276 118584
rect 79324 118260 79376 118312
rect 81164 118260 81216 118312
rect 342260 118192 342312 118244
rect 345756 118192 345808 118244
rect 343640 117920 343692 117972
rect 347872 117920 347924 117972
rect 33784 117240 33836 117292
rect 113640 117240 113692 117292
rect 176016 117240 176068 117292
rect 176660 117240 176712 117292
rect 76288 116016 76340 116068
rect 77944 116016 77996 116068
rect 29644 115880 29696 115932
rect 113548 115880 113600 115932
rect 81164 114452 81216 114504
rect 82820 114452 82872 114504
rect 340420 114452 340472 114504
rect 342260 114520 342312 114572
rect 341524 113704 341576 113756
rect 343640 113704 343692 113756
rect 37924 113092 37976 113144
rect 113640 113092 113692 113144
rect 95884 112412 95936 112464
rect 108304 112412 108356 112464
rect 333980 112412 334032 112464
rect 340420 112412 340472 112464
rect 77944 112276 77996 112328
rect 79968 112276 80020 112328
rect 15844 111732 15896 111784
rect 113640 111732 113692 111784
rect 82820 111052 82872 111104
rect 88248 111052 88300 111104
rect 324320 111052 324372 111104
rect 333980 111052 334032 111104
rect 23480 110372 23532 110424
rect 113640 110372 113692 110424
rect 108304 108944 108356 108996
rect 113640 108944 113692 108996
rect 80060 107584 80112 107636
rect 113640 107584 113692 107636
rect 102140 107516 102192 107568
rect 106188 107516 106240 107568
rect 106188 106224 106240 106276
rect 113548 106224 113600 106276
rect 178040 106224 178092 106276
rect 341524 106224 341576 106276
rect 88248 104864 88300 104916
rect 113640 104796 113692 104848
rect 178040 104796 178092 104848
rect 324228 104796 324280 104848
rect 106924 104728 106976 104780
rect 108396 104728 108448 104780
rect 88984 103844 89036 103896
rect 95240 103844 95292 103896
rect 178040 103436 178092 103488
rect 410524 103436 410576 103488
rect 178040 102076 178092 102128
rect 409144 102076 409196 102128
rect 178040 100648 178092 100700
rect 407764 100648 407816 100700
rect 175924 99356 175976 99408
rect 580080 99356 580132 99408
rect 178040 99288 178092 99340
rect 566464 99288 566516 99340
rect 95240 98676 95292 98728
rect 98644 98676 98696 98728
rect 73804 98608 73856 98660
rect 77944 98608 77996 98660
rect 178040 97928 178092 97980
rect 406384 97928 406436 97980
rect 108396 96636 108448 96688
rect 110972 96568 111024 96620
rect 178040 95140 178092 95192
rect 405004 95140 405056 95192
rect 178040 93780 178092 93832
rect 403624 93780 403676 93832
rect 178040 92420 178092 92472
rect 400864 92420 400916 92472
rect 320824 91740 320876 91792
rect 338764 91740 338816 91792
rect 178040 90992 178092 91044
rect 417424 90992 417476 91044
rect 178040 89632 178092 89684
rect 414664 89632 414716 89684
rect 110972 88272 111024 88324
rect 113824 88272 113876 88324
rect 178040 88272 178092 88324
rect 552664 88272 552716 88324
rect 77944 86980 77996 87032
rect 83556 86912 83608 86964
rect 178040 86912 178092 86964
rect 413284 86912 413336 86964
rect 179236 85552 179288 85604
rect 580080 85552 580132 85604
rect 178040 85484 178092 85536
rect 188344 85484 188396 85536
rect 307760 84804 307812 84856
rect 320824 84804 320876 84856
rect 3332 84192 3384 84244
rect 116584 84192 116636 84244
rect 178040 84124 178092 84176
rect 185584 84124 185636 84176
rect 98644 82832 98696 82884
rect 104164 82832 104216 82884
rect 178040 82764 178092 82816
rect 184204 82764 184256 82816
rect 113824 81608 113876 81660
rect 114560 81608 114612 81660
rect 83556 79976 83608 80028
rect 84844 79976 84896 80028
rect 299388 77936 299440 77988
rect 307760 77936 307812 77988
rect 178040 75896 178092 75948
rect 562324 75896 562376 75948
rect 114468 75692 114520 75744
rect 175924 75692 175976 75744
rect 114560 75624 114612 75676
rect 118608 75624 118660 75676
rect 170680 75624 170732 75676
rect 29736 75216 29788 75268
rect 172244 75284 172296 75336
rect 141792 74876 141844 74928
rect 170404 75216 170456 75268
rect 150624 74876 150676 74928
rect 145104 74808 145156 74860
rect 164424 74876 164476 74928
rect 170496 75148 170548 75200
rect 170588 75080 170640 75132
rect 175372 75148 175424 75200
rect 299388 75148 299440 75200
rect 259460 75080 259512 75132
rect 170864 75012 170916 75064
rect 195980 75012 196032 75064
rect 170404 74944 170456 74996
rect 302240 74944 302292 74996
rect 165068 74876 165120 74928
rect 146760 74672 146812 74724
rect 168104 74740 168156 74792
rect 153384 74400 153436 74452
rect 168104 74604 168156 74656
rect 169392 74604 169444 74656
rect 169760 74876 169812 74928
rect 170772 74876 170824 74928
rect 324320 74876 324372 74928
rect 170680 74808 170732 74860
rect 172244 74808 172296 74860
rect 374000 74808 374052 74860
rect 172152 74740 172204 74792
rect 396724 74740 396776 74792
rect 170404 74672 170456 74724
rect 170680 74604 170732 74656
rect 172060 74672 172112 74724
rect 396816 74672 396868 74724
rect 462412 74604 462464 74656
rect 164424 74536 164476 74588
rect 170404 74536 170456 74588
rect 170496 74536 170548 74588
rect 550640 74536 550692 74588
rect 161664 74468 161716 74520
rect 167644 74468 167696 74520
rect 168564 74468 168616 74520
rect 175372 74468 175424 74520
rect 167092 74400 167144 74452
rect 580540 74468 580592 74520
rect 111064 74332 111116 74384
rect 113916 74332 113968 74384
rect 157524 74332 157576 74384
rect 164424 74332 164476 74384
rect 167184 74332 167236 74384
rect 580448 74400 580500 74452
rect 115204 74264 115256 74316
rect 170036 74264 170088 74316
rect 140964 74196 141016 74248
rect 249800 74196 249852 74248
rect 143724 74128 143776 74180
rect 284300 74128 284352 74180
rect 146484 74060 146536 74112
rect 320180 74060 320232 74112
rect 147864 73992 147916 74044
rect 338120 73992 338172 74044
rect 152004 73924 152056 73976
rect 390560 73924 390612 73976
rect 116584 73856 116636 73908
rect 157800 73788 157852 73840
rect 161664 73788 161716 73840
rect 112444 73720 112496 73772
rect 168380 73856 168432 73908
rect 462320 73856 462372 73908
rect 164424 73788 164476 73840
rect 465172 73788 465224 73840
rect 5264 73652 5316 73704
rect 170128 73720 170180 73772
rect 44824 73584 44876 73636
rect 169944 73652 169996 73704
rect 167736 73584 167788 73636
rect 172152 73584 172204 73636
rect 161664 73516 161716 73568
rect 167460 73516 167512 73568
rect 167552 73516 167604 73568
rect 172060 73516 172112 73568
rect 169668 73448 169720 73500
rect 169852 73380 169904 73432
rect 152004 73312 152056 73364
rect 152188 73312 152240 73364
rect 84844 73176 84896 73228
rect 152188 73176 152240 73228
rect 152740 73176 152792 73228
rect 162400 73244 162452 73296
rect 92480 73108 92532 73160
rect 118608 73108 118660 73160
rect 120080 73108 120132 73160
rect 120908 73108 120960 73160
rect 127900 73108 127952 73160
rect 136824 73108 136876 73160
rect 161664 73108 161716 73160
rect 137652 73040 137704 73092
rect 207020 73176 207072 73228
rect 164424 73108 164476 73160
rect 166724 73108 166776 73160
rect 172888 73108 172940 73160
rect 165068 73040 165120 73092
rect 167736 73040 167788 73092
rect 167828 73040 167880 73092
rect 580724 73040 580776 73092
rect 120724 72972 120776 73024
rect 128176 72972 128228 73024
rect 136272 72972 136324 73024
rect 168104 72972 168156 73024
rect 168472 72972 168524 73024
rect 397460 72972 397512 73024
rect 120816 72904 120868 72956
rect 129280 72904 129332 72956
rect 141608 72904 141660 72956
rect 146760 72904 146812 72956
rect 154396 72904 154448 72956
rect 422300 72904 422352 72956
rect 121092 72836 121144 72888
rect 130384 72836 130436 72888
rect 142160 72836 142212 72888
rect 152740 72836 152792 72888
rect 156052 72836 156104 72888
rect 443000 72836 443052 72888
rect 149152 72768 149204 72820
rect 154396 72768 154448 72820
rect 156604 72768 156656 72820
rect 449900 72768 449952 72820
rect 121000 72700 121052 72752
rect 129832 72700 129884 72752
rect 140504 72700 140556 72752
rect 151636 72700 151688 72752
rect 152004 72700 152056 72752
rect 121368 72632 121420 72684
rect 132684 72632 132736 72684
rect 138848 72632 138900 72684
rect 146484 72632 146536 72684
rect 150256 72632 150308 72684
rect 132316 72564 132368 72616
rect 137744 72564 137796 72616
rect 139216 72564 139268 72616
rect 60740 72496 60792 72548
rect 126336 72496 126388 72548
rect 134708 72496 134760 72548
rect 149152 72496 149204 72548
rect 151268 72564 151320 72616
rect 154212 72564 154264 72616
rect 153108 72496 153160 72548
rect 157432 72700 157484 72752
rect 158812 72700 158864 72752
rect 158260 72632 158312 72684
rect 164424 72700 164476 72752
rect 166356 72700 166408 72752
rect 167736 72700 167788 72752
rect 460940 72700 460992 72752
rect 471980 72632 472032 72684
rect 158260 72496 158312 72548
rect 25504 72428 25556 72480
rect 123116 72428 123168 72480
rect 135720 72428 135772 72480
rect 116584 72360 116636 72412
rect 124864 72360 124916 72412
rect 137652 72360 137704 72412
rect 118148 72292 118200 72344
rect 124312 72292 124364 72344
rect 86224 72224 86276 72276
rect 122380 72224 122432 72276
rect 117964 72156 118016 72208
rect 123760 72156 123812 72208
rect 118056 72088 118108 72140
rect 123024 72088 123076 72140
rect 157524 72428 157576 72480
rect 150808 72360 150860 72412
rect 152924 72360 152976 72412
rect 162492 72564 162544 72616
rect 514760 72564 514812 72616
rect 158812 72496 158864 72548
rect 165068 72496 165120 72548
rect 170588 72496 170640 72548
rect 558920 72496 558972 72548
rect 166632 72428 166684 72480
rect 581000 72428 581052 72480
rect 167368 72360 167420 72412
rect 167920 72360 167972 72412
rect 217324 72360 217376 72412
rect 152188 72292 152240 72344
rect 167460 72292 167512 72344
rect 145472 72224 145524 72276
rect 146484 72156 146536 72208
rect 150164 72156 150216 72208
rect 153844 72224 153896 72276
rect 168288 72224 168340 72276
rect 154396 72156 154448 72208
rect 142712 72088 142764 72140
rect 146024 72020 146076 72072
rect 154948 72088 155000 72140
rect 167736 72156 167788 72208
rect 153016 72020 153068 72072
rect 153292 72020 153344 72072
rect 167552 72088 167604 72140
rect 151912 71952 151964 72004
rect 155776 71952 155828 72004
rect 146760 71884 146812 71936
rect 151544 71884 151596 71936
rect 151820 71884 151872 71936
rect 157156 71884 157208 71936
rect 157524 71884 157576 71936
rect 165252 71884 165304 71936
rect 119344 71816 119396 71868
rect 122748 71816 122800 71868
rect 132500 71816 132552 71868
rect 136272 71816 136324 71868
rect 136640 71816 136692 71868
rect 122380 71748 122432 71800
rect 127348 71748 127400 71800
rect 133972 71748 134024 71800
rect 137652 71748 137704 71800
rect 151360 71816 151412 71868
rect 158444 71816 158496 71868
rect 143172 71748 143224 71800
rect 145840 71748 145892 71800
rect 147312 71748 147364 71800
rect 149704 71748 149756 71800
rect 156972 71748 157024 71800
rect 3516 71680 3568 71732
rect 178868 72020 178920 72072
rect 167092 71952 167144 72004
rect 580172 71952 580224 72004
rect 6920 71612 6972 71664
rect 169024 71612 169076 71664
rect 92480 71544 92532 71596
rect 168656 71544 168708 71596
rect 104164 71476 104216 71528
rect 168932 71476 168984 71528
rect 113916 71408 113968 71460
rect 168748 71408 168800 71460
rect 120080 71340 120132 71392
rect 168840 71340 168892 71392
rect 166908 71000 166960 71052
rect 580264 71000 580316 71052
rect 122932 70048 122984 70100
rect 124128 70048 124180 70100
rect 131212 70048 131264 70100
rect 131580 70048 131632 70100
rect 121552 69980 121604 70032
rect 122564 69980 122616 70032
rect 123024 69980 123076 70032
rect 123852 69980 123904 70032
rect 124312 69980 124364 70032
rect 125232 69980 125284 70032
rect 128544 69980 128596 70032
rect 129372 69980 129424 70032
rect 123208 69912 123260 69964
rect 123668 69912 123720 69964
rect 129188 69912 129240 69964
rect 130108 69912 130160 69964
rect 130384 69912 130436 69964
rect 121460 69844 121512 69896
rect 122012 69844 122064 69896
rect 122104 69844 122156 69896
rect 122564 69844 122616 69896
rect 123576 69844 123628 69896
rect 124128 69844 124180 69896
rect 124588 69844 124640 69896
rect 125232 69844 125284 69896
rect 121736 69776 121788 69828
rect 122196 69776 122248 69828
rect 123944 69776 123996 69828
rect 124496 69776 124548 69828
rect 124956 69776 125008 69828
rect 127072 69776 127124 69828
rect 127716 69776 127768 69828
rect 125692 69708 125744 69760
rect 126612 69708 126664 69760
rect 130476 69776 130528 69828
rect 138112 69776 138164 69828
rect 138848 69776 138900 69828
rect 130016 69708 130068 69760
rect 125784 69640 125836 69692
rect 126428 69640 126480 69692
rect 129188 69640 129240 69692
rect 130476 69640 130528 69692
rect 130936 69640 130988 69692
rect 131120 69640 131172 69692
rect 131764 69640 131816 69692
rect 122104 69572 122156 69624
rect 122656 69572 122708 69624
rect 123484 69572 123536 69624
rect 127164 69572 127216 69624
rect 127440 69572 127492 69624
rect 128820 69572 128872 69624
rect 129280 69572 129332 69624
rect 130200 69572 130252 69624
rect 130568 69572 130620 69624
rect 123116 69504 123168 69556
rect 123760 69504 123812 69556
rect 127348 69504 127400 69556
rect 127624 69504 127676 69556
rect 130108 69504 130160 69556
rect 130844 69504 130896 69556
rect 131304 69504 131356 69556
rect 124864 69436 124916 69488
rect 125416 69436 125468 69488
rect 131580 69368 131632 69420
rect 126428 69300 126480 69352
rect 126796 69300 126848 69352
rect 127440 69300 127492 69352
rect 127900 69300 127952 69352
rect 131396 69300 131448 69352
rect 127348 69232 127400 69284
rect 128268 69232 128320 69284
rect 126060 69164 126112 69216
rect 126520 69164 126572 69216
rect 131580 69164 131632 69216
rect 127716 69096 127768 69148
rect 128084 69096 128136 69148
rect 121644 68212 121696 68264
rect 122288 68212 122340 68264
rect 125968 67804 126020 67856
rect 126244 67804 126296 67856
rect 129924 67600 129976 67652
rect 130752 67600 130804 67652
rect 125784 67532 125836 67584
rect 125968 67532 126020 67584
rect 126060 67532 126112 67584
rect 126704 67532 126756 67584
rect 124680 67328 124732 67380
rect 125324 67328 125376 67380
rect 5540 66852 5592 66904
rect 121460 66852 121512 66904
rect 124772 65900 124824 65952
rect 125048 65900 125100 65952
rect 128820 65628 128872 65680
rect 129464 65628 129516 65680
rect 128912 65560 128964 65612
rect 129188 65560 129240 65612
rect 129096 65492 129148 65544
rect 129556 65492 129608 65544
rect 128636 65424 128688 65476
rect 129188 65424 129240 65476
rect 128636 65288 128688 65340
rect 129648 65288 129700 65340
rect 114376 60664 114428 60716
rect 580172 60664 580224 60716
rect 163504 58624 163556 58676
rect 326344 58624 326396 58676
rect 15200 54476 15252 54528
rect 119344 54476 119396 54528
rect 113180 51076 113232 51128
rect 121092 51076 121144 51128
rect 178684 46860 178736 46912
rect 580172 46860 580224 46912
rect 3516 45500 3568 45552
rect 170220 45500 170272 45552
rect 106280 43392 106332 43444
rect 121000 43392 121052 43444
rect 153108 40672 153160 40724
rect 226340 40672 226392 40724
rect 158444 36660 158496 36712
rect 382280 36660 382332 36712
rect 155776 36592 155828 36644
rect 390652 36592 390704 36644
rect 152464 36524 152516 36576
rect 397460 36524 397512 36576
rect 145564 35844 145616 35896
rect 307760 35844 307812 35896
rect 147312 35776 147364 35828
rect 311900 35776 311952 35828
rect 146392 35708 146444 35760
rect 318800 35708 318852 35760
rect 146668 35640 146720 35692
rect 322940 35640 322992 35692
rect 146944 35572 146996 35624
rect 325700 35572 325752 35624
rect 147772 35504 147824 35556
rect 336740 35504 336792 35556
rect 148600 35436 148652 35488
rect 347780 35436 347832 35488
rect 154488 35368 154540 35420
rect 354680 35368 354732 35420
rect 149428 35300 149480 35352
rect 357440 35300 357492 35352
rect 158352 35232 158404 35284
rect 368480 35232 368532 35284
rect 157800 35164 157852 35216
rect 456800 35164 456852 35216
rect 145288 35096 145340 35148
rect 305000 35096 305052 35148
rect 138848 34416 138900 34468
rect 212540 34416 212592 34468
rect 138388 34348 138440 34400
rect 216680 34348 216732 34400
rect 138664 34280 138716 34332
rect 219440 34280 219492 34332
rect 139768 34212 139820 34264
rect 234620 34212 234672 34264
rect 140872 34144 140924 34196
rect 248420 34144 248472 34196
rect 141424 34076 141476 34128
rect 255320 34076 255372 34128
rect 142528 34008 142580 34060
rect 269120 34008 269172 34060
rect 143080 33940 143132 33992
rect 276020 33940 276072 33992
rect 143632 33872 143684 33924
rect 284392 33872 284444 33924
rect 144184 33804 144236 33856
rect 291200 33804 291252 33856
rect 145012 33736 145064 33788
rect 300860 33736 300912 33788
rect 2872 33056 2924 33108
rect 175280 33056 175332 33108
rect 135352 32920 135404 32972
rect 176660 32920 176712 32972
rect 135628 32852 135680 32904
rect 180800 32852 180852 32904
rect 135904 32784 135956 32836
rect 184940 32784 184992 32836
rect 136732 32716 136784 32768
rect 194600 32716 194652 32768
rect 137008 32648 137060 32700
rect 198740 32648 198792 32700
rect 137560 32580 137612 32632
rect 205640 32580 205692 32632
rect 142252 32512 142304 32564
rect 266360 32512 266412 32564
rect 164332 32444 164384 32496
rect 549260 32444 549312 32496
rect 166264 32376 166316 32428
rect 574100 32376 574152 32428
rect 157616 31696 157668 31748
rect 463700 31696 463752 31748
rect 158168 31628 158220 31680
rect 470600 31628 470652 31680
rect 158720 31560 158772 31612
rect 477500 31560 477552 31612
rect 159088 31492 159140 31544
rect 481640 31492 481692 31544
rect 161112 31424 161164 31476
rect 490012 31424 490064 31476
rect 160192 31356 160244 31408
rect 496820 31356 496872 31408
rect 160744 31288 160796 31340
rect 503720 31288 503772 31340
rect 162584 31220 162636 31272
rect 510620 31220 510672 31272
rect 161848 31152 161900 31204
rect 517520 31152 517572 31204
rect 166356 31084 166408 31136
rect 524420 31084 524472 31136
rect 162124 31016 162176 31068
rect 521660 31016 521712 31068
rect 154304 30268 154356 30320
rect 307852 30268 307904 30320
rect 144920 30200 144972 30252
rect 299480 30200 299532 30252
rect 145196 30132 145248 30184
rect 303620 30132 303672 30184
rect 150716 30064 150768 30116
rect 374092 30064 374144 30116
rect 154212 29996 154264 30048
rect 382372 29996 382424 30048
rect 157248 29928 157300 29980
rect 389180 29928 389232 29980
rect 155132 29860 155184 29912
rect 431960 29860 432012 29912
rect 157064 29792 157116 29844
rect 438860 29792 438912 29844
rect 155960 29724 156012 29776
rect 441620 29724 441672 29776
rect 156236 29656 156288 29708
rect 445760 29656 445812 29708
rect 156788 29588 156840 29640
rect 452660 29588 452712 29640
rect 139400 28908 139452 28960
rect 229100 28908 229152 28960
rect 151636 28840 151688 28892
rect 242900 28840 242952 28892
rect 140228 28772 140280 28824
rect 240140 28772 240192 28824
rect 140780 28704 140832 28756
rect 247040 28704 247092 28756
rect 151544 28636 151596 28688
rect 258080 28636 258132 28688
rect 141056 28568 141108 28620
rect 251180 28568 251232 28620
rect 152832 28500 152884 28552
rect 264980 28500 265032 28552
rect 153016 28432 153068 28484
rect 271880 28432 271932 28484
rect 150440 28364 150492 28416
rect 371240 28364 371292 28416
rect 152924 28296 152976 28348
rect 375380 28296 375432 28348
rect 165988 28228 166040 28280
rect 571340 28228 571392 28280
rect 138296 28160 138348 28212
rect 215300 28160 215352 28212
rect 138112 28092 138164 28144
rect 211160 28092 211212 28144
rect 150164 28024 150216 28076
rect 222200 28024 222252 28076
rect 143172 27548 143224 27600
rect 193220 27548 193272 27600
rect 136088 27480 136140 27532
rect 186320 27480 186372 27532
rect 136916 27412 136968 27464
rect 197360 27412 197412 27464
rect 146024 27344 146076 27396
rect 208400 27344 208452 27396
rect 137192 27276 137244 27328
rect 201500 27276 201552 27328
rect 137468 27208 137520 27260
rect 204260 27208 204312 27260
rect 138572 27140 138624 27192
rect 218060 27140 218112 27192
rect 139676 27072 139728 27124
rect 233240 27072 233292 27124
rect 148324 27004 148376 27056
rect 343640 27004 343692 27056
rect 154580 26936 154632 26988
rect 423680 26936 423732 26988
rect 157984 26868 158036 26920
rect 467840 26868 467892 26920
rect 135536 26188 135588 26240
rect 179420 26188 179472 26240
rect 135812 26120 135864 26172
rect 183560 26120 183612 26172
rect 139952 26052 140004 26104
rect 236000 26052 236052 26104
rect 141884 25984 141936 26036
rect 260840 25984 260892 26036
rect 144368 25916 144420 25968
rect 292580 25916 292632 25968
rect 149336 25848 149388 25900
rect 357532 25848 357584 25900
rect 150532 25780 150584 25832
rect 372620 25780 372672 25832
rect 153752 25712 153804 25764
rect 414020 25712 414072 25764
rect 164792 25644 164844 25696
rect 556160 25644 556212 25696
rect 165620 25576 165672 25628
rect 565820 25576 565872 25628
rect 81440 25508 81492 25560
rect 120908 25508 120960 25560
rect 166172 25508 166224 25560
rect 572720 25508 572772 25560
rect 135260 25440 135312 25492
rect 176752 25440 176804 25492
rect 141332 24760 141384 24812
rect 253940 24760 253992 24812
rect 143540 24692 143592 24744
rect 282920 24692 282972 24744
rect 153200 24624 153252 24676
rect 407212 24624 407264 24676
rect 162860 24556 162912 24608
rect 531320 24556 531372 24608
rect 163136 24488 163188 24540
rect 534080 24488 534132 24540
rect 163412 24420 163464 24472
rect 538220 24420 538272 24472
rect 163688 24352 163740 24404
rect 540980 24352 541032 24404
rect 164240 24284 164292 24336
rect 547880 24284 547932 24336
rect 164516 24216 164568 24268
rect 552020 24216 552072 24268
rect 165712 24148 165764 24200
rect 567200 24148 567252 24200
rect 165896 24080 165948 24132
rect 569960 24080 570012 24132
rect 157340 23400 157392 23452
rect 459560 23400 459612 23452
rect 160100 23332 160152 23384
rect 495440 23332 495492 23384
rect 160376 23264 160428 23316
rect 498292 23264 498344 23316
rect 160652 23196 160704 23248
rect 502340 23196 502392 23248
rect 160928 23128 160980 23180
rect 506480 23128 506532 23180
rect 161480 23060 161532 23112
rect 513380 23060 513432 23112
rect 161756 22992 161808 23044
rect 516140 22992 516192 23044
rect 162032 22924 162084 22976
rect 520280 22924 520332 22976
rect 162308 22856 162360 22908
rect 523040 22856 523092 22908
rect 165160 22788 165212 22840
rect 560300 22788 560352 22840
rect 114468 22720 114520 22772
rect 580172 22720 580224 22772
rect 3516 22652 3568 22704
rect 170312 22652 170364 22704
rect 148048 22040 148100 22092
rect 340880 22040 340932 22092
rect 156972 21972 157024 22024
rect 361580 21972 361632 22024
rect 154672 21904 154724 21956
rect 425060 21904 425112 21956
rect 155040 21836 155092 21888
rect 430580 21836 430632 21888
rect 155224 21768 155276 21820
rect 432052 21768 432104 21820
rect 156328 21700 156380 21752
rect 447140 21700 447192 21752
rect 156420 21632 156472 21684
rect 448520 21632 448572 21684
rect 158996 21564 159048 21616
rect 481732 21564 481784 21616
rect 159272 21496 159324 21548
rect 484400 21496 484452 21548
rect 159548 21428 159600 21480
rect 488540 21428 488592 21480
rect 159824 21360 159876 21412
rect 491300 21360 491352 21412
rect 139492 20408 139544 20460
rect 230480 20408 230532 20460
rect 140044 20340 140096 20392
rect 237380 20340 237432 20392
rect 141700 20272 141752 20324
rect 259552 20272 259604 20324
rect 147220 20204 147272 20256
rect 329840 20204 329892 20256
rect 152280 20136 152332 20188
rect 394700 20136 394752 20188
rect 152556 20068 152608 20120
rect 398840 20068 398892 20120
rect 153660 20000 153712 20052
rect 412640 20000 412692 20052
rect 158076 19932 158128 19984
rect 469220 19932 469272 19984
rect 141148 19048 141200 19100
rect 251272 19048 251324 19100
rect 163780 18980 163832 19032
rect 312544 18980 312596 19032
rect 149520 18912 149572 18964
rect 358820 18912 358872 18964
rect 150900 18844 150952 18896
rect 376760 18844 376812 18896
rect 151176 18776 151228 18828
rect 380900 18776 380952 18828
rect 156696 18708 156748 18760
rect 451280 18708 451332 18760
rect 163228 18640 163280 18692
rect 535460 18640 535512 18692
rect 35900 18572 35952 18624
rect 118148 18572 118200 18624
rect 164608 18572 164660 18624
rect 553400 18572 553452 18624
rect 142804 17620 142856 17672
rect 273260 17620 273312 17672
rect 147036 17552 147088 17604
rect 327080 17552 327132 17604
rect 154856 17484 154908 17536
rect 427820 17484 427872 17536
rect 155316 17416 155368 17468
rect 433340 17416 433392 17468
rect 155408 17348 155460 17400
rect 434720 17348 434772 17400
rect 155592 17280 155644 17332
rect 437480 17280 437532 17332
rect 164884 17212 164936 17264
rect 556252 17212 556304 17264
rect 142896 16328 142948 16380
rect 274824 16328 274876 16380
rect 143908 16260 143960 16312
rect 287336 16260 287388 16312
rect 144000 16192 144052 16244
rect 288992 16192 289044 16244
rect 144276 16124 144328 16176
rect 292672 16124 292724 16176
rect 148508 16056 148560 16108
rect 346952 16056 347004 16108
rect 149060 15988 149112 16040
rect 353576 15988 353628 16040
rect 153936 15920 153988 15972
rect 415492 15920 415544 15972
rect 162952 15852 163004 15904
rect 532056 15852 532108 15904
rect 141240 14832 141292 14884
rect 253480 14832 253532 14884
rect 141516 14764 141568 14816
rect 256700 14764 256752 14816
rect 142344 14696 142396 14748
rect 267740 14696 267792 14748
rect 142620 14628 142672 14680
rect 270776 14628 270828 14680
rect 149612 14560 149664 14612
rect 361120 14560 361172 14612
rect 151452 14492 151504 14544
rect 384304 14492 384356 14544
rect 157892 14424 157944 14476
rect 467472 14424 467524 14476
rect 139584 13404 139636 13456
rect 231860 13404 231912 13456
rect 140136 13336 140188 13388
rect 239312 13336 239364 13388
rect 146852 13268 146904 13320
rect 324412 13268 324464 13320
rect 147128 13200 147180 13252
rect 328736 13200 328788 13252
rect 149796 13132 149848 13184
rect 363512 13132 363564 13184
rect 14280 13064 14332 13116
rect 122104 13064 122156 13116
rect 150992 13064 151044 13116
rect 378416 13064 378468 13116
rect 157708 12248 157760 12300
rect 169024 12248 169076 12300
rect 138204 12180 138256 12232
rect 214472 12180 214524 12232
rect 138480 12112 138532 12164
rect 218152 12112 218204 12164
rect 138756 12044 138808 12096
rect 221096 12044 221148 12096
rect 146576 11976 146628 12028
rect 322112 11976 322164 12028
rect 148232 11908 148284 11960
rect 342904 11908 342956 11960
rect 131396 11840 131448 11892
rect 148416 11840 148468 11892
rect 345296 11840 345348 11892
rect 131120 11636 131172 11688
rect 131304 11636 131356 11688
rect 131120 11500 131172 11552
rect 149244 11772 149296 11824
rect 356336 11772 356388 11824
rect 159364 11704 159416 11756
rect 486424 11704 486476 11756
rect 176660 11636 176712 11688
rect 177856 11636 177908 11688
rect 218060 11636 218112 11688
rect 219256 11636 219308 11688
rect 242900 11636 242952 11688
rect 244096 11636 244148 11688
rect 259460 11636 259512 11688
rect 260656 11636 260708 11688
rect 110512 10956 110564 11008
rect 130384 10956 130436 11008
rect 102140 10888 102192 10940
rect 129096 10888 129148 10940
rect 95792 10820 95844 10872
rect 129004 10820 129056 10872
rect 134800 10820 134852 10872
rect 170312 10820 170364 10872
rect 92480 10752 92532 10804
rect 129188 10752 129240 10804
rect 137100 10752 137152 10804
rect 200304 10752 200356 10804
rect 75000 10684 75052 10736
rect 122196 10684 122248 10736
rect 137376 10684 137428 10736
rect 203432 10684 203484 10736
rect 78128 10616 78180 10668
rect 127808 10616 127860 10668
rect 142988 10616 143040 10668
rect 276112 10616 276164 10668
rect 67640 10548 67692 10600
rect 126428 10548 126480 10600
rect 144460 10548 144512 10600
rect 294880 10548 294932 10600
rect 64328 10480 64380 10532
rect 126336 10480 126388 10532
rect 145932 10480 145984 10532
rect 313832 10480 313884 10532
rect 46664 10412 46716 10464
rect 125048 10412 125100 10464
rect 146300 10412 146352 10464
rect 318064 10412 318116 10464
rect 31944 10344 31996 10396
rect 123668 10344 123720 10396
rect 152648 10344 152700 10396
rect 398932 10344 398984 10396
rect 25320 10276 25372 10328
rect 123576 10276 123628 10328
rect 156512 10276 156564 10328
rect 448612 10276 448664 10328
rect 117320 10208 117372 10260
rect 130568 10208 130620 10260
rect 120632 10140 120684 10192
rect 130476 10140 130528 10192
rect 116400 9596 116452 9648
rect 130200 9596 130252 9648
rect 134892 9596 134944 9648
rect 171968 9596 172020 9648
rect 112812 9528 112864 9580
rect 130292 9528 130344 9580
rect 135444 9528 135496 9580
rect 179052 9528 179104 9580
rect 60832 9460 60884 9512
rect 126152 9460 126204 9512
rect 135996 9460 136048 9512
rect 186136 9460 186188 9512
rect 57244 9392 57296 9444
rect 126244 9392 126296 9444
rect 145380 9392 145432 9444
rect 306748 9392 306800 9444
rect 43076 9324 43128 9376
rect 116584 9324 116636 9376
rect 145656 9324 145708 9376
rect 310244 9324 310296 9376
rect 50160 9256 50212 9308
rect 124864 9256 124916 9308
rect 145748 9256 145800 9308
rect 311440 9256 311492 9308
rect 45468 9188 45520 9240
rect 124772 9188 124824 9240
rect 147956 9188 148008 9240
rect 339868 9188 339920 9240
rect 41880 9120 41932 9172
rect 124956 9120 125008 9172
rect 148140 9120 148192 9172
rect 342168 9120 342220 9172
rect 31300 9052 31352 9104
rect 123484 9052 123536 9104
rect 152096 9052 152148 9104
rect 393044 9052 393096 9104
rect 24216 8984 24268 9036
rect 123392 8984 123444 9036
rect 153476 8984 153528 9036
rect 410800 8984 410852 9036
rect 9956 8916 10008 8968
rect 122012 8916 122064 8968
rect 153568 8916 153620 8968
rect 411904 8916 411956 8968
rect 98644 8236 98696 8288
rect 128912 8236 128964 8288
rect 481640 8236 481692 8288
rect 482468 8236 482520 8288
rect 95148 8168 95200 8220
rect 128728 8168 128780 8220
rect 84476 8100 84528 8152
rect 127716 8100 127768 8152
rect 80888 8032 80940 8084
rect 127440 8032 127492 8084
rect 77392 7964 77444 8016
rect 127532 7964 127584 8016
rect 73804 7896 73856 7948
rect 127624 7896 127676 7948
rect 142436 7896 142488 7948
rect 268844 7896 268896 7948
rect 66720 7828 66772 7880
rect 126060 7828 126112 7880
rect 144092 7828 144144 7880
rect 290188 7828 290240 7880
rect 63224 7760 63276 7812
rect 125968 7760 126020 7812
rect 147680 7760 147732 7812
rect 336280 7760 336332 7812
rect 27712 7692 27764 7744
rect 123208 7692 123260 7744
rect 154028 7692 154080 7744
rect 417884 7692 417936 7744
rect 19432 7624 19484 7676
rect 118056 7624 118108 7676
rect 119896 7624 119948 7676
rect 130108 7624 130160 7676
rect 164700 7624 164752 7676
rect 554964 7624 555016 7676
rect 23020 7556 23072 7608
rect 123300 7556 123352 7608
rect 164976 7556 165028 7608
rect 558552 7556 558604 7608
rect 102232 7488 102284 7540
rect 128820 7488 128872 7540
rect 115204 6808 115256 6860
rect 130016 6808 130068 6860
rect 562324 6808 562376 6860
rect 580172 6808 580224 6860
rect 99840 6740 99892 6792
rect 120816 6740 120868 6792
rect 139860 6740 139912 6792
rect 235816 6740 235868 6792
rect 59636 6672 59688 6724
rect 125876 6672 125928 6724
rect 143816 6672 143868 6724
rect 286600 6672 286652 6724
rect 11152 6604 11204 6656
rect 86224 6604 86276 6656
rect 104532 6604 104584 6656
rect 128636 6604 128688 6656
rect 151084 6604 151136 6656
rect 379980 6604 380032 6656
rect 48964 6536 49016 6588
rect 124680 6536 124732 6588
rect 152372 6536 152424 6588
rect 396540 6536 396592 6588
rect 44272 6468 44324 6520
rect 124496 6468 124548 6520
rect 167276 6468 167328 6520
rect 436744 6468 436796 6520
rect 40684 6400 40736 6452
rect 124588 6400 124640 6452
rect 161572 6400 161624 6452
rect 514760 6400 514812 6452
rect 30104 6332 30156 6384
rect 123116 6332 123168 6384
rect 163596 6332 163648 6384
rect 540796 6332 540848 6384
rect 13544 6264 13596 6316
rect 121736 6264 121788 6316
rect 163872 6264 163924 6316
rect 544384 6264 544436 6316
rect 8760 6196 8812 6248
rect 121828 6196 121880 6248
rect 165804 6196 165856 6248
rect 569132 6196 569184 6248
rect 4068 6128 4120 6180
rect 121920 6128 121972 6180
rect 166080 6128 166132 6180
rect 572720 6128 572772 6180
rect 97448 5448 97500 5500
rect 129372 5448 129424 5500
rect 93952 5380 94004 5432
rect 129280 5380 129332 5432
rect 132592 5380 132644 5432
rect 142436 5380 142488 5432
rect 85672 5312 85724 5364
rect 120724 5312 120776 5364
rect 132776 5312 132828 5364
rect 144736 5312 144788 5364
rect 86868 5244 86920 5296
rect 127348 5244 127400 5296
rect 134524 5244 134576 5296
rect 167184 5244 167236 5296
rect 76196 5176 76248 5228
rect 127164 5176 127216 5228
rect 137284 5176 137336 5228
rect 202696 5176 202748 5228
rect 72608 5108 72660 5160
rect 127256 5108 127308 5160
rect 133052 5108 133104 5160
rect 148324 5108 148376 5160
rect 149888 5108 149940 5160
rect 364616 5108 364668 5160
rect 65524 5040 65576 5092
rect 125784 5040 125836 5092
rect 133144 5040 133196 5092
rect 149520 5040 149572 5092
rect 160468 5040 160520 5092
rect 500592 5040 500644 5092
rect 33600 4972 33652 5024
rect 123024 4972 123076 5024
rect 133420 4972 133472 5024
rect 153016 4972 153068 5024
rect 160560 4972 160612 5024
rect 501788 4972 501840 5024
rect 28908 4904 28960 4956
rect 117964 4904 118016 4956
rect 118792 4904 118844 4956
rect 129924 4904 129976 4956
rect 133328 4904 133380 4956
rect 151820 4904 151872 4956
rect 161940 4904 161992 4956
rect 519544 4904 519596 4956
rect 5264 4836 5316 4888
rect 22744 4836 22796 4888
rect 26516 4836 26568 4888
rect 124128 4836 124180 4888
rect 133880 4836 133932 4888
rect 158904 4836 158956 4888
rect 162216 4836 162268 4888
rect 523040 4836 523092 4888
rect 21824 4768 21876 4820
rect 123760 4768 123812 4820
rect 134248 4768 134300 4820
rect 163688 4768 163740 4820
rect 166816 4768 166868 4820
rect 577412 4768 577464 4820
rect 111616 4700 111668 4752
rect 129832 4700 129884 4752
rect 117228 4632 117280 4684
rect 128544 4632 128596 4684
rect 101036 4088 101088 4140
rect 117228 4088 117280 4140
rect 121368 4088 121420 4140
rect 143540 4088 143592 4140
rect 168104 4088 168156 4140
rect 189724 4088 189776 4140
rect 276020 4088 276072 4140
rect 276756 4088 276808 4140
rect 284300 4088 284352 4140
rect 285036 4088 285088 4140
rect 292580 4088 292632 4140
rect 293316 4088 293368 4140
rect 312544 4088 312596 4140
rect 543188 4088 543240 4140
rect 83280 4020 83332 4072
rect 127992 4020 128044 4072
rect 131856 4020 131908 4072
rect 132960 4020 133012 4072
rect 79692 3952 79744 4004
rect 127072 3952 127124 4004
rect 132868 3952 132920 4004
rect 134064 3952 134116 4004
rect 146944 4020 146996 4072
rect 160100 4020 160152 4072
rect 167460 4020 167512 4072
rect 401324 4020 401376 4072
rect 69112 3884 69164 3936
rect 126888 3884 126940 3936
rect 132040 3884 132092 3936
rect 135260 3884 135312 3936
rect 145932 3952 145984 4004
rect 167552 3952 167604 4004
rect 408408 3952 408460 4004
rect 161296 3884 161348 3936
rect 168196 3884 168248 3936
rect 409604 3884 409656 3936
rect 58440 3816 58492 3868
rect 126520 3816 126572 3868
rect 134156 3816 134208 3868
rect 162492 3816 162544 3868
rect 168288 3816 168340 3868
rect 415400 3816 415452 3868
rect 51356 3748 51408 3800
rect 125508 3748 125560 3800
rect 134340 3748 134392 3800
rect 164884 3748 164936 3800
rect 167644 3748 167696 3800
rect 427268 3748 427320 3800
rect 47860 3680 47912 3732
rect 124312 3680 124364 3732
rect 134432 3680 134484 3732
rect 166080 3680 166132 3732
rect 167736 3680 167788 3732
rect 429660 3680 429712 3732
rect 445116 3680 445168 3732
rect 546684 3680 546736 3732
rect 39580 3612 39632 3664
rect 125232 3612 125284 3664
rect 134616 3612 134668 3664
rect 168380 3612 168432 3664
rect 169024 3612 169076 3664
rect 465172 3612 465224 3664
rect 12348 3544 12400 3596
rect 122472 3544 122524 3596
rect 125876 3544 125928 3596
rect 131120 3544 131172 3596
rect 133052 3544 133104 3596
rect 147128 3544 147180 3596
rect 159180 3544 159232 3596
rect 484032 3544 484084 3596
rect 7656 3476 7708 3528
rect 122564 3476 122616 3528
rect 129372 3476 129424 3528
rect 131212 3476 131264 3528
rect 133236 3476 133288 3528
rect 150624 3476 150676 3528
rect 159456 3476 159508 3528
rect 478052 3476 478104 3528
rect 2872 3408 2924 3460
rect 122196 3408 122248 3460
rect 126980 3408 127032 3460
rect 131396 3408 131448 3460
rect 133512 3408 133564 3460
rect 154212 3408 154264 3460
rect 159732 3408 159784 3460
rect 491116 3408 491168 3460
rect 102140 3340 102192 3392
rect 103336 3340 103388 3392
rect 122288 3340 122340 3392
rect 131028 3340 131080 3392
rect 131948 3340 132000 3392
rect 134156 3340 134208 3392
rect 137744 3340 137796 3392
rect 146944 3340 146996 3392
rect 167368 3340 167420 3392
rect 394240 3340 394292 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 415492 3340 415544 3392
rect 416688 3340 416740 3392
rect 432052 3340 432104 3392
rect 433248 3340 433300 3392
rect 440332 3340 440384 3392
rect 441528 3340 441580 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 456800 3340 456852 3392
rect 458088 3340 458140 3392
rect 473360 3340 473412 3392
rect 474188 3340 474240 3392
rect 478052 3340 478104 3392
rect 487620 3340 487672 3392
rect 130568 3272 130620 3324
rect 131488 3272 131540 3324
rect 132132 3272 132184 3324
rect 136456 3272 136508 3324
rect 149152 3272 149204 3324
rect 169576 3272 169628 3324
rect 169668 3272 169720 3324
rect 175464 3272 175516 3324
rect 193220 3272 193272 3324
rect 194416 3272 194468 3324
rect 226340 3272 226392 3324
rect 227536 3272 227588 3324
rect 299480 3272 299532 3324
rect 300768 3272 300820 3324
rect 307760 3272 307812 3324
rect 309048 3272 309100 3324
rect 316040 3272 316092 3324
rect 317328 3272 317380 3324
rect 324412 3272 324464 3324
rect 325608 3272 325660 3324
rect 332600 3272 332652 3324
rect 333888 3272 333940 3324
rect 20628 3204 20680 3256
rect 25504 3204 25556 3256
rect 165252 3204 165304 3256
rect 182548 3204 182600 3256
rect 326436 3204 326488 3256
rect 539600 3272 539652 3324
rect 349160 3204 349212 3256
rect 350448 3204 350500 3256
rect 357440 3204 357492 3256
rect 358728 3204 358780 3256
rect 365720 3204 365772 3256
rect 367008 3204 367060 3256
rect 374092 3204 374144 3256
rect 375288 3204 375340 3256
rect 382280 3204 382332 3256
rect 383568 3204 383620 3256
rect 390560 3204 390612 3256
rect 391848 3204 391900 3256
rect 128176 3136 128228 3188
rect 131580 3136 131632 3188
rect 136180 2932 136232 2984
rect 141240 2932 141292 2984
rect 423680 1232 423732 1284
rect 424968 1232 425020 1284
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3330 566944 3386 566953
rect 3330 566879 3386 566888
rect 3344 565894 3372 566879
rect 3332 565888 3384 565894
rect 3332 565830 3384 565836
rect 2778 553888 2834 553897
rect 2778 553823 2780 553832
rect 2832 553823 2834 553832
rect 2780 553794 2832 553800
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 2778 501800 2834 501809
rect 2778 501735 2834 501744
rect 2792 501090 2820 501735
rect 2780 501084 2832 501090
rect 2780 501026 2832 501032
rect 2778 462632 2834 462641
rect 2778 462567 2780 462576
rect 2832 462567 2834 462576
rect 2780 462538 2832 462544
rect 2778 449576 2834 449585
rect 2778 449511 2834 449520
rect 2792 448866 2820 449511
rect 2780 448860 2832 448866
rect 2780 448802 2832 448808
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 410106 3188 410479
rect 3148 410100 3200 410106
rect 3148 410042 3200 410048
rect 2780 397520 2832 397526
rect 2778 397488 2780 397497
rect 2832 397488 2834 397497
rect 2778 397423 2834 397432
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3344 357474 3372 358391
rect 3332 357468 3384 357474
rect 3332 357410 3384 357416
rect 2778 345400 2834 345409
rect 2778 345335 2834 345344
rect 2792 345234 2820 345335
rect 2780 345228 2832 345234
rect 2780 345170 2832 345176
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 3238 293176 3294 293185
rect 3238 293111 3294 293120
rect 3252 292602 3280 293111
rect 3240 292596 3292 292602
rect 3240 292538 3292 292544
rect 3238 267200 3294 267209
rect 3238 267135 3294 267144
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3160 253978 3188 254079
rect 3148 253972 3200 253978
rect 3148 253914 3200 253920
rect 3054 241088 3110 241097
rect 3054 241023 3110 241032
rect 3068 240174 3096 241023
rect 3056 240168 3108 240174
rect 3056 240110 3108 240116
rect 3146 214976 3202 214985
rect 3146 214911 3202 214920
rect 3160 213994 3188 214911
rect 3148 213988 3200 213994
rect 3148 213930 3200 213936
rect 2962 201920 3018 201929
rect 2962 201855 3018 201864
rect 2976 201550 3004 201855
rect 2964 201544 3016 201550
rect 2964 201486 3016 201492
rect 3146 188864 3202 188873
rect 3146 188799 3202 188808
rect 3160 187746 3188 188799
rect 3148 187740 3200 187746
rect 3148 187682 3200 187688
rect 3148 162920 3200 162926
rect 3146 162888 3148 162897
rect 3200 162888 3202 162897
rect 3146 162823 3202 162832
rect 3146 149832 3202 149841
rect 3146 149767 3202 149776
rect 3160 149122 3188 149767
rect 3148 149116 3200 149122
rect 3148 149058 3200 149064
rect 3252 136134 3280 267135
rect 3240 136128 3292 136134
rect 3240 136070 3292 136076
rect 3344 136066 3372 319223
rect 3436 138378 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3606 632088 3662 632097
rect 3606 632023 3662 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3424 138372 3476 138378
rect 3424 138314 3476 138320
rect 3422 136776 3478 136785
rect 3422 136711 3478 136720
rect 3436 136678 3464 136711
rect 3424 136672 3476 136678
rect 3424 136614 3476 136620
rect 3332 136060 3384 136066
rect 3332 136002 3384 136008
rect 3424 131164 3476 131170
rect 3424 131106 3476 131112
rect 3330 84688 3386 84697
rect 3330 84623 3386 84632
rect 3344 84250 3372 84623
rect 3332 84244 3384 84250
rect 3332 84186 3384 84192
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 3436 19417 3464 131106
rect 3528 73817 3556 606047
rect 3620 134706 3648 632023
rect 3698 580000 3754 580009
rect 3698 579935 3754 579944
rect 3712 136202 3740 579935
rect 4804 553852 4856 553858
rect 4804 553794 4856 553800
rect 3790 527912 3846 527921
rect 3790 527847 3846 527856
rect 3804 136338 3832 527847
rect 3974 475688 4030 475697
rect 3974 475623 4030 475632
rect 3882 423600 3938 423609
rect 3882 423535 3938 423544
rect 3792 136332 3844 136338
rect 3792 136274 3844 136280
rect 3896 136270 3924 423535
rect 3988 227050 4016 475623
rect 4066 371376 4122 371385
rect 4066 371311 4122 371320
rect 3976 227044 4028 227050
rect 3976 226986 4028 226992
rect 4080 142154 4108 371311
rect 3988 142126 4108 142154
rect 3988 136406 4016 142126
rect 4068 138372 4120 138378
rect 4068 138314 4120 138320
rect 3976 136400 4028 136406
rect 3976 136342 4028 136348
rect 3884 136264 3936 136270
rect 3884 136206 3936 136212
rect 3700 136196 3752 136202
rect 3700 136138 3752 136144
rect 3608 134700 3660 134706
rect 3608 134642 3660 134648
rect 4080 134638 4108 138314
rect 4068 134632 4120 134638
rect 4068 134574 4120 134580
rect 3792 133952 3844 133958
rect 3792 133894 3844 133900
rect 3608 128376 3660 128382
rect 3608 128318 3660 128324
rect 3514 73808 3570 73817
rect 3514 73743 3570 73752
rect 3516 71732 3568 71738
rect 3516 71674 3568 71680
rect 3528 71641 3556 71674
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 3620 58585 3648 128318
rect 3700 127016 3752 127022
rect 3700 126958 3752 126964
rect 3712 97617 3740 126958
rect 3804 110673 3832 133894
rect 3790 110664 3846 110673
rect 3790 110599 3846 110608
rect 3698 97608 3754 97617
rect 3698 97543 3754 97552
rect 4816 73681 4844 553794
rect 4896 501084 4948 501090
rect 4896 501026 4948 501032
rect 4908 75177 4936 501026
rect 5080 462596 5132 462602
rect 5080 462538 5132 462544
rect 4988 448860 5040 448866
rect 4988 448802 5040 448808
rect 4894 75168 4950 75177
rect 4894 75103 4950 75112
rect 5000 74089 5028 448802
rect 5092 118658 5120 462538
rect 5172 397520 5224 397526
rect 5172 397462 5224 397468
rect 5080 118652 5132 118658
rect 5080 118594 5132 118600
rect 5184 75313 5212 397462
rect 5264 345228 5316 345234
rect 5264 345170 5316 345176
rect 5170 75304 5226 75313
rect 5170 75239 5226 75248
rect 4986 74080 5042 74089
rect 4986 74015 5042 74024
rect 5276 73710 5304 345170
rect 5264 73704 5316 73710
rect 4802 73672 4858 73681
rect 5264 73646 5316 73652
rect 4802 73607 4858 73616
rect 6932 71670 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 15844 670744 15896 670750
rect 15844 670686 15896 670692
rect 8944 410100 8996 410106
rect 8944 410042 8996 410048
rect 8956 120086 8984 410042
rect 10324 357468 10376 357474
rect 10324 357410 10376 357416
rect 10336 121446 10364 357410
rect 10324 121440 10376 121446
rect 10324 121382 10376 121388
rect 8944 120080 8996 120086
rect 8944 120022 8996 120028
rect 15856 111790 15884 670686
rect 22744 253972 22796 253978
rect 22744 253914 22796 253920
rect 22756 124166 22784 253914
rect 22836 201544 22888 201550
rect 22836 201486 22888 201492
rect 22848 125594 22876 201486
rect 22836 125588 22888 125594
rect 22836 125530 22888 125536
rect 22744 124160 22796 124166
rect 22744 124102 22796 124108
rect 15844 111784 15896 111790
rect 15844 111726 15896 111732
rect 23492 110430 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 37924 618316 37976 618322
rect 37924 618258 37976 618264
rect 29644 565888 29696 565894
rect 29644 565830 29696 565836
rect 24124 305040 24176 305046
rect 24124 304982 24176 304988
rect 24136 122806 24164 304982
rect 25504 149116 25556 149122
rect 25504 149058 25556 149064
rect 25516 126954 25544 149058
rect 25504 126948 25556 126954
rect 25504 126890 25556 126896
rect 24124 122800 24176 122806
rect 24124 122742 24176 122748
rect 29656 115938 29684 565830
rect 33784 514820 33836 514826
rect 33784 514762 33836 514768
rect 29736 292596 29788 292602
rect 29736 292538 29788 292544
rect 29644 115932 29696 115938
rect 29644 115874 29696 115880
rect 23480 110424 23532 110430
rect 23480 110366 23532 110372
rect 29748 75274 29776 292538
rect 33796 117298 33824 514762
rect 33784 117292 33836 117298
rect 33784 117234 33836 117240
rect 37936 113150 37964 618258
rect 40052 136474 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 59268 609272 59320 609278
rect 59268 609214 59320 609220
rect 59280 606490 59308 609214
rect 53104 606484 53156 606490
rect 53104 606426 53156 606432
rect 59268 606484 59320 606490
rect 59268 606426 59320 606432
rect 53116 559774 53144 606426
rect 46204 559768 46256 559774
rect 46204 559710 46256 559716
rect 53104 559768 53156 559774
rect 53104 559710 53156 559716
rect 46216 517546 46244 559710
rect 62672 537532 62724 537538
rect 62672 537474 62724 537480
rect 62684 533050 62712 537474
rect 61384 533044 61436 533050
rect 61384 532986 61436 532992
rect 62672 533044 62724 533050
rect 62672 532986 62724 532992
rect 45100 517540 45152 517546
rect 45100 517482 45152 517488
rect 46204 517540 46256 517546
rect 46204 517482 46256 517488
rect 45008 240780 45060 240786
rect 45008 240722 45060 240728
rect 44824 240168 44876 240174
rect 44824 240110 44876 240116
rect 44732 239760 44784 239766
rect 44732 239702 44784 239708
rect 44744 227730 44772 239702
rect 44732 227724 44784 227730
rect 44732 227666 44784 227672
rect 40040 136468 40092 136474
rect 40040 136410 40092 136416
rect 37924 113144 37976 113150
rect 37924 113086 37976 113092
rect 29736 75268 29788 75274
rect 29736 75210 29788 75216
rect 44836 73642 44864 240110
rect 44916 238808 44968 238814
rect 44916 238750 44968 238756
rect 44928 232966 44956 238750
rect 44916 232960 44968 232966
rect 44916 232902 44968 232908
rect 45020 232830 45048 240722
rect 45008 232824 45060 232830
rect 45008 232766 45060 232772
rect 45112 221134 45140 517482
rect 61396 376650 61424 532986
rect 58624 376644 58676 376650
rect 58624 376586 58676 376592
rect 61384 376644 61436 376650
rect 61384 376586 61436 376592
rect 58636 346390 58664 376586
rect 69664 356720 69716 356726
rect 69664 356662 69716 356668
rect 56876 346384 56928 346390
rect 56876 346326 56928 346332
rect 58624 346384 58676 346390
rect 58624 346326 58676 346332
rect 56888 338298 56916 346326
rect 69676 339726 69704 356662
rect 68284 339720 68336 339726
rect 68284 339662 68336 339668
rect 69664 339720 69716 339726
rect 69664 339662 69716 339668
rect 55864 338292 55916 338298
rect 55864 338234 55916 338240
rect 56876 338292 56928 338298
rect 56876 338234 56928 338240
rect 48964 331900 49016 331906
rect 48964 331842 49016 331848
rect 48976 302258 49004 331842
rect 55876 323406 55904 338234
rect 66260 336048 66312 336054
rect 66260 335990 66312 335996
rect 66272 331906 66300 335990
rect 66260 331900 66312 331906
rect 66260 331842 66312 331848
rect 53104 323400 53156 323406
rect 53104 323342 53156 323348
rect 55864 323400 55916 323406
rect 55864 323342 55916 323348
rect 53116 305046 53144 323342
rect 62764 313948 62816 313954
rect 62764 313890 62816 313896
rect 51724 305040 51776 305046
rect 51724 304982 51776 304988
rect 53104 305040 53156 305046
rect 53104 304982 53156 304988
rect 46204 302252 46256 302258
rect 46204 302194 46256 302200
rect 48964 302252 49016 302258
rect 48964 302194 49016 302200
rect 46216 273222 46244 302194
rect 45376 273216 45428 273222
rect 45376 273158 45428 273164
rect 46204 273216 46256 273222
rect 46204 273158 46256 273164
rect 45388 248414 45416 273158
rect 51080 266416 51132 266422
rect 51080 266358 51132 266364
rect 50344 262880 50396 262886
rect 50344 262822 50396 262828
rect 47584 260500 47636 260506
rect 47584 260442 47636 260448
rect 47492 256760 47544 256766
rect 47492 256702 47544 256708
rect 47504 253978 47532 256702
rect 45836 253972 45888 253978
rect 45836 253914 45888 253920
rect 47492 253972 47544 253978
rect 47492 253914 47544 253920
rect 45848 248414 45876 253914
rect 46940 249484 46992 249490
rect 46940 249426 46992 249432
rect 45296 248386 45416 248414
rect 45756 248386 45876 248414
rect 45192 242276 45244 242282
rect 45192 242218 45244 242224
rect 45204 231130 45232 242218
rect 45296 231946 45324 248386
rect 45560 241392 45612 241398
rect 45560 241334 45612 241340
rect 45376 240848 45428 240854
rect 45376 240790 45428 240796
rect 45284 231940 45336 231946
rect 45284 231882 45336 231888
rect 45388 231878 45416 240790
rect 45468 239420 45520 239426
rect 45468 239362 45520 239368
rect 45480 231878 45508 239362
rect 45376 231872 45428 231878
rect 45376 231814 45428 231820
rect 45468 231872 45520 231878
rect 45468 231814 45520 231820
rect 45192 231124 45244 231130
rect 45192 231066 45244 231072
rect 45100 221128 45152 221134
rect 45100 221070 45152 221076
rect 45572 172514 45600 241334
rect 45652 241324 45704 241330
rect 45652 241266 45704 241272
rect 45664 217326 45692 241266
rect 45756 238814 45784 248386
rect 46952 242282 46980 249426
rect 46940 242276 46992 242282
rect 46940 242218 46992 242224
rect 45836 241460 45888 241466
rect 45836 241402 45888 241408
rect 45744 238808 45796 238814
rect 45744 238750 45796 238756
rect 45848 232898 45876 241402
rect 47596 241330 47624 260442
rect 49240 259004 49292 259010
rect 49240 258946 49292 258952
rect 49252 256766 49280 258946
rect 49240 256760 49292 256766
rect 49240 256702 49292 256708
rect 50356 252618 50384 262822
rect 50896 261248 50948 261254
rect 50896 261190 50948 261196
rect 50908 259010 50936 261190
rect 51092 260506 51120 266358
rect 51080 260500 51132 260506
rect 51080 260442 51132 260448
rect 50896 259004 50948 259010
rect 50896 258946 50948 258952
rect 48688 252612 48740 252618
rect 48688 252554 48740 252560
rect 50344 252612 50396 252618
rect 50344 252554 50396 252560
rect 47676 251864 47728 251870
rect 47676 251806 47728 251812
rect 47688 241398 47716 251806
rect 48700 249490 48728 252554
rect 48688 249484 48740 249490
rect 48688 249426 48740 249432
rect 51736 245682 51764 304982
rect 57244 301504 57296 301510
rect 57244 301446 57296 301452
rect 57256 288386 57284 301446
rect 62776 301102 62804 313890
rect 61384 301096 61436 301102
rect 61384 301038 61436 301044
rect 62764 301096 62816 301102
rect 62764 301038 62816 301044
rect 55864 288380 55916 288386
rect 55864 288322 55916 288328
rect 57244 288380 57296 288386
rect 57244 288322 57296 288328
rect 55876 272950 55904 288322
rect 61396 280838 61424 301038
rect 68296 300218 68324 339662
rect 66904 300212 66956 300218
rect 66904 300154 66956 300160
rect 68284 300212 68336 300218
rect 68284 300154 68336 300160
rect 60004 280832 60056 280838
rect 60004 280774 60056 280780
rect 61384 280832 61436 280838
rect 61384 280774 61436 280780
rect 60016 274718 60044 280774
rect 57980 274712 58032 274718
rect 57980 274654 58032 274660
rect 60004 274712 60056 274718
rect 60004 274654 60056 274660
rect 54484 272944 54536 272950
rect 54484 272886 54536 272892
rect 55864 272944 55916 272950
rect 55864 272886 55916 272892
rect 52368 269136 52420 269142
rect 52368 269078 52420 269084
rect 52380 261254 52408 269078
rect 54496 266422 54524 272886
rect 57992 270586 58020 274654
rect 57900 270558 58020 270586
rect 57900 269142 57928 270558
rect 57888 269136 57940 269142
rect 57888 269078 57940 269084
rect 66916 266422 66944 300154
rect 54484 266416 54536 266422
rect 54484 266358 54536 266364
rect 63500 266416 63552 266422
rect 63500 266358 63552 266364
rect 66904 266416 66956 266422
rect 66904 266358 66956 266364
rect 63512 262886 63540 266358
rect 63500 262880 63552 262886
rect 63500 262822 63552 262828
rect 52368 261248 52420 261254
rect 52368 261190 52420 261196
rect 71792 251870 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 78588 362228 78640 362234
rect 78588 362170 78640 362176
rect 78600 357814 78628 362170
rect 75184 357808 75236 357814
rect 75184 357750 75236 357756
rect 78588 357808 78640 357814
rect 78588 357750 78640 357756
rect 75196 336054 75224 357750
rect 75184 336048 75236 336054
rect 75184 335990 75236 335996
rect 88352 318170 88380 702406
rect 103520 365696 103572 365702
rect 103520 365638 103572 365644
rect 103532 362234 103560 365638
rect 103520 362228 103572 362234
rect 103520 362170 103572 362176
rect 103520 355836 103572 355842
rect 103520 355778 103572 355784
rect 103532 351898 103560 355778
rect 98644 351892 98696 351898
rect 98644 351834 98696 351840
rect 103520 351892 103572 351898
rect 103520 351834 103572 351840
rect 98656 340950 98684 351834
rect 94504 340944 94556 340950
rect 94504 340886 94556 340892
rect 98644 340944 98696 340950
rect 98644 340886 98696 340892
rect 85580 318164 85632 318170
rect 85580 318106 85632 318112
rect 88340 318164 88392 318170
rect 88340 318106 88392 318112
rect 85592 313410 85620 318106
rect 79324 313404 79376 313410
rect 79324 313346 79376 313352
rect 85580 313404 85632 313410
rect 85580 313346 85632 313352
rect 79336 301510 79364 313346
rect 94516 311574 94544 340886
rect 104912 313954 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 134524 672104 134576 672110
rect 134524 672046 134576 672052
rect 134536 651914 134564 672046
rect 131764 651908 131816 651914
rect 131764 651850 131816 651856
rect 134524 651908 134576 651914
rect 134524 651850 134576 651856
rect 131776 621042 131804 651850
rect 136548 638920 136600 638926
rect 136548 638862 136600 638868
rect 136560 635594 136588 638862
rect 134524 635588 134576 635594
rect 134524 635530 134576 635536
rect 136548 635588 136600 635594
rect 136548 635530 136600 635536
rect 123484 621036 123536 621042
rect 123484 620978 123536 620984
rect 131764 621036 131816 621042
rect 131764 620978 131816 620984
rect 123496 609278 123524 620978
rect 123484 609272 123536 609278
rect 123484 609214 123536 609220
rect 134536 597582 134564 635530
rect 131764 597576 131816 597582
rect 131764 597518 131816 597524
rect 134524 597576 134576 597582
rect 134524 597518 134576 597524
rect 131776 533390 131804 597518
rect 130384 533384 130436 533390
rect 130384 533326 130436 533332
rect 131764 533384 131816 533390
rect 131764 533326 131816 533332
rect 130396 527202 130424 533326
rect 129004 527196 129056 527202
rect 129004 527138 129056 527144
rect 130384 527196 130436 527202
rect 130384 527138 130436 527144
rect 117964 508564 118016 508570
rect 117964 508506 118016 508512
rect 117976 487218 118004 508506
rect 129016 500954 129044 527138
rect 136652 508570 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 699718 154160 703520
rect 170324 702434 170352 703520
rect 169772 702406 170352 702434
rect 155224 700324 155276 700330
rect 155224 700266 155276 700272
rect 153016 699712 153068 699718
rect 153016 699654 153068 699660
rect 154120 699712 154172 699718
rect 154120 699654 154172 699660
rect 153028 697746 153056 699654
rect 149704 697740 149756 697746
rect 149704 697682 149756 697688
rect 153016 697740 153068 697746
rect 153016 697682 153068 697688
rect 140780 675504 140832 675510
rect 140780 675446 140832 675452
rect 140792 672110 140820 675446
rect 149716 673538 149744 697682
rect 155236 675510 155264 700266
rect 155224 675504 155276 675510
rect 155224 675446 155276 675452
rect 149704 673532 149756 673538
rect 149704 673474 149756 673480
rect 145564 673464 145616 673470
rect 145564 673406 145616 673412
rect 140780 672104 140832 672110
rect 140780 672046 140832 672052
rect 145576 658170 145604 673406
rect 143172 658164 143224 658170
rect 143172 658106 143224 658112
rect 145564 658164 145616 658170
rect 145564 658106 145616 658112
rect 143184 655586 143212 658106
rect 141424 655580 141476 655586
rect 141424 655522 141476 655528
rect 143172 655580 143224 655586
rect 143172 655522 143224 655528
rect 141436 641782 141464 655522
rect 139400 641776 139452 641782
rect 139400 641718 139452 641724
rect 141424 641776 141476 641782
rect 141424 641718 141476 641724
rect 139412 638994 139440 641718
rect 139400 638988 139452 638994
rect 139400 638930 139452 638936
rect 169772 537538 169800 702406
rect 202800 700330 202828 703520
rect 202788 700324 202840 700330
rect 202788 700266 202840 700272
rect 218072 683114 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 217980 683086 218100 683114
rect 217980 673538 218008 683086
rect 217968 673532 218020 673538
rect 217968 673474 218020 673480
rect 212540 673464 212592 673470
rect 212540 673406 212592 673412
rect 212552 667962 212580 673406
rect 212540 667956 212592 667962
rect 212540 667898 212592 667904
rect 211068 667888 211120 667894
rect 211068 667830 211120 667836
rect 211080 663814 211108 667830
rect 234632 665854 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 695162 267688 703520
rect 283852 696386 283880 703520
rect 282184 696380 282236 696386
rect 282184 696322 282236 696328
rect 283840 696380 283892 696386
rect 283840 696322 283892 696328
rect 264244 695156 264296 695162
rect 264244 695098 264296 695104
rect 267648 695156 267700 695162
rect 267648 695098 267700 695104
rect 226984 665848 227036 665854
rect 226984 665790 227036 665796
rect 234620 665848 234672 665854
rect 234620 665790 234672 665796
rect 209044 663808 209096 663814
rect 209044 663750 209096 663756
rect 211068 663808 211120 663814
rect 211068 663750 211120 663756
rect 209056 644502 209084 663750
rect 209044 644496 209096 644502
rect 209044 644438 209096 644444
rect 204904 644428 204956 644434
rect 204904 644370 204956 644376
rect 204916 630698 204944 644370
rect 226996 640354 227024 665790
rect 264256 658238 264284 695098
rect 282196 687274 282224 696322
rect 299492 694822 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 700330 332548 703520
rect 332508 700324 332560 700330
rect 332508 700266 332560 700272
rect 340144 700324 340196 700330
rect 340144 700266 340196 700272
rect 299480 694816 299532 694822
rect 299480 694758 299532 694764
rect 309784 694816 309836 694822
rect 309784 694758 309836 694764
rect 282184 687268 282236 687274
rect 282184 687210 282236 687216
rect 278688 687200 278740 687206
rect 278688 687142 278740 687148
rect 278700 684554 278728 687142
rect 309796 685166 309824 694758
rect 309784 685160 309836 685166
rect 309784 685102 309836 685108
rect 327724 685160 327776 685166
rect 327724 685102 327776 685108
rect 276664 684548 276716 684554
rect 276664 684490 276716 684496
rect 278688 684548 278740 684554
rect 278688 684490 278740 684496
rect 258724 658232 258776 658238
rect 258724 658174 258776 658180
rect 264244 658232 264296 658238
rect 264244 658174 264296 658180
rect 224224 640348 224276 640354
rect 224224 640290 224276 640296
rect 226984 640348 227036 640354
rect 226984 640290 227036 640296
rect 224236 634098 224264 640290
rect 258736 634098 258764 658174
rect 211804 634092 211856 634098
rect 211804 634034 211856 634040
rect 224224 634092 224276 634098
rect 224224 634034 224276 634040
rect 247040 634092 247092 634098
rect 247040 634034 247092 634040
rect 258724 634092 258776 634098
rect 258724 634034 258776 634040
rect 203524 630692 203576 630698
rect 203524 630634 203576 630640
rect 204904 630692 204956 630698
rect 204904 630634 204956 630640
rect 203536 610570 203564 630634
rect 211816 623830 211844 634034
rect 247052 629678 247080 634034
rect 276676 630698 276704 684490
rect 327736 655518 327764 685102
rect 327724 655512 327776 655518
rect 327724 655454 327776 655460
rect 332692 655512 332744 655518
rect 332692 655454 332744 655460
rect 332704 650010 332732 655454
rect 332692 650004 332744 650010
rect 332692 649946 332744 649952
rect 337384 650004 337436 650010
rect 337384 649946 337436 649952
rect 337396 642190 337424 649946
rect 337384 642184 337436 642190
rect 337384 642126 337436 642132
rect 340156 641034 340184 700266
rect 348804 696250 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 696244 348844 696250
rect 348792 696186 348844 696192
rect 359464 696244 359516 696250
rect 359464 696186 359516 696192
rect 359476 686526 359504 696186
rect 359464 686520 359516 686526
rect 359464 686462 359516 686468
rect 364352 683806 364380 702406
rect 371884 686520 371936 686526
rect 371884 686462 371936 686468
rect 364340 683800 364392 683806
rect 364340 683742 364392 683748
rect 371896 679658 371924 686462
rect 375380 683800 375432 683806
rect 375380 683742 375432 683748
rect 371884 679652 371936 679658
rect 371884 679594 371936 679600
rect 375392 678298 375420 683742
rect 381544 679652 381596 679658
rect 381544 679594 381596 679600
rect 375380 678292 375432 678298
rect 375380 678234 375432 678240
rect 381556 646542 381584 679594
rect 388444 678292 388496 678298
rect 388444 678234 388496 678240
rect 388456 671158 388484 678234
rect 388444 671152 388496 671158
rect 388444 671094 388496 671100
rect 391940 671152 391992 671158
rect 391940 671094 391992 671100
rect 391952 665242 391980 671094
rect 391940 665236 391992 665242
rect 391940 665178 391992 665184
rect 395344 665236 395396 665242
rect 395344 665178 395396 665184
rect 381544 646536 381596 646542
rect 381544 646478 381596 646484
rect 343640 642184 343692 642190
rect 343640 642126 343692 642132
rect 340144 641028 340196 641034
rect 340144 640970 340196 640976
rect 343652 639606 343680 642126
rect 352564 641028 352616 641034
rect 352564 640970 352616 640976
rect 343640 639600 343692 639606
rect 343640 639542 343692 639548
rect 349160 639600 349212 639606
rect 349160 639542 349212 639548
rect 349172 637566 349200 639542
rect 349160 637560 349212 637566
rect 349160 637502 349212 637508
rect 275376 630692 275428 630698
rect 275376 630634 275428 630640
rect 276664 630692 276716 630698
rect 276664 630634 276716 630640
rect 243544 629672 243596 629678
rect 243544 629614 243596 629620
rect 247040 629672 247092 629678
rect 247040 629614 247092 629620
rect 209044 623824 209096 623830
rect 209044 623766 209096 623772
rect 211804 623824 211856 623830
rect 211804 623766 211856 623772
rect 200764 610564 200816 610570
rect 200764 610506 200816 610512
rect 203524 610564 203576 610570
rect 203524 610506 203576 610512
rect 200776 593366 200804 610506
rect 195244 593360 195296 593366
rect 195244 593302 195296 593308
rect 200764 593360 200816 593366
rect 200764 593302 200816 593308
rect 195256 560318 195284 593302
rect 209056 583778 209084 623766
rect 243556 613426 243584 629614
rect 275388 628794 275416 630634
rect 273904 628788 273956 628794
rect 273904 628730 273956 628736
rect 275376 628788 275428 628794
rect 275376 628730 275428 628736
rect 273916 622470 273944 628730
rect 352576 623082 352604 640970
rect 352656 637560 352708 637566
rect 352656 637502 352708 637508
rect 352668 624442 352696 637502
rect 352656 624436 352708 624442
rect 352656 624378 352708 624384
rect 370504 624436 370556 624442
rect 370504 624378 370556 624384
rect 352564 623076 352616 623082
rect 352564 623018 352616 623024
rect 360200 623076 360252 623082
rect 360200 623018 360252 623024
rect 271144 622464 271196 622470
rect 271144 622406 271196 622412
rect 273904 622464 273956 622470
rect 273904 622406 273956 622412
rect 233148 613420 233200 613426
rect 233148 613362 233200 613368
rect 243544 613420 243596 613426
rect 243544 613362 243596 613368
rect 233160 609278 233188 613362
rect 271156 612814 271184 622406
rect 360212 619614 360240 623018
rect 360200 619608 360252 619614
rect 360200 619550 360252 619556
rect 362960 619608 363012 619614
rect 362960 619550 363012 619556
rect 362972 616146 363000 619550
rect 362960 616140 363012 616146
rect 362960 616082 363012 616088
rect 268384 612808 268436 612814
rect 268384 612750 268436 612756
rect 271144 612808 271196 612814
rect 271144 612750 271196 612756
rect 224224 609272 224276 609278
rect 224224 609214 224276 609220
rect 233148 609272 233200 609278
rect 233148 609214 233200 609220
rect 224236 591326 224264 609214
rect 268396 604518 268424 612750
rect 267004 604512 267056 604518
rect 267004 604454 267056 604460
rect 268384 604512 268436 604518
rect 268384 604454 268436 604460
rect 214564 591320 214616 591326
rect 214564 591262 214616 591268
rect 224224 591320 224276 591326
rect 224224 591262 224276 591268
rect 214576 585206 214604 591262
rect 211804 585200 211856 585206
rect 211804 585142 211856 585148
rect 214564 585200 214616 585206
rect 214564 585142 214616 585148
rect 200764 583772 200816 583778
rect 200764 583714 200816 583720
rect 209044 583772 209096 583778
rect 209044 583714 209096 583720
rect 200776 565010 200804 583714
rect 198004 565004 198056 565010
rect 198004 564946 198056 564952
rect 200764 565004 200816 565010
rect 200764 564946 200816 564952
rect 193956 560312 194008 560318
rect 193956 560254 194008 560260
rect 195244 560312 195296 560318
rect 195244 560254 195296 560260
rect 193968 558618 193996 560254
rect 192484 558612 192536 558618
rect 192484 558554 192536 558560
rect 193956 558612 194008 558618
rect 193956 558554 194008 558560
rect 192496 546514 192524 558554
rect 191104 546508 191156 546514
rect 191104 546450 191156 546456
rect 192484 546508 192536 546514
rect 192484 546450 192536 546456
rect 189724 538892 189776 538898
rect 189724 538834 189776 538840
rect 169760 537532 169812 537538
rect 169760 537474 169812 537480
rect 188344 535152 188396 535158
rect 188344 535094 188396 535100
rect 153200 511284 153252 511290
rect 153200 511226 153252 511232
rect 136640 508564 136692 508570
rect 136640 508506 136692 508512
rect 153212 507890 153240 511226
rect 150440 507884 150492 507890
rect 150440 507826 150492 507832
rect 153200 507884 153252 507890
rect 153200 507826 153252 507832
rect 150452 501770 150480 507826
rect 143540 501764 143592 501770
rect 143540 501706 143592 501712
rect 150440 501764 150492 501770
rect 150440 501706 150492 501712
rect 126980 500948 127032 500954
rect 126980 500890 127032 500896
rect 129004 500948 129056 500954
rect 129004 500890 129056 500896
rect 126992 496874 127020 500890
rect 126980 496868 127032 496874
rect 126980 496810 127032 496816
rect 124864 496800 124916 496806
rect 124864 496742 124916 496748
rect 116584 487212 116636 487218
rect 116584 487154 116636 487160
rect 117964 487212 118016 487218
rect 117964 487154 118016 487160
rect 116596 473006 116624 487154
rect 124876 474026 124904 496742
rect 143552 496738 143580 501706
rect 180064 498840 180116 498846
rect 180064 498782 180116 498788
rect 140044 496732 140096 496738
rect 140044 496674 140096 496680
rect 143540 496732 143592 496738
rect 143540 496674 143592 496680
rect 140056 487218 140084 496674
rect 136456 487212 136508 487218
rect 136456 487154 136508 487160
rect 140044 487212 140096 487218
rect 140044 487154 140096 487160
rect 136468 481506 136496 487154
rect 180076 482050 180104 498782
rect 175924 482044 175976 482050
rect 175924 481986 175976 481992
rect 180064 482044 180116 482050
rect 180064 481986 180116 481992
rect 133144 481500 133196 481506
rect 133144 481442 133196 481448
rect 136456 481500 136508 481506
rect 136456 481442 136508 481448
rect 123484 474020 123536 474026
rect 123484 473962 123536 473968
rect 124864 474020 124916 474026
rect 124864 473962 124916 473968
rect 115204 473000 115256 473006
rect 115204 472942 115256 472948
rect 116584 473000 116636 473006
rect 116584 472942 116636 472948
rect 113916 405476 113968 405482
rect 113916 405418 113968 405424
rect 113928 398546 113956 405418
rect 112444 398540 112496 398546
rect 112444 398482 112496 398488
rect 113916 398540 113968 398546
rect 113916 398482 113968 398488
rect 112456 392018 112484 398482
rect 110420 392012 110472 392018
rect 110420 391954 110472 391960
rect 112444 392012 112496 392018
rect 112444 391954 112496 391960
rect 110432 384674 110460 391954
rect 112444 385688 112496 385694
rect 112444 385630 112496 385636
rect 106924 384668 106976 384674
rect 106924 384610 106976 384616
rect 110420 384668 110472 384674
rect 110420 384610 110472 384616
rect 106936 357610 106964 384610
rect 112456 365702 112484 385630
rect 112444 365696 112496 365702
rect 112444 365638 112496 365644
rect 105268 357604 105320 357610
rect 105268 357546 105320 357552
rect 106924 357604 106976 357610
rect 106924 357546 106976 357552
rect 105280 355842 105308 357546
rect 115216 356726 115244 472942
rect 123496 465050 123524 473962
rect 122104 465044 122156 465050
rect 122104 464986 122156 464992
rect 123484 465044 123536 465050
rect 123484 464986 123536 464992
rect 122116 446214 122144 464986
rect 133156 449954 133184 481442
rect 175936 460222 175964 481986
rect 163504 460216 163556 460222
rect 163504 460158 163556 460164
rect 175924 460216 175976 460222
rect 175924 460158 175976 460164
rect 127624 449948 127676 449954
rect 127624 449890 127676 449896
rect 133144 449948 133196 449954
rect 133144 449890 133196 449896
rect 119436 446208 119488 446214
rect 119436 446150 119488 446156
rect 122104 446208 122156 446214
rect 122104 446150 122156 446156
rect 119448 433294 119476 446150
rect 117964 433288 118016 433294
rect 117964 433230 118016 433236
rect 119436 433288 119488 433294
rect 119436 433230 119488 433236
rect 117976 416770 118004 433230
rect 127636 432614 127664 449890
rect 163516 447030 163544 460158
rect 188356 455462 188384 535094
rect 189736 511290 189764 538834
rect 191116 535158 191144 546450
rect 198016 538898 198044 564946
rect 211816 549302 211844 585142
rect 267016 572762 267044 604454
rect 370516 602410 370544 624378
rect 373264 616140 373316 616146
rect 373264 616082 373316 616088
rect 370504 602404 370556 602410
rect 370504 602346 370556 602352
rect 373276 599622 373304 616082
rect 387064 602404 387116 602410
rect 387064 602346 387116 602352
rect 373264 599616 373316 599622
rect 373264 599558 373316 599564
rect 387076 574054 387104 602346
rect 387064 574048 387116 574054
rect 387064 573990 387116 573996
rect 393964 574048 394016 574054
rect 393964 573990 394016 573996
rect 265716 572756 265768 572762
rect 265716 572698 265768 572704
rect 267004 572756 267056 572762
rect 267004 572698 267056 572704
rect 265728 570722 265756 572698
rect 264244 570716 264296 570722
rect 264244 570658 264296 570664
rect 265716 570716 265768 570722
rect 265716 570658 265768 570664
rect 264256 553450 264284 570658
rect 393976 562698 394004 573990
rect 393964 562692 394016 562698
rect 393964 562634 394016 562640
rect 261484 553444 261536 553450
rect 261484 553386 261536 553392
rect 264244 553444 264296 553450
rect 264244 553386 264296 553392
rect 206284 549296 206336 549302
rect 206284 549238 206336 549244
rect 211804 549296 211856 549302
rect 211804 549238 211856 549244
rect 198004 538892 198056 538898
rect 198004 538834 198056 538840
rect 191104 535152 191156 535158
rect 191104 535094 191156 535100
rect 206296 524482 206324 549238
rect 261496 531282 261524 553386
rect 260104 531276 260156 531282
rect 260104 531218 260156 531224
rect 261484 531276 261536 531282
rect 261484 531218 261536 531224
rect 200764 524476 200816 524482
rect 200764 524418 200816 524424
rect 206284 524476 206336 524482
rect 206284 524418 206336 524424
rect 189724 511284 189776 511290
rect 189724 511226 189776 511232
rect 200776 505782 200804 524418
rect 260116 518974 260144 531218
rect 257344 518968 257396 518974
rect 257344 518910 257396 518916
rect 260104 518968 260156 518974
rect 260104 518910 260156 518916
rect 192484 505776 192536 505782
rect 192484 505718 192536 505724
rect 200764 505776 200816 505782
rect 200764 505718 200816 505724
rect 192496 498846 192524 505718
rect 257356 502382 257384 518910
rect 257344 502376 257396 502382
rect 257344 502318 257396 502324
rect 253940 502308 253992 502314
rect 253940 502250 253992 502256
rect 192484 498840 192536 498846
rect 192484 498782 192536 498788
rect 253952 498234 253980 502250
rect 253940 498228 253992 498234
rect 253940 498170 253992 498176
rect 249524 498160 249576 498166
rect 249524 498102 249576 498108
rect 249536 495514 249564 498102
rect 246304 495508 246356 495514
rect 246304 495450 246356 495456
rect 249524 495508 249576 495514
rect 249524 495450 249576 495456
rect 246316 472054 246344 495450
rect 246304 472048 246356 472054
rect 246304 471990 246356 471996
rect 239404 471980 239456 471986
rect 239404 471922 239456 471928
rect 188344 455456 188396 455462
rect 188344 455398 188396 455404
rect 182824 455388 182876 455394
rect 182824 455330 182876 455336
rect 160744 447024 160796 447030
rect 160744 446966 160796 446972
rect 163504 447024 163556 447030
rect 163504 446966 163556 446972
rect 119344 432608 119396 432614
rect 119344 432550 119396 432556
rect 127624 432608 127676 432614
rect 127624 432550 127676 432556
rect 116584 416764 116636 416770
rect 116584 416706 116636 416712
rect 117964 416764 118016 416770
rect 117964 416706 118016 416712
rect 116596 407250 116624 416706
rect 115296 407244 115348 407250
rect 115296 407186 115348 407192
rect 116584 407244 116636 407250
rect 116584 407186 116636 407192
rect 115308 405482 115336 407186
rect 115296 405476 115348 405482
rect 115296 405418 115348 405424
rect 119356 385694 119384 432550
rect 119344 385688 119396 385694
rect 119344 385630 119396 385636
rect 160756 379574 160784 446966
rect 182836 438938 182864 455330
rect 239416 451314 239444 471922
rect 238024 451308 238076 451314
rect 238024 451250 238076 451256
rect 239404 451308 239456 451314
rect 239404 451250 239456 451256
rect 181444 438932 181496 438938
rect 181444 438874 181496 438880
rect 182824 438932 182876 438938
rect 182824 438874 182876 438880
rect 181456 414050 181484 438874
rect 238036 427854 238064 451250
rect 236644 427848 236696 427854
rect 236644 427790 236696 427796
rect 238024 427848 238076 427854
rect 238024 427790 238076 427796
rect 179328 414044 179380 414050
rect 179328 413986 179380 413992
rect 181444 414044 181496 414050
rect 181444 413986 181496 413992
rect 179340 409902 179368 413986
rect 177304 409896 177356 409902
rect 177304 409838 177356 409844
rect 179328 409896 179380 409902
rect 179328 409838 179380 409844
rect 157984 379568 158036 379574
rect 157984 379510 158036 379516
rect 160744 379568 160796 379574
rect 160744 379510 160796 379516
rect 115204 356720 115256 356726
rect 115204 356662 115256 356668
rect 105268 355836 105320 355842
rect 105268 355778 105320 355784
rect 104900 313948 104952 313954
rect 104900 313890 104952 313896
rect 93124 311568 93176 311574
rect 93124 311510 93176 311516
rect 94504 311568 94556 311574
rect 94504 311510 94556 311516
rect 79324 301504 79376 301510
rect 79324 301446 79376 301452
rect 93136 289814 93164 311510
rect 157340 305040 157392 305046
rect 157340 304982 157392 304988
rect 157352 302326 157380 304982
rect 155960 302320 156012 302326
rect 155960 302262 156012 302268
rect 157340 302320 157392 302326
rect 157340 302262 157392 302268
rect 155224 302252 155276 302258
rect 155224 302194 155276 302200
rect 152004 298580 152056 298586
rect 152004 298522 152056 298528
rect 150440 295996 150492 296002
rect 150440 295938 150492 295944
rect 150452 292602 150480 295938
rect 152016 294098 152044 298522
rect 155236 296002 155264 302194
rect 155972 300914 156000 302262
rect 157996 302258 158024 379510
rect 177316 375358 177344 409838
rect 236656 404326 236684 427790
rect 233884 404320 233936 404326
rect 233884 404262 233936 404268
rect 236644 404320 236696 404326
rect 236644 404262 236696 404268
rect 175280 375352 175332 375358
rect 175280 375294 175332 375300
rect 177304 375352 177356 375358
rect 177304 375294 177356 375300
rect 175292 371278 175320 375294
rect 175280 371272 175332 371278
rect 175280 371214 175332 371220
rect 173164 371204 173216 371210
rect 173164 371146 173216 371152
rect 173176 349178 173204 371146
rect 233896 349518 233924 404262
rect 231124 349512 231176 349518
rect 231124 349454 231176 349460
rect 233884 349512 233936 349518
rect 233884 349454 233936 349460
rect 172152 349172 172204 349178
rect 172152 349114 172204 349120
rect 173164 349172 173216 349178
rect 173164 349114 173216 349120
rect 172164 345098 172192 349114
rect 170404 345092 170456 345098
rect 170404 345034 170456 345040
rect 172152 345092 172204 345098
rect 172152 345034 172204 345040
rect 170416 330410 170444 345034
rect 167644 330404 167696 330410
rect 167644 330346 167696 330352
rect 170404 330404 170456 330410
rect 170404 330346 170456 330352
rect 167656 322998 167684 330346
rect 165620 322992 165672 322998
rect 165620 322934 165672 322940
rect 167644 322992 167696 322998
rect 167644 322934 167696 322940
rect 165632 320482 165660 322934
rect 231136 321638 231164 349454
rect 231124 321632 231176 321638
rect 231124 321574 231176 321580
rect 228364 321564 228416 321570
rect 228364 321506 228416 321512
rect 162124 320476 162176 320482
rect 162124 320418 162176 320424
rect 165620 320476 165672 320482
rect 165620 320418 165672 320424
rect 162136 307834 162164 320418
rect 228376 307834 228404 321506
rect 160100 307828 160152 307834
rect 160100 307770 160152 307776
rect 162124 307828 162176 307834
rect 162124 307770 162176 307776
rect 228364 307828 228416 307834
rect 228364 307770 228416 307776
rect 160112 305046 160140 307770
rect 221464 307760 221516 307766
rect 221464 307702 221516 307708
rect 160100 305040 160152 305046
rect 160100 304982 160152 304988
rect 157984 302252 158036 302258
rect 157984 302194 158036 302200
rect 155880 300886 156000 300914
rect 155880 298586 155908 300886
rect 221476 299470 221504 307702
rect 220084 299464 220136 299470
rect 220084 299406 220136 299412
rect 221464 299464 221516 299470
rect 221464 299406 221516 299412
rect 155868 298580 155920 298586
rect 155868 298522 155920 298528
rect 155224 295996 155276 296002
rect 155224 295938 155276 295944
rect 151084 294092 151136 294098
rect 151084 294034 151136 294040
rect 152004 294092 152056 294098
rect 152004 294034 152056 294040
rect 146944 292596 146996 292602
rect 146944 292538 146996 292544
rect 150440 292596 150492 292602
rect 150440 292538 150492 292544
rect 91836 289808 91888 289814
rect 91836 289750 91888 289756
rect 93124 289808 93176 289814
rect 93124 289750 93176 289756
rect 91848 280226 91876 289750
rect 146956 282198 146984 292538
rect 135904 282192 135956 282198
rect 135904 282134 135956 282140
rect 146944 282192 146996 282198
rect 146944 282134 146996 282140
rect 91836 280220 91888 280226
rect 91836 280162 91888 280168
rect 88984 280152 89036 280158
rect 88984 280094 89036 280100
rect 88996 258738 89024 280094
rect 135916 262886 135944 282134
rect 151096 269074 151124 294034
rect 220096 274786 220124 299406
rect 218060 274780 218112 274786
rect 218060 274722 218112 274728
rect 220084 274780 220136 274786
rect 220084 274722 220136 274728
rect 218072 271114 218100 274722
rect 215944 271108 215996 271114
rect 215944 271050 215996 271056
rect 218060 271108 218112 271114
rect 218060 271050 218112 271056
rect 149060 269068 149112 269074
rect 149060 269010 149112 269016
rect 151084 269068 151136 269074
rect 151084 269010 151136 269016
rect 149072 262954 149100 269010
rect 146944 262948 146996 262954
rect 146944 262890 146996 262896
rect 149060 262948 149112 262954
rect 149060 262890 149112 262896
rect 121460 262880 121512 262886
rect 121460 262822 121512 262828
rect 135904 262880 135956 262886
rect 135904 262822 135956 262828
rect 121472 258738 121500 262822
rect 81716 258732 81768 258738
rect 81716 258674 81768 258680
rect 88984 258732 89036 258738
rect 88984 258674 89036 258680
rect 117228 258732 117280 258738
rect 117228 258674 117280 258680
rect 121460 258732 121512 258738
rect 121460 258674 121512 258680
rect 81728 253978 81756 258674
rect 117240 253978 117268 258674
rect 146956 253978 146984 262890
rect 215956 256766 215984 271050
rect 215944 256760 215996 256766
rect 215944 256702 215996 256708
rect 210424 256692 210476 256698
rect 210424 256634 210476 256640
rect 210436 253978 210464 256634
rect 79324 253972 79376 253978
rect 79324 253914 79376 253920
rect 81716 253972 81768 253978
rect 81716 253914 81768 253920
rect 113824 253972 113876 253978
rect 113824 253914 113876 253920
rect 117228 253972 117280 253978
rect 117228 253914 117280 253920
rect 145564 253972 145616 253978
rect 145564 253914 145616 253920
rect 146944 253972 146996 253978
rect 146944 253914 146996 253920
rect 209044 253972 209096 253978
rect 209044 253914 209096 253920
rect 210424 253972 210476 253978
rect 210424 253914 210476 253920
rect 71780 251864 71832 251870
rect 71780 251806 71832 251812
rect 79336 247110 79364 253914
rect 113836 247722 113864 253914
rect 97264 247716 97316 247722
rect 97264 247658 97316 247664
rect 113824 247716 113876 247722
rect 113824 247658 113876 247664
rect 76196 247104 76248 247110
rect 76196 247046 76248 247052
rect 79324 247104 79376 247110
rect 79324 247046 79376 247052
rect 49700 245676 49752 245682
rect 49700 245618 49752 245624
rect 51724 245676 51776 245682
rect 51724 245618 51776 245624
rect 49712 242978 49740 245618
rect 49620 242950 49740 242978
rect 49620 241466 49648 242950
rect 49608 241460 49660 241466
rect 49608 241402 49660 241408
rect 47676 241392 47728 241398
rect 47676 241334 47728 241340
rect 47584 241324 47636 241330
rect 47584 241266 47636 241272
rect 76208 240922 76236 247046
rect 46848 240916 46900 240922
rect 46848 240858 46900 240864
rect 76196 240916 76248 240922
rect 76196 240858 76248 240864
rect 46860 239766 46888 240858
rect 46848 239760 46900 239766
rect 46848 239702 46900 239708
rect 97276 239426 97304 247658
rect 145576 247110 145604 253914
rect 143172 247104 143224 247110
rect 143172 247046 143224 247052
rect 145564 247104 145616 247110
rect 145564 247046 145616 247052
rect 143184 242962 143212 247046
rect 143172 242956 143224 242962
rect 143172 242898 143224 242904
rect 136088 242888 136140 242894
rect 136088 242830 136140 242836
rect 136100 240854 136128 242830
rect 136088 240848 136140 240854
rect 136088 240790 136140 240796
rect 209056 240786 209084 253914
rect 209044 240780 209096 240786
rect 209044 240722 209096 240728
rect 395356 240145 395384 665178
rect 395528 646536 395580 646542
rect 395528 646478 395580 646484
rect 395436 562692 395488 562698
rect 395436 562634 395488 562640
rect 395342 240136 395398 240145
rect 395448 240106 395476 562634
rect 395342 240071 395398 240080
rect 395436 240100 395488 240106
rect 395436 240042 395488 240048
rect 395540 240009 395568 646478
rect 396724 378208 396776 378214
rect 396724 378150 396776 378156
rect 396540 240100 396592 240106
rect 396540 240042 396592 240048
rect 395526 240000 395582 240009
rect 395526 239935 395582 239944
rect 97264 239420 97316 239426
rect 97264 239362 97316 239368
rect 396552 238882 396580 240042
rect 396540 238876 396592 238882
rect 396540 238818 396592 238824
rect 396540 238740 396592 238746
rect 396540 238682 396592 238688
rect 45836 232892 45888 232898
rect 45836 232834 45888 232840
rect 45744 232824 45796 232830
rect 45744 232766 45796 232772
rect 45756 230450 45784 232766
rect 64144 232416 64196 232422
rect 64144 232358 64196 232364
rect 85764 232416 85816 232422
rect 85764 232358 85816 232364
rect 392582 232384 392638 232393
rect 46848 231940 46900 231946
rect 46848 231882 46900 231888
rect 46664 231872 46716 231878
rect 46664 231814 46716 231820
rect 46860 231826 46888 231882
rect 45744 230444 45796 230450
rect 45744 230386 45796 230392
rect 46676 229090 46704 231814
rect 46860 231798 46980 231826
rect 46664 229084 46716 229090
rect 46664 229026 46716 229032
rect 46204 227724 46256 227730
rect 46204 227666 46256 227672
rect 46216 223310 46244 227666
rect 46952 224398 46980 231798
rect 48320 231804 48372 231810
rect 48320 231746 48372 231752
rect 48332 229158 48360 231746
rect 60740 231124 60792 231130
rect 60740 231066 60792 231072
rect 51908 230444 51960 230450
rect 51908 230386 51960 230392
rect 48320 229152 48372 229158
rect 48320 229094 48372 229100
rect 48228 229084 48280 229090
rect 48228 229026 48280 229032
rect 46940 224392 46992 224398
rect 46940 224334 46992 224340
rect 46204 223304 46256 223310
rect 46204 223246 46256 223252
rect 47676 223304 47728 223310
rect 47676 223246 47728 223252
rect 46940 221128 46992 221134
rect 46940 221070 46992 221076
rect 45652 217320 45704 217326
rect 45652 217262 45704 217268
rect 46952 216714 46980 221070
rect 47688 218074 47716 223246
rect 48240 222154 48268 229026
rect 51920 227798 51948 230386
rect 55864 229084 55916 229090
rect 55864 229026 55916 229032
rect 51908 227792 51960 227798
rect 51908 227734 51960 227740
rect 50344 224392 50396 224398
rect 50344 224334 50396 224340
rect 48228 222148 48280 222154
rect 48228 222090 48280 222096
rect 47676 218068 47728 218074
rect 47676 218010 47728 218016
rect 46940 216708 46992 216714
rect 46940 216650 46992 216656
rect 50356 198014 50384 224334
rect 55876 224194 55904 229026
rect 55864 224188 55916 224194
rect 55864 224130 55916 224136
rect 51448 222148 51500 222154
rect 51448 222090 51500 222096
rect 51460 213926 51488 222090
rect 53840 218000 53892 218006
rect 53840 217942 53892 217948
rect 51724 216708 51776 216714
rect 51724 216650 51776 216656
rect 51448 213920 51500 213926
rect 51448 213862 51500 213868
rect 51736 200802 51764 216650
rect 53852 211206 53880 217942
rect 54484 213920 54536 213926
rect 54484 213862 54536 213868
rect 53840 211200 53892 211206
rect 53840 211142 53892 211148
rect 54496 208214 54524 213862
rect 54484 208208 54536 208214
rect 54484 208150 54536 208156
rect 55864 208208 55916 208214
rect 55864 208150 55916 208156
rect 51724 200796 51776 200802
rect 51724 200738 51776 200744
rect 50344 198008 50396 198014
rect 50344 197950 50396 197956
rect 53840 198008 53892 198014
rect 53840 197950 53892 197956
rect 53852 192506 53880 197950
rect 53840 192500 53892 192506
rect 53840 192442 53892 192448
rect 55876 177206 55904 208150
rect 56612 195838 56640 230588
rect 60752 230178 60780 231066
rect 60740 230172 60792 230178
rect 60740 230114 60792 230120
rect 62764 230172 62816 230178
rect 62764 230114 62816 230120
rect 60004 227724 60056 227730
rect 60004 227666 60056 227672
rect 60016 224194 60044 227666
rect 57244 224188 57296 224194
rect 57244 224130 57296 224136
rect 60004 224188 60056 224194
rect 60004 224130 60056 224136
rect 62120 224188 62172 224194
rect 62120 224130 62172 224136
rect 57256 215830 57284 224130
rect 62132 221270 62160 224130
rect 62776 221474 62804 230114
rect 64156 227118 64184 232358
rect 85776 230722 85804 232358
rect 392582 232319 392638 232328
rect 380162 231160 380218 231169
rect 380162 231095 380218 231104
rect 85764 230716 85816 230722
rect 85764 230658 85816 230664
rect 93768 230716 93820 230722
rect 93768 230658 93820 230664
rect 64144 227112 64196 227118
rect 64144 227054 64196 227060
rect 62764 221468 62816 221474
rect 62764 221410 62816 221416
rect 69020 221468 69072 221474
rect 69020 221410 69072 221416
rect 62120 221264 62172 221270
rect 62120 221206 62172 221212
rect 66260 221264 66312 221270
rect 66260 221206 66312 221212
rect 58256 217320 58308 217326
rect 58256 217262 58308 217268
rect 57244 215824 57296 215830
rect 57244 215766 57296 215772
rect 58268 212498 58296 217262
rect 66272 216714 66300 221206
rect 69032 219502 69060 221410
rect 69020 219496 69072 219502
rect 69020 219438 69072 219444
rect 72424 219428 72476 219434
rect 72424 219370 72476 219376
rect 66260 216708 66312 216714
rect 66260 216650 66312 216656
rect 68284 216708 68336 216714
rect 68284 216650 68336 216656
rect 58716 215824 58768 215830
rect 58716 215766 58768 215772
rect 58728 213926 58756 215766
rect 58716 213920 58768 213926
rect 58716 213862 58768 213868
rect 60004 213920 60056 213926
rect 60004 213862 60056 213868
rect 58256 212492 58308 212498
rect 58256 212434 58308 212440
rect 56692 211132 56744 211138
rect 56692 211074 56744 211080
rect 56704 207806 56732 211074
rect 56692 207800 56744 207806
rect 56692 207742 56744 207748
rect 60016 206990 60044 213862
rect 61936 212492 61988 212498
rect 61936 212434 61988 212440
rect 60004 206984 60056 206990
rect 60004 206926 60056 206932
rect 61948 204950 61976 212434
rect 62028 207800 62080 207806
rect 62028 207742 62080 207748
rect 62040 206938 62068 207742
rect 66168 206984 66220 206990
rect 62040 206910 62160 206938
rect 66168 206926 66220 206932
rect 61936 204944 61988 204950
rect 61936 204886 61988 204892
rect 62132 204270 62160 206910
rect 62120 204264 62172 204270
rect 62120 204206 62172 204212
rect 64144 204264 64196 204270
rect 64144 204206 64196 204212
rect 64156 195974 64184 204206
rect 66180 200114 66208 206926
rect 66180 200086 66484 200114
rect 66456 199442 66484 200086
rect 66444 199436 66496 199442
rect 66444 199378 66496 199384
rect 68296 197402 68324 216650
rect 72436 215286 72464 219370
rect 72424 215280 72476 215286
rect 72424 215222 72476 215228
rect 75184 215280 75236 215286
rect 75184 215222 75236 215228
rect 71044 204944 71096 204950
rect 71044 204886 71096 204892
rect 68284 197396 68336 197402
rect 68284 197338 68336 197344
rect 64144 195968 64196 195974
rect 64144 195910 64196 195916
rect 65524 195968 65576 195974
rect 65524 195910 65576 195916
rect 56600 195832 56652 195838
rect 56600 195774 56652 195780
rect 60372 192500 60424 192506
rect 60372 192442 60424 192448
rect 60384 189106 60412 192442
rect 60372 189100 60424 189106
rect 60372 189042 60424 189048
rect 62764 189100 62816 189106
rect 62764 189042 62816 189048
rect 62776 180062 62804 189042
rect 65536 182170 65564 195910
rect 65524 182164 65576 182170
rect 65524 182106 65576 182112
rect 66904 182164 66956 182170
rect 66904 182106 66956 182112
rect 62764 180056 62816 180062
rect 62764 179998 62816 180004
rect 63776 180056 63828 180062
rect 63776 179998 63828 180004
rect 63788 178022 63816 179998
rect 63776 178016 63828 178022
rect 63776 177958 63828 177964
rect 65524 178016 65576 178022
rect 65524 177958 65576 177964
rect 55864 177200 55916 177206
rect 55864 177142 55916 177148
rect 56876 177200 56928 177206
rect 56876 177142 56928 177148
rect 56888 175302 56916 177142
rect 56876 175296 56928 175302
rect 56876 175238 56928 175244
rect 62120 175228 62172 175234
rect 62120 175170 62172 175176
rect 62132 173058 62160 175170
rect 62120 173052 62172 173058
rect 62120 172994 62172 173000
rect 65248 173052 65300 173058
rect 65248 172994 65300 173000
rect 45560 172508 45612 172514
rect 45560 172450 45612 172456
rect 46940 172508 46992 172514
rect 46940 172450 46992 172456
rect 46952 169046 46980 172450
rect 46940 169040 46992 169046
rect 46940 168982 46992 168988
rect 50988 169040 51040 169046
rect 50988 168982 51040 168988
rect 51000 162178 51028 168982
rect 65260 165578 65288 172994
rect 65248 165572 65300 165578
rect 65248 165514 65300 165520
rect 65536 165510 65564 177958
rect 65524 165504 65576 165510
rect 65524 165446 65576 165452
rect 50988 162172 51040 162178
rect 50988 162114 51040 162120
rect 60556 162172 60608 162178
rect 60556 162114 60608 162120
rect 60568 159050 60596 162114
rect 60556 159044 60608 159050
rect 60556 158986 60608 158992
rect 66916 141302 66944 182106
rect 71056 180130 71084 204886
rect 75196 202910 75224 215222
rect 75184 202904 75236 202910
rect 75184 202846 75236 202852
rect 80704 202836 80756 202842
rect 80704 202778 80756 202784
rect 73160 200796 73212 200802
rect 73160 200738 73212 200744
rect 73172 198014 73200 200738
rect 75460 199436 75512 199442
rect 75460 199378 75512 199384
rect 73160 198008 73212 198014
rect 73160 197950 73212 197956
rect 71780 197328 71832 197334
rect 71780 197270 71832 197276
rect 71792 194546 71820 197270
rect 75472 194546 75500 199378
rect 77944 198008 77996 198014
rect 77944 197950 77996 197956
rect 71780 194540 71832 194546
rect 71780 194482 71832 194488
rect 75184 194540 75236 194546
rect 75184 194482 75236 194488
rect 75460 194540 75512 194546
rect 75460 194482 75512 194488
rect 76564 194540 76616 194546
rect 76564 194482 76616 194488
rect 71044 180124 71096 180130
rect 71044 180066 71096 180072
rect 68284 165572 68336 165578
rect 68284 165514 68336 165520
rect 66996 159044 67048 159050
rect 66996 158986 67048 158992
rect 67008 153202 67036 158986
rect 66996 153196 67048 153202
rect 66996 153138 67048 153144
rect 68296 146266 68324 165514
rect 73804 165504 73856 165510
rect 73804 165446 73856 165452
rect 73816 158710 73844 165446
rect 73804 158704 73856 158710
rect 73804 158646 73856 158652
rect 71044 153196 71096 153202
rect 71044 153138 71096 153144
rect 68284 146260 68336 146266
rect 68284 146202 68336 146208
rect 69664 146260 69716 146266
rect 69664 146202 69716 146208
rect 69676 143546 69704 146202
rect 69664 143540 69716 143546
rect 69664 143482 69716 143488
rect 71056 143070 71084 153138
rect 75196 143546 75224 194482
rect 76576 188630 76604 194482
rect 76564 188624 76616 188630
rect 76564 188566 76616 188572
rect 76748 158704 76800 158710
rect 76748 158646 76800 158652
rect 76760 155990 76788 158646
rect 76748 155984 76800 155990
rect 76748 155926 76800 155932
rect 77956 151094 77984 197950
rect 79968 188624 80020 188630
rect 79968 188566 80020 188572
rect 79980 186386 80008 188566
rect 80716 187950 80744 202778
rect 86972 195906 87000 230588
rect 93780 228970 93808 230658
rect 93780 228942 93900 228970
rect 93872 226506 93900 228942
rect 117240 228410 117268 230588
rect 146312 230574 146510 230602
rect 117228 228404 117280 228410
rect 117228 228346 117280 228352
rect 138664 228404 138716 228410
rect 138664 228346 138716 228352
rect 95884 227112 95936 227118
rect 95884 227054 95936 227060
rect 93860 226500 93912 226506
rect 93860 226442 93912 226448
rect 95896 218754 95924 227054
rect 98000 226500 98052 226506
rect 98000 226442 98052 226448
rect 98012 224194 98040 226442
rect 98000 224188 98052 224194
rect 98000 224130 98052 224136
rect 100024 224188 100076 224194
rect 100024 224130 100076 224136
rect 95884 218748 95936 218754
rect 95884 218690 95936 218696
rect 100036 218006 100064 224130
rect 106188 218748 106240 218754
rect 106188 218690 106240 218696
rect 100024 218000 100076 218006
rect 100024 217942 100076 217948
rect 106004 218000 106056 218006
rect 106004 217942 106056 217948
rect 106016 215354 106044 217942
rect 106004 215348 106056 215354
rect 106004 215290 106056 215296
rect 106200 214674 106228 218690
rect 115848 218068 115900 218074
rect 115848 218010 115900 218016
rect 110420 215280 110472 215286
rect 110420 215222 110472 215228
rect 106188 214668 106240 214674
rect 106188 214610 106240 214616
rect 107844 214668 107896 214674
rect 107844 214610 107896 214616
rect 107856 210458 107884 214610
rect 110432 210526 110460 215222
rect 110420 210520 110472 210526
rect 110420 210462 110472 210468
rect 113180 210520 113232 210526
rect 113180 210462 113232 210468
rect 107844 210452 107896 210458
rect 107844 210394 107896 210400
rect 113192 206038 113220 210462
rect 113180 206032 113232 206038
rect 113180 205974 113232 205980
rect 115112 206032 115164 206038
rect 115112 205974 115164 205980
rect 115124 201482 115152 205974
rect 115112 201476 115164 201482
rect 115112 201418 115164 201424
rect 86960 195900 87012 195906
rect 86960 195842 87012 195848
rect 80704 187944 80756 187950
rect 80704 187886 80756 187892
rect 82176 187944 82228 187950
rect 82176 187886 82228 187892
rect 79968 186380 80020 186386
rect 79968 186322 80020 186328
rect 82188 183530 82216 187886
rect 112444 187740 112496 187746
rect 112444 187682 112496 187688
rect 86224 186312 86276 186318
rect 86224 186254 86276 186260
rect 82176 183524 82228 183530
rect 82176 183466 82228 183472
rect 83556 183524 83608 183530
rect 83556 183466 83608 183472
rect 81440 180124 81492 180130
rect 81440 180066 81492 180072
rect 81452 175234 81480 180066
rect 83568 176662 83596 183466
rect 83556 176656 83608 176662
rect 83556 176598 83608 176604
rect 84936 176656 84988 176662
rect 84936 176598 84988 176604
rect 81440 175228 81492 175234
rect 81440 175170 81492 175176
rect 84844 175228 84896 175234
rect 84844 175170 84896 175176
rect 84856 167686 84884 175170
rect 84948 170134 84976 176598
rect 84936 170128 84988 170134
rect 84936 170070 84988 170076
rect 84844 167680 84896 167686
rect 84844 167622 84896 167628
rect 86236 165578 86264 186254
rect 88248 170128 88300 170134
rect 88248 170070 88300 170076
rect 87696 167680 87748 167686
rect 87696 167622 87748 167628
rect 86224 165572 86276 165578
rect 86224 165514 86276 165520
rect 87708 164218 87736 167622
rect 88260 167074 88288 170070
rect 88248 167068 88300 167074
rect 88248 167010 88300 167016
rect 91100 167000 91152 167006
rect 91100 166942 91152 166948
rect 88984 165572 89036 165578
rect 88984 165514 89036 165520
rect 87696 164212 87748 164218
rect 87696 164154 87748 164160
rect 84844 155916 84896 155922
rect 84844 155858 84896 155864
rect 84856 153270 84884 155858
rect 84844 153264 84896 153270
rect 84844 153206 84896 153212
rect 87604 153196 87656 153202
rect 87604 153138 87656 153144
rect 77944 151088 77996 151094
rect 77944 151030 77996 151036
rect 81440 151088 81492 151094
rect 81440 151030 81492 151036
rect 81452 145586 81480 151030
rect 81440 145580 81492 145586
rect 81440 145522 81492 145528
rect 71136 143540 71188 143546
rect 71136 143482 71188 143488
rect 75184 143540 75236 143546
rect 75184 143482 75236 143488
rect 76564 143540 76616 143546
rect 76564 143482 76616 143488
rect 71044 143064 71096 143070
rect 71044 143006 71096 143012
rect 66904 141296 66956 141302
rect 66904 141238 66956 141244
rect 68376 141296 68428 141302
rect 68376 141238 68428 141244
rect 68388 137902 68416 141238
rect 68376 137896 68428 137902
rect 68376 137838 68428 137844
rect 69664 137896 69716 137902
rect 69664 137838 69716 137844
rect 69676 120018 69704 137838
rect 71148 135250 71176 143482
rect 71136 135244 71188 135250
rect 71136 135186 71188 135192
rect 72424 135244 72476 135250
rect 72424 135186 72476 135192
rect 72436 121514 72464 135186
rect 76576 127634 76604 143482
rect 76656 143064 76708 143070
rect 76656 143006 76708 143012
rect 76668 133210 76696 143006
rect 87616 134774 87644 153138
rect 88996 151570 89024 165514
rect 91112 164218 91140 166942
rect 90364 164212 90416 164218
rect 90364 164154 90416 164160
rect 91100 164212 91152 164218
rect 91100 164154 91152 164160
rect 93124 164212 93176 164218
rect 93124 164154 93176 164160
rect 88984 151564 89036 151570
rect 88984 151506 89036 151512
rect 90376 138038 90404 164154
rect 93136 151842 93164 164154
rect 93124 151836 93176 151842
rect 93124 151778 93176 151784
rect 95240 151768 95292 151774
rect 95240 151710 95292 151716
rect 90456 151564 90508 151570
rect 90456 151506 90508 151512
rect 90364 138032 90416 138038
rect 90364 137974 90416 137980
rect 90468 137970 90496 151506
rect 95252 146266 95280 151710
rect 95240 146260 95292 146266
rect 95240 146202 95292 146208
rect 97264 146260 97316 146266
rect 97264 146202 97316 146208
rect 91744 145580 91796 145586
rect 91744 145522 91796 145528
rect 91756 141574 91784 145522
rect 91744 141568 91796 141574
rect 91744 141510 91796 141516
rect 94044 141568 94096 141574
rect 94044 141510 94096 141516
rect 93124 138032 93176 138038
rect 93124 137974 93176 137980
rect 90456 137964 90508 137970
rect 90456 137906 90508 137912
rect 87604 134768 87656 134774
rect 87604 134710 87656 134716
rect 76656 133204 76708 133210
rect 76656 133146 76708 133152
rect 86224 133204 86276 133210
rect 86224 133146 86276 133152
rect 76564 127628 76616 127634
rect 76564 127570 76616 127576
rect 79324 127628 79376 127634
rect 79324 127570 79376 127576
rect 72424 121508 72476 121514
rect 72424 121450 72476 121456
rect 73804 121508 73856 121514
rect 73804 121450 73856 121456
rect 69664 120012 69716 120018
rect 69664 119954 69716 119960
rect 70492 120012 70544 120018
rect 70492 119954 70544 119960
rect 70504 118590 70532 119954
rect 70492 118584 70544 118590
rect 70492 118526 70544 118532
rect 73816 98666 73844 121450
rect 76288 118584 76340 118590
rect 76288 118526 76340 118532
rect 76300 116074 76328 118526
rect 79336 118318 79364 127570
rect 86236 121514 86264 133146
rect 93136 128314 93164 137974
rect 94056 135930 94084 141510
rect 94688 137964 94740 137970
rect 94688 137906 94740 137912
rect 94044 135924 94096 135930
rect 94044 135866 94096 135872
rect 94700 133890 94728 137906
rect 94688 133884 94740 133890
rect 94688 133826 94740 133832
rect 95608 133884 95660 133890
rect 95608 133826 95660 133832
rect 95620 131782 95648 133826
rect 95608 131776 95660 131782
rect 95608 131718 95660 131724
rect 97276 131646 97304 146202
rect 105544 135924 105596 135930
rect 105544 135866 105596 135872
rect 97540 131776 97592 131782
rect 97540 131718 97592 131724
rect 97264 131640 97316 131646
rect 97264 131582 97316 131588
rect 93124 128308 93176 128314
rect 93124 128250 93176 128256
rect 95884 128308 95936 128314
rect 95884 128250 95936 128256
rect 86224 121508 86276 121514
rect 86224 121450 86276 121456
rect 88984 121508 89036 121514
rect 88984 121450 89036 121456
rect 79324 118312 79376 118318
rect 79324 118254 79376 118260
rect 81164 118312 81216 118318
rect 81164 118254 81216 118260
rect 76288 116068 76340 116074
rect 76288 116010 76340 116016
rect 77944 116068 77996 116074
rect 77944 116010 77996 116016
rect 77956 112334 77984 116010
rect 81176 114510 81204 118254
rect 81164 114504 81216 114510
rect 81164 114446 81216 114452
rect 82820 114504 82872 114510
rect 82820 114446 82872 114452
rect 77944 112328 77996 112334
rect 77944 112270 77996 112276
rect 79968 112328 80020 112334
rect 79968 112270 80020 112276
rect 79980 111738 80008 112270
rect 79980 111710 80100 111738
rect 80072 107642 80100 111710
rect 82832 111110 82860 114446
rect 82820 111104 82872 111110
rect 82820 111046 82872 111052
rect 88248 111104 88300 111110
rect 88248 111046 88300 111052
rect 80060 107636 80112 107642
rect 80060 107578 80112 107584
rect 88260 104922 88288 111046
rect 88248 104916 88300 104922
rect 88248 104858 88300 104864
rect 88996 103902 89024 121450
rect 95896 112470 95924 128250
rect 97552 124098 97580 131718
rect 99288 131640 99340 131646
rect 99288 131582 99340 131588
rect 99300 128330 99328 131582
rect 99300 128302 99420 128330
rect 99392 126886 99420 128302
rect 105556 127634 105584 135866
rect 105544 127628 105596 127634
rect 105544 127570 105596 127576
rect 111064 127628 111116 127634
rect 111064 127570 111116 127576
rect 99380 126880 99432 126886
rect 99380 126822 99432 126828
rect 101496 126880 101548 126886
rect 101496 126822 101548 126828
rect 97540 124092 97592 124098
rect 97540 124034 97592 124040
rect 99288 124092 99340 124098
rect 99288 124034 99340 124040
rect 99300 122834 99328 124034
rect 99300 122806 99420 122834
rect 99392 121310 99420 122806
rect 101508 121378 101536 126822
rect 101496 121372 101548 121378
rect 101496 121314 101548 121320
rect 104900 121372 104952 121378
rect 104900 121314 104952 121320
rect 99380 121304 99432 121310
rect 99380 121246 99432 121252
rect 102048 121304 102100 121310
rect 102048 121246 102100 121252
rect 102060 115818 102088 121246
rect 104912 119678 104940 121314
rect 104900 119672 104952 119678
rect 104900 119614 104952 119620
rect 106924 119672 106976 119678
rect 106924 119614 106976 119620
rect 102060 115790 102180 115818
rect 95884 112464 95936 112470
rect 95884 112406 95936 112412
rect 102152 107574 102180 115790
rect 102140 107568 102192 107574
rect 102140 107510 102192 107516
rect 106188 107568 106240 107574
rect 106188 107510 106240 107516
rect 106200 106282 106228 107510
rect 106188 106276 106240 106282
rect 106188 106218 106240 106224
rect 106936 104786 106964 119614
rect 108304 112464 108356 112470
rect 108304 112406 108356 112412
rect 108316 109002 108344 112406
rect 108304 108996 108356 109002
rect 108304 108938 108356 108944
rect 106924 104780 106976 104786
rect 106924 104722 106976 104728
rect 108396 104780 108448 104786
rect 108396 104722 108448 104728
rect 88984 103896 89036 103902
rect 88984 103838 89036 103844
rect 95240 103896 95292 103902
rect 95240 103838 95292 103844
rect 95252 98734 95280 103838
rect 95240 98728 95292 98734
rect 95240 98670 95292 98676
rect 98644 98728 98696 98734
rect 98644 98670 98696 98676
rect 73804 98660 73856 98666
rect 73804 98602 73856 98608
rect 77944 98660 77996 98666
rect 77944 98602 77996 98608
rect 77956 87038 77984 98602
rect 77944 87032 77996 87038
rect 77944 86974 77996 86980
rect 83556 86964 83608 86970
rect 83556 86906 83608 86912
rect 83568 80034 83596 86906
rect 98656 82890 98684 98670
rect 108408 96694 108436 104722
rect 108396 96688 108448 96694
rect 108396 96630 108448 96636
rect 110972 96620 111024 96626
rect 110972 96562 111024 96568
rect 110984 88330 111012 96562
rect 110972 88324 111024 88330
rect 110972 88266 111024 88272
rect 98644 82884 98696 82890
rect 98644 82826 98696 82832
rect 104164 82884 104216 82890
rect 104164 82826 104216 82832
rect 83556 80028 83608 80034
rect 83556 79970 83608 79976
rect 84844 80028 84896 80034
rect 84844 79970 84896 79976
rect 44824 73636 44876 73642
rect 44824 73578 44876 73584
rect 84856 73234 84884 79970
rect 84844 73228 84896 73234
rect 84844 73170 84896 73176
rect 92480 73160 92532 73166
rect 92480 73102 92532 73108
rect 22742 72584 22798 72593
rect 22742 72519 22798 72528
rect 60740 72548 60792 72554
rect 6920 71664 6972 71670
rect 6920 71606 6972 71612
rect 5540 66904 5592 66910
rect 5540 66846 5592 66852
rect 3606 58576 3662 58585
rect 3606 58511 3662 58520
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 3516 22704 3568 22710
rect 3516 22646 3568 22652
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3528 6497 3556 22646
rect 5552 16574 5580 66846
rect 15200 54528 15252 54534
rect 15200 54470 15252 54476
rect 15212 16574 15240 54470
rect 5552 16546 6040 16574
rect 15212 16546 15976 16574
rect 3514 6488 3570 6497
rect 3514 6423 3570 6432
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 2872 3460 2924 3466
rect 570 3360 626 3369
rect 570 3295 626 3304
rect 584 480 612 3295
rect 1688 480 1716 3431
rect 2872 3402 2924 3408
rect 2884 480 2912 3402
rect 4080 480 4108 6122
rect 5264 4888 5316 4894
rect 5264 4830 5316 4836
rect 5276 480 5304 4830
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6012 354 6040 16546
rect 14280 13116 14332 13122
rect 14280 13058 14332 13064
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7668 480 7696 3470
rect 8772 480 8800 6190
rect 9968 480 9996 8910
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11164 480 11192 6598
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12360 480 12388 3538
rect 13556 480 13584 6258
rect 6430 354 6542 480
rect 6012 326 6542 354
rect 6430 -960 6542 326
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 13058
rect 15948 480 15976 16546
rect 19432 7676 19484 7682
rect 19432 7618 19484 7624
rect 18234 6216 18290 6225
rect 18234 6151 18290 6160
rect 17038 3632 17094 3641
rect 17038 3567 17094 3576
rect 17052 480 17080 3567
rect 18248 480 18276 6151
rect 19444 480 19472 7618
rect 22756 4894 22784 72519
rect 60740 72490 60792 72496
rect 25504 72480 25556 72486
rect 25504 72422 25556 72428
rect 25320 10328 25372 10334
rect 25320 10270 25372 10276
rect 24216 9036 24268 9042
rect 24216 8978 24268 8984
rect 23020 7608 23072 7614
rect 23020 7550 23072 7556
rect 22744 4888 22796 4894
rect 22744 4830 22796 4836
rect 21824 4820 21876 4826
rect 21824 4762 21876 4768
rect 20628 3256 20680 3262
rect 20628 3198 20680 3204
rect 20640 480 20668 3198
rect 21836 480 21864 4762
rect 23032 480 23060 7550
rect 24228 480 24256 8978
rect 25332 480 25360 10270
rect 25516 3262 25544 72422
rect 35900 18624 35952 18630
rect 35900 18566 35952 18572
rect 35912 16574 35940 18566
rect 60752 16574 60780 72490
rect 86224 72276 86276 72282
rect 86224 72218 86276 72224
rect 81440 25560 81492 25566
rect 81440 25502 81492 25508
rect 81452 16574 81480 25502
rect 35912 16546 36032 16574
rect 60752 16546 61608 16574
rect 81452 16546 81664 16574
rect 31944 10396 31996 10402
rect 31944 10338 31996 10344
rect 31300 9104 31352 9110
rect 31300 9046 31352 9052
rect 27712 7744 27764 7750
rect 27712 7686 27764 7692
rect 26516 4888 26568 4894
rect 26516 4830 26568 4836
rect 25504 3256 25556 3262
rect 25504 3198 25556 3204
rect 26528 480 26556 4830
rect 27724 480 27752 7686
rect 30104 6384 30156 6390
rect 30104 6326 30156 6332
rect 28908 4956 28960 4962
rect 28908 4898 28960 4904
rect 28920 480 28948 4898
rect 30116 480 30144 6326
rect 31312 480 31340 9046
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 31956 354 31984 10338
rect 34794 8936 34850 8945
rect 34794 8871 34850 8880
rect 33600 5024 33652 5030
rect 33600 4966 33652 4972
rect 33612 480 33640 4966
rect 34808 480 34836 8871
rect 36004 480 36032 16546
rect 46664 10464 46716 10470
rect 46664 10406 46716 10412
rect 43076 9376 43128 9382
rect 43076 9318 43128 9324
rect 41880 9172 41932 9178
rect 41880 9114 41932 9120
rect 38382 9072 38438 9081
rect 38382 9007 38438 9016
rect 37186 4856 37242 4865
rect 37186 4791 37242 4800
rect 37200 480 37228 4791
rect 38396 480 38424 9007
rect 40684 6452 40736 6458
rect 40684 6394 40736 6400
rect 39580 3664 39632 3670
rect 39580 3606 39632 3612
rect 39592 480 39620 3606
rect 40696 480 40724 6394
rect 41892 480 41920 9114
rect 43088 480 43116 9318
rect 45468 9240 45520 9246
rect 45468 9182 45520 9188
rect 44272 6520 44324 6526
rect 44272 6462 44324 6468
rect 44284 480 44312 6462
rect 45480 480 45508 9182
rect 46676 480 46704 10406
rect 60832 9512 60884 9518
rect 60832 9454 60884 9460
rect 57244 9444 57296 9450
rect 57244 9386 57296 9392
rect 50160 9308 50212 9314
rect 50160 9250 50212 9256
rect 48964 6588 49016 6594
rect 48964 6530 49016 6536
rect 47860 3732 47912 3738
rect 47860 3674 47912 3680
rect 47872 480 47900 3674
rect 48976 480 49004 6530
rect 50172 480 50200 9250
rect 53746 9208 53802 9217
rect 53746 9143 53802 9152
rect 52550 6352 52606 6361
rect 52550 6287 52606 6296
rect 51356 3800 51408 3806
rect 51356 3742 51408 3748
rect 51368 480 51396 3742
rect 52564 480 52592 6287
rect 53760 480 53788 9143
rect 56046 6488 56102 6497
rect 56046 6423 56102 6432
rect 54942 3768 54998 3777
rect 54942 3703 54998 3712
rect 54956 480 54984 3703
rect 56060 480 56088 6423
rect 57256 480 57284 9386
rect 59636 6724 59688 6730
rect 59636 6666 59688 6672
rect 58440 3868 58492 3874
rect 58440 3810 58492 3816
rect 58452 480 58480 3810
rect 59648 480 59676 6666
rect 60844 480 60872 9454
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 75000 10736 75052 10742
rect 75000 10678 75052 10684
rect 67640 10600 67692 10606
rect 67640 10542 67692 10548
rect 64328 10532 64380 10538
rect 64328 10474 64380 10480
rect 63224 7812 63276 7818
rect 63224 7754 63276 7760
rect 63236 480 63264 7754
rect 64340 480 64368 10474
rect 66720 7880 66772 7886
rect 66720 7822 66772 7828
rect 65524 5092 65576 5098
rect 65524 5034 65576 5040
rect 65536 480 65564 5034
rect 66732 480 66760 7822
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 10542
rect 71502 10296 71558 10305
rect 71502 10231 71558 10240
rect 70306 7576 70362 7585
rect 70306 7511 70362 7520
rect 69112 3936 69164 3942
rect 69112 3878 69164 3884
rect 69124 480 69152 3878
rect 70320 480 70348 7511
rect 71516 480 71544 10231
rect 73804 7948 73856 7954
rect 73804 7890 73856 7896
rect 72608 5160 72660 5166
rect 72608 5102 72660 5108
rect 72620 480 72648 5102
rect 73816 480 73844 7890
rect 75012 480 75040 10678
rect 78128 10668 78180 10674
rect 78128 10610 78180 10616
rect 77392 8016 77444 8022
rect 77392 7958 77444 7964
rect 76196 5228 76248 5234
rect 76196 5170 76248 5176
rect 76208 480 76236 5170
rect 77404 480 77432 7958
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78140 354 78168 10610
rect 80888 8084 80940 8090
rect 80888 8026 80940 8032
rect 79692 4004 79744 4010
rect 79692 3946 79744 3952
rect 79704 480 79732 3946
rect 80900 480 80928 8026
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 78558 -960 78670 326
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 84476 8152 84528 8158
rect 84476 8094 84528 8100
rect 83280 4072 83332 4078
rect 83280 4014 83332 4020
rect 83292 480 83320 4014
rect 84488 480 84516 8094
rect 86236 6662 86264 72218
rect 92492 71602 92520 73102
rect 92480 71596 92532 71602
rect 92480 71538 92532 71544
rect 104176 71534 104204 82826
rect 111076 74390 111104 127570
rect 111064 74384 111116 74390
rect 111064 74326 111116 74332
rect 112456 73778 112484 187682
rect 114468 178084 114520 178090
rect 114468 178026 114520 178032
rect 114006 138680 114062 138689
rect 114006 138615 114062 138624
rect 113824 137420 113876 137426
rect 113824 137362 113876 137368
rect 113732 134564 113784 134570
rect 113732 134506 113784 134512
rect 113638 131200 113694 131209
rect 113638 131135 113640 131144
rect 113692 131135 113694 131144
rect 113640 131106 113692 131112
rect 113546 129024 113602 129033
rect 113546 128959 113602 128968
rect 113560 128382 113588 128959
rect 113548 128376 113600 128382
rect 113548 128318 113600 128324
rect 113546 127528 113602 127537
rect 113546 127463 113602 127472
rect 113560 127022 113588 127463
rect 113548 127016 113600 127022
rect 113548 126958 113600 126964
rect 113640 126948 113692 126954
rect 113640 126890 113692 126896
rect 113652 126857 113680 126890
rect 113638 126848 113694 126857
rect 113638 126783 113694 126792
rect 113640 125588 113692 125594
rect 113640 125530 113692 125536
rect 113652 125497 113680 125530
rect 113638 125488 113694 125497
rect 113638 125423 113694 125432
rect 113640 124160 113692 124166
rect 113640 124102 113692 124108
rect 113652 123865 113680 124102
rect 113638 123856 113694 123865
rect 113638 123791 113694 123800
rect 113640 122800 113692 122806
rect 113638 122768 113640 122777
rect 113692 122768 113694 122777
rect 113638 122703 113694 122712
rect 113640 121440 113692 121446
rect 113640 121382 113692 121388
rect 113652 121281 113680 121382
rect 113638 121272 113694 121281
rect 113638 121207 113694 121216
rect 113640 120080 113692 120086
rect 113640 120022 113692 120028
rect 113652 119785 113680 120022
rect 113638 119776 113694 119785
rect 113638 119711 113694 119720
rect 113640 118652 113692 118658
rect 113640 118594 113692 118600
rect 113652 118289 113680 118594
rect 113638 118280 113694 118289
rect 113638 118215 113694 118224
rect 113640 117292 113692 117298
rect 113640 117234 113692 117240
rect 113652 116793 113680 117234
rect 113638 116784 113694 116793
rect 113638 116719 113694 116728
rect 113548 115932 113600 115938
rect 113548 115874 113600 115880
rect 113560 115297 113588 115874
rect 113546 115288 113602 115297
rect 113546 115223 113602 115232
rect 113640 113144 113692 113150
rect 113638 113112 113640 113121
rect 113692 113112 113694 113121
rect 113638 113047 113694 113056
rect 113640 111784 113692 111790
rect 113638 111752 113640 111761
rect 113692 111752 113694 111761
rect 113638 111687 113694 111696
rect 113640 110424 113692 110430
rect 113638 110392 113640 110401
rect 113692 110392 113694 110401
rect 113638 110327 113694 110336
rect 113640 108996 113692 109002
rect 113640 108938 113692 108944
rect 113652 108905 113680 108938
rect 113638 108896 113694 108905
rect 113638 108831 113694 108840
rect 113640 107636 113692 107642
rect 113640 107578 113692 107584
rect 113652 107545 113680 107578
rect 113638 107536 113694 107545
rect 113638 107471 113694 107480
rect 113548 106276 113600 106282
rect 113548 106218 113600 106224
rect 113560 105913 113588 106218
rect 113546 105904 113602 105913
rect 113546 105839 113602 105848
rect 113640 104848 113692 104854
rect 113638 104816 113640 104825
rect 113692 104816 113694 104825
rect 113638 104751 113694 104760
rect 113744 103193 113772 134506
rect 113730 103184 113786 103193
rect 113730 103119 113786 103128
rect 113836 101833 113864 137362
rect 113916 135924 113968 135930
rect 113916 135866 113968 135872
rect 113822 101824 113878 101833
rect 113822 101759 113878 101768
rect 113928 91089 113956 135866
rect 113914 91080 113970 91089
rect 113914 91015 113970 91024
rect 114020 89729 114048 138615
rect 114376 138032 114428 138038
rect 114376 137974 114428 137980
rect 114100 137624 114152 137630
rect 114100 137566 114152 137572
rect 114006 89720 114062 89729
rect 114006 89655 114062 89664
rect 113824 88324 113876 88330
rect 113824 88266 113876 88272
rect 113836 81666 113864 88266
rect 114112 88233 114140 137566
rect 114192 137556 114244 137562
rect 114192 137498 114244 137504
rect 114098 88224 114154 88233
rect 114098 88159 114154 88168
rect 114204 86873 114232 137498
rect 114284 137488 114336 137494
rect 114284 137430 114336 137436
rect 114190 86864 114246 86873
rect 114190 86799 114246 86808
rect 114296 85377 114324 137430
rect 114282 85368 114338 85377
rect 114282 85303 114338 85312
rect 113824 81660 113876 81666
rect 113824 81602 113876 81608
rect 114388 80889 114416 137974
rect 114480 82385 114508 178026
rect 115756 174344 115808 174350
rect 115756 174286 115808 174292
rect 115664 142860 115716 142866
rect 115664 142802 115716 142808
rect 115112 137352 115164 137358
rect 115112 137294 115164 137300
rect 115294 137320 115350 137329
rect 115124 132734 115152 137294
rect 115294 137255 115350 137264
rect 115388 137284 115440 137290
rect 115204 136672 115256 136678
rect 115204 136614 115256 136620
rect 115112 132728 115164 132734
rect 115112 132670 115164 132676
rect 114466 82376 114522 82385
rect 114466 82311 114522 82320
rect 114560 81660 114612 81666
rect 114560 81602 114612 81608
rect 114374 80880 114430 80889
rect 114374 80815 114430 80824
rect 114466 78704 114522 78713
rect 114466 78639 114522 78648
rect 114374 76664 114430 76673
rect 114374 76599 114430 76608
rect 113916 74384 113968 74390
rect 113916 74326 113968 74332
rect 112444 73772 112496 73778
rect 112444 73714 112496 73720
rect 104164 71528 104216 71534
rect 104164 71470 104216 71476
rect 113928 71466 113956 74326
rect 113916 71460 113968 71466
rect 113916 71402 113968 71408
rect 114388 60722 114416 76599
rect 114480 75750 114508 78639
rect 114468 75744 114520 75750
rect 114468 75686 114520 75692
rect 114572 75682 114600 81602
rect 114560 75676 114612 75682
rect 114560 75618 114612 75624
rect 114466 75440 114522 75449
rect 114466 75375 114522 75384
rect 114376 60716 114428 60722
rect 114376 60658 114428 60664
rect 113180 51128 113232 51134
rect 113180 51070 113232 51076
rect 106280 43444 106332 43450
rect 106280 43386 106332 43392
rect 106292 16574 106320 43386
rect 113192 16574 113220 51070
rect 114480 22778 114508 75375
rect 115216 74322 115244 136614
rect 115308 132818 115336 137255
rect 115388 137226 115440 137232
rect 115400 132954 115428 137226
rect 115480 135992 115532 135998
rect 115480 135934 115532 135940
rect 115492 133090 115520 135934
rect 115572 134836 115624 134842
rect 115572 134778 115624 134784
rect 115584 133249 115612 134778
rect 115570 133240 115626 133249
rect 115570 133175 115626 133184
rect 115492 133062 115612 133090
rect 115400 132926 115520 132954
rect 115308 132790 115428 132818
rect 115296 132728 115348 132734
rect 115296 132670 115348 132676
rect 115308 100337 115336 132670
rect 115294 100328 115350 100337
rect 115294 100263 115350 100272
rect 115400 98841 115428 132790
rect 115386 98832 115442 98841
rect 115386 98767 115442 98776
rect 115492 93809 115520 132926
rect 115478 93800 115534 93809
rect 115478 93735 115534 93744
rect 115584 92449 115612 133062
rect 115676 95237 115704 142802
rect 115768 96733 115796 174286
rect 115754 96724 115810 96733
rect 115754 96659 115810 96668
rect 115662 95228 115718 95237
rect 115662 95163 115718 95172
rect 115570 92440 115626 92449
rect 115570 92375 115626 92384
rect 115860 83269 115888 218010
rect 116584 210452 116636 210458
rect 116584 210394 116636 210400
rect 116596 194546 116624 210394
rect 116860 201476 116912 201482
rect 116860 201418 116912 201424
rect 116872 197878 116900 201418
rect 116860 197872 116912 197878
rect 116860 197814 116912 197820
rect 119988 197872 120040 197878
rect 119988 197814 120040 197820
rect 120000 195922 120028 197814
rect 138676 195974 138704 228346
rect 146312 197418 146340 230574
rect 176672 229770 176700 230588
rect 167644 229764 167696 229770
rect 167644 229706 167696 229712
rect 176660 229764 176712 229770
rect 176660 229706 176712 229712
rect 157984 228472 158036 228478
rect 157984 228414 158036 228420
rect 155960 199436 156012 199442
rect 155960 199378 156012 199384
rect 148968 198008 149020 198014
rect 148968 197950 149020 197956
rect 146142 197390 146340 197418
rect 148980 197404 149008 197950
rect 155972 197470 156000 199378
rect 154488 197464 154540 197470
rect 154146 197412 154488 197418
rect 154146 197406 154540 197412
rect 155960 197464 156012 197470
rect 155960 197406 156012 197412
rect 154146 197390 154528 197406
rect 157996 197334 158024 228414
rect 152740 197328 152792 197334
rect 152582 197276 152740 197282
rect 152582 197270 152792 197276
rect 157984 197328 158036 197334
rect 157984 197270 158036 197276
rect 152582 197254 152780 197270
rect 167656 196790 167684 229706
rect 176660 227044 176712 227050
rect 176660 226986 176712 226992
rect 147956 196784 148008 196790
rect 147798 196732 147956 196738
rect 147798 196726 148008 196732
rect 167644 196784 167696 196790
rect 167644 196726 167696 196732
rect 147798 196710 147996 196726
rect 160836 196716 160888 196722
rect 160836 196658 160888 196664
rect 151176 196648 151228 196654
rect 150926 196596 151176 196602
rect 150926 196590 151228 196596
rect 150926 196574 151216 196590
rect 140424 196030 140530 196058
rect 157366 196030 157564 196058
rect 138664 195968 138716 195974
rect 138110 195936 138166 195945
rect 120000 195894 120120 195922
rect 116584 194540 116636 194546
rect 116584 194482 116636 194488
rect 120092 192506 120120 195894
rect 140424 195945 140452 196030
rect 157536 195974 157564 196030
rect 141424 195968 141476 195974
rect 138664 195910 138716 195916
rect 140410 195936 140466 195945
rect 138110 195871 138166 195880
rect 139400 195900 139452 195906
rect 138124 195838 138152 195871
rect 140410 195871 140466 195880
rect 141422 195936 141424 195945
rect 157524 195968 157576 195974
rect 141476 195936 141478 195945
rect 158916 195937 158944 196044
rect 160848 195945 160876 196658
rect 157524 195910 157576 195916
rect 158902 195928 158958 195937
rect 141422 195871 141478 195880
rect 157432 195900 157484 195906
rect 139400 195842 139452 195848
rect 158902 195863 158958 195872
rect 160834 195936 160890 195945
rect 160834 195871 160890 195880
rect 157432 195842 157484 195848
rect 138112 195832 138164 195838
rect 138112 195774 138164 195780
rect 139412 195537 139440 195842
rect 157154 195664 157210 195673
rect 157444 195650 157472 195842
rect 157210 195622 157472 195650
rect 157154 195599 157210 195608
rect 139398 195528 139454 195537
rect 139398 195463 139454 195472
rect 124864 194540 124916 194546
rect 124864 194482 124916 194488
rect 120080 192500 120132 192506
rect 120080 192442 120132 192448
rect 117320 180124 117372 180130
rect 117320 180066 117372 180072
rect 117332 134994 117360 180066
rect 120724 178696 120776 178702
rect 120724 178638 120776 178644
rect 120080 177336 120132 177342
rect 120080 177278 120132 177284
rect 120092 151814 120120 177278
rect 120092 151786 120488 151814
rect 119344 137964 119396 137970
rect 119344 137906 119396 137912
rect 117332 134966 117806 134994
rect 119356 134980 119384 137906
rect 120460 134994 120488 151786
rect 120736 137970 120764 178638
rect 122840 176112 122892 176118
rect 122840 176054 122892 176060
rect 121460 175976 121512 175982
rect 121460 175918 121512 175924
rect 121472 151814 121500 175918
rect 122852 151814 122880 176054
rect 124876 173874 124904 194482
rect 128360 192500 128412 192506
rect 128360 192442 128412 192448
rect 128372 189106 128400 192442
rect 140870 191856 140926 191865
rect 140870 191791 140926 191800
rect 140778 190904 140834 190913
rect 140778 190839 140834 190848
rect 128360 189100 128412 189106
rect 128360 189042 128412 189048
rect 130384 189100 130436 189106
rect 130384 189042 130436 189048
rect 130396 179450 130424 189042
rect 135260 184204 135312 184210
rect 135260 184146 135312 184152
rect 130384 179444 130436 179450
rect 130384 179386 130436 179392
rect 135168 179376 135220 179382
rect 135168 179318 135220 179324
rect 134708 177812 134760 177818
rect 134708 177754 134760 177760
rect 134720 176118 134748 177754
rect 134708 176112 134760 176118
rect 134708 176054 134760 176060
rect 125600 174548 125652 174554
rect 125600 174490 125652 174496
rect 124864 173868 124916 173874
rect 124864 173810 124916 173816
rect 121472 151786 122144 151814
rect 122852 151786 123616 151814
rect 120724 137964 120776 137970
rect 120724 137906 120776 137912
rect 122116 134994 122144 151786
rect 123588 134994 123616 151786
rect 120460 134966 120934 134994
rect 122116 134966 122498 134994
rect 123588 134966 124062 134994
rect 125612 134980 125640 174490
rect 134524 174480 134576 174486
rect 134524 174422 134576 174428
rect 129740 173936 129792 173942
rect 129740 173878 129792 173884
rect 128268 173868 128320 173874
rect 128268 173810 128320 173816
rect 126980 173256 127032 173262
rect 126980 173198 127032 173204
rect 126992 134994 127020 173198
rect 128280 164898 128308 173810
rect 128360 171148 128412 171154
rect 128360 171090 128412 171096
rect 128268 164892 128320 164898
rect 128268 164834 128320 164840
rect 127624 153196 127676 153202
rect 127624 153138 127676 153144
rect 126992 134966 127190 134994
rect 127636 134842 127664 153138
rect 128372 134994 128400 171090
rect 129752 151814 129780 173878
rect 133880 172168 133932 172174
rect 133880 172110 133932 172116
rect 131120 171896 131172 171902
rect 131120 171838 131172 171844
rect 129832 155916 129884 155922
rect 129832 155858 129884 155864
rect 129844 153270 129872 155858
rect 129832 153264 129884 153270
rect 129832 153206 129884 153212
rect 131132 151814 131160 171838
rect 132500 171556 132552 171562
rect 132500 171498 132552 171504
rect 132512 151814 132540 171498
rect 133892 151814 133920 172110
rect 134536 155922 134564 174422
rect 135180 173194 135208 179318
rect 135168 173188 135220 173194
rect 135168 173130 135220 173136
rect 134524 155916 134576 155922
rect 134524 155858 134576 155864
rect 135272 151814 135300 184146
rect 140792 182617 140820 190839
rect 140884 184249 140912 191791
rect 140962 191720 141018 191729
rect 140962 191655 141018 191664
rect 140976 184385 141004 191655
rect 144550 191040 144606 191049
rect 144302 190998 144550 191026
rect 144550 190975 144606 190984
rect 144458 190632 144514 190641
rect 144394 190590 144458 190618
rect 144458 190567 144514 190576
rect 145838 189816 145894 189825
rect 145894 189774 145958 189802
rect 145838 189751 145894 189760
rect 166106 189366 166212 189394
rect 159560 185910 159588 188428
rect 166184 187678 166212 189366
rect 166172 187672 166224 187678
rect 166172 187614 166224 187620
rect 159548 185904 159600 185910
rect 159548 185846 159600 185852
rect 159916 185564 159968 185570
rect 159916 185506 159968 185512
rect 140962 184376 141018 184385
rect 140962 184311 141018 184320
rect 142436 184272 142488 184278
rect 140870 184240 140926 184249
rect 142436 184214 142488 184220
rect 142448 184212 142476 184214
rect 140870 184175 140926 184184
rect 144734 183832 144790 183841
rect 144734 183767 144790 183776
rect 144642 183696 144698 183705
rect 144642 183631 144698 183640
rect 140778 182608 140834 182617
rect 140778 182543 140834 182552
rect 136376 182158 136758 182186
rect 136376 180130 136404 182158
rect 144656 181558 144684 183631
rect 144644 181552 144696 181558
rect 144644 181494 144696 181500
rect 144748 181150 144776 183767
rect 145196 181552 145248 181558
rect 145196 181494 145248 181500
rect 145208 181257 145236 181494
rect 145194 181248 145250 181257
rect 159928 181218 159956 185506
rect 145194 181183 145250 181192
rect 157248 181212 157300 181218
rect 157248 181154 157300 181160
rect 159916 181212 159968 181218
rect 159916 181154 159968 181160
rect 144736 181144 144788 181150
rect 144736 181086 144788 181092
rect 150900 181076 150952 181082
rect 150900 181018 150952 181024
rect 144642 180976 144698 180985
rect 136468 180934 136758 180962
rect 144578 180934 144642 180962
rect 136364 180124 136416 180130
rect 136364 180066 136416 180072
rect 136468 178702 136496 180934
rect 144642 180911 144698 180920
rect 150912 180130 150940 181018
rect 157260 180674 157288 181154
rect 157248 180668 157300 180674
rect 157248 180610 157300 180616
rect 150900 180124 150952 180130
rect 150900 180066 150952 180072
rect 153936 180124 153988 180130
rect 153936 180066 153988 180072
rect 157248 180124 157300 180130
rect 157248 180066 157300 180072
rect 136560 179982 136758 180010
rect 136456 178696 136508 178702
rect 136456 178638 136508 178644
rect 136364 178424 136416 178430
rect 136364 178366 136416 178372
rect 136376 175982 136404 178366
rect 136560 177970 136588 179982
rect 153948 179602 153976 180066
rect 153948 179586 154436 179602
rect 153948 179580 154448 179586
rect 153948 179574 154396 179580
rect 154396 179522 154448 179528
rect 149334 179480 149390 179489
rect 149334 179415 149390 179424
rect 148046 179344 148102 179353
rect 148046 179279 148102 179288
rect 142666 179072 142722 179081
rect 136744 178838 136772 179044
rect 142666 179007 142722 179016
rect 144090 178936 144146 178945
rect 144090 178871 144146 178880
rect 136732 178832 136784 178838
rect 136732 178774 136784 178780
rect 141606 178800 141662 178809
rect 141606 178735 141662 178744
rect 136468 177942 136588 177970
rect 136468 177342 136496 177942
rect 136744 177834 136772 177956
rect 136652 177818 136772 177834
rect 136640 177812 136772 177818
rect 136692 177806 136772 177812
rect 136640 177754 136692 177760
rect 136456 177336 136508 177342
rect 136456 177278 136508 177284
rect 136468 177126 136758 177154
rect 136364 175976 136416 175982
rect 136364 175918 136416 175924
rect 136468 174554 136496 177126
rect 136560 175902 136758 175930
rect 136456 174548 136508 174554
rect 136456 174490 136508 174496
rect 136560 173262 136588 175902
rect 140502 175672 140558 175681
rect 140502 175607 140558 175616
rect 136548 173256 136600 173262
rect 136548 173198 136600 173204
rect 136744 171154 136772 174964
rect 140516 174418 140544 175607
rect 141620 175370 141648 178735
rect 141608 175364 141660 175370
rect 141608 175306 141660 175312
rect 144104 174758 144132 178871
rect 148060 177274 148088 179279
rect 144460 177268 144512 177274
rect 144460 177210 144512 177216
rect 148048 177268 148100 177274
rect 148048 177210 148100 177216
rect 144092 174752 144144 174758
rect 144092 174694 144144 174700
rect 140504 174412 140556 174418
rect 140504 174354 140556 174360
rect 137376 173936 137428 173942
rect 137428 173884 137586 173890
rect 137376 173878 137586 173884
rect 137388 173862 137586 173878
rect 138676 171902 138704 173196
rect 138664 171896 138716 171902
rect 138664 171838 138716 171844
rect 139688 171562 139716 173196
rect 140792 172174 140820 173196
rect 142436 172780 142488 172786
rect 142436 172722 142488 172728
rect 140780 172168 140832 172174
rect 140780 172110 140832 172116
rect 139676 171556 139728 171562
rect 139676 171498 139728 171504
rect 136732 171148 136784 171154
rect 136732 171090 136784 171096
rect 140780 171148 140832 171154
rect 140780 171090 140832 171096
rect 137284 164892 137336 164898
rect 137284 164834 137336 164840
rect 137296 154562 137324 164834
rect 137284 154556 137336 154562
rect 137284 154498 137336 154504
rect 140688 154556 140740 154562
rect 140688 154498 140740 154504
rect 129752 151786 129872 151814
rect 131132 151786 131528 151814
rect 132512 151786 133000 151814
rect 133892 151786 134656 151814
rect 135272 151786 136128 151814
rect 129844 134994 129872 151786
rect 131500 134994 131528 151786
rect 132972 134994 133000 151786
rect 134628 134994 134656 151786
rect 136100 134994 136128 151786
rect 140700 148374 140728 154498
rect 140792 151814 140820 171090
rect 140792 151786 140912 151814
rect 140688 148368 140740 148374
rect 140688 148310 140740 148316
rect 139674 138000 139730 138009
rect 139674 137935 139730 137944
rect 138112 136740 138164 136746
rect 138112 136682 138164 136688
rect 128372 134966 128754 134994
rect 129844 134966 130318 134994
rect 131500 134966 131882 134994
rect 132972 134966 133446 134994
rect 134628 134966 135010 134994
rect 136100 134966 136574 134994
rect 138124 134980 138152 136682
rect 139688 134980 139716 137935
rect 140884 134994 140912 151786
rect 142448 137970 142476 172722
rect 142632 161474 142660 173196
rect 143448 172916 143500 172922
rect 143448 172858 143500 172864
rect 142540 161446 142660 161474
rect 142436 137964 142488 137970
rect 142436 137906 142488 137912
rect 142540 136746 142568 161446
rect 143460 142154 143488 172858
rect 143540 172848 143592 172854
rect 143540 172790 143592 172796
rect 143552 151814 143580 172790
rect 143552 151786 144040 151814
rect 143184 142126 143488 142154
rect 142528 136740 142580 136746
rect 142528 136682 142580 136688
rect 143184 134994 143212 142126
rect 140884 134966 141266 134994
rect 142830 134966 143212 134994
rect 144012 134994 144040 151786
rect 144472 137698 144500 177210
rect 149348 175409 149376 179415
rect 157260 178566 157288 180066
rect 158628 179648 158680 179654
rect 157798 179616 157854 179625
rect 157798 179551 157800 179560
rect 157852 179551 157854 179560
rect 158534 179616 158590 179625
rect 158590 179596 158628 179602
rect 158590 179590 158680 179596
rect 166540 179648 166592 179654
rect 166540 179590 166592 179596
rect 158590 179574 158668 179590
rect 158534 179551 158590 179560
rect 157800 179522 157852 179528
rect 154396 178560 154448 178566
rect 153948 178508 154396 178514
rect 153948 178502 154448 178508
rect 157248 178560 157300 178566
rect 157248 178502 157300 178508
rect 153948 178498 154436 178502
rect 153108 178492 153160 178498
rect 153108 178434 153160 178440
rect 153936 178492 154436 178498
rect 153988 178486 154436 178492
rect 153936 178434 153988 178440
rect 153120 176458 153148 178434
rect 157798 178120 157854 178129
rect 153948 178090 154436 178106
rect 153936 178084 154448 178090
rect 153988 178078 154396 178084
rect 153936 178026 153988 178032
rect 157798 178055 157800 178064
rect 154396 178026 154448 178032
rect 157852 178055 157854 178064
rect 158534 178120 158590 178129
rect 158628 178084 158680 178090
rect 158590 178064 158628 178072
rect 158534 178055 158628 178064
rect 158548 178044 158628 178055
rect 157800 178026 157852 178032
rect 158628 178026 158680 178032
rect 153108 176452 153160 176458
rect 153108 176394 153160 176400
rect 153108 175432 153160 175438
rect 149334 175400 149390 175409
rect 153108 175374 153160 175380
rect 154578 175400 154634 175409
rect 149334 175335 149390 175344
rect 153120 174894 153148 175374
rect 153936 175364 153988 175370
rect 154634 175358 154974 175386
rect 154578 175335 154634 175344
rect 153936 175306 153988 175312
rect 153948 175250 153976 175306
rect 154396 175296 154448 175302
rect 153948 175244 154396 175250
rect 153948 175238 154448 175244
rect 156512 175296 156564 175302
rect 156512 175238 156564 175244
rect 153948 175222 154436 175238
rect 153108 174888 153160 174894
rect 153108 174830 153160 174836
rect 145472 174752 145524 174758
rect 145472 174694 145524 174700
rect 145484 174486 145512 174694
rect 145472 174480 145524 174486
rect 145472 174422 145524 174428
rect 155500 174480 155552 174486
rect 155500 174422 155552 174428
rect 147494 174176 147550 174185
rect 147494 174111 147550 174120
rect 144932 171154 144960 173196
rect 145668 172922 145696 173196
rect 145656 172916 145708 172922
rect 145656 172858 145708 172864
rect 146484 172916 146536 172922
rect 146484 172858 146536 172864
rect 144920 171148 144972 171154
rect 144920 171090 144972 171096
rect 146496 151814 146524 172858
rect 146680 172854 146708 173196
rect 146668 172848 146720 172854
rect 146668 172790 146720 172796
rect 147508 159322 147536 174111
rect 155512 173942 155540 174422
rect 155500 173936 155552 173942
rect 155500 173878 155552 173884
rect 147600 172786 147628 173196
rect 148612 172922 148640 173196
rect 148600 172916 148652 172922
rect 148600 172858 148652 172864
rect 147588 172780 147640 172786
rect 147588 172722 147640 172728
rect 149624 161474 149652 173196
rect 150636 171134 150664 173196
rect 149532 161446 149652 161474
rect 150452 171106 150664 171134
rect 147496 159316 147548 159322
rect 147496 159258 147548 159264
rect 146496 151786 147168 151814
rect 145932 137964 145984 137970
rect 145932 137906 145984 137912
rect 144460 137692 144512 137698
rect 144460 137634 144512 137640
rect 144012 134966 144394 134994
rect 145944 134980 145972 137906
rect 147140 134994 147168 151786
rect 149532 142154 149560 161446
rect 149704 159316 149756 159322
rect 149704 159258 149756 159264
rect 149716 146266 149744 159258
rect 149704 146260 149756 146266
rect 149704 146202 149756 146208
rect 149440 142126 149560 142154
rect 149440 134994 149468 142126
rect 147140 134966 147522 134994
rect 149086 134966 149468 134994
rect 150452 134994 150480 171106
rect 151648 161474 151676 173196
rect 152660 161474 152688 173196
rect 150544 161446 151676 161474
rect 152476 161446 152688 161474
rect 153488 173182 153686 173210
rect 150544 137970 150572 161446
rect 150532 137964 150584 137970
rect 150532 137906 150584 137912
rect 152188 137964 152240 137970
rect 152188 137906 152240 137912
rect 150452 134966 150650 134994
rect 152200 134980 152228 137906
rect 152476 137222 152504 161446
rect 152648 146260 152700 146266
rect 152648 146202 152700 146208
rect 152660 143546 152688 146202
rect 152648 143540 152700 143546
rect 152648 143482 152700 143488
rect 152464 137216 152516 137222
rect 152464 137158 152516 137164
rect 153488 136746 153516 173182
rect 156524 172922 156552 175238
rect 162492 174548 162544 174554
rect 162492 174490 162544 174496
rect 159456 173052 159508 173058
rect 159456 172994 159508 173000
rect 156512 172916 156564 172922
rect 156512 172858 156564 172864
rect 158444 172916 158496 172922
rect 158444 172858 158496 172864
rect 154856 143540 154908 143546
rect 154856 143482 154908 143488
rect 154868 137766 154896 143482
rect 154856 137760 154908 137766
rect 154856 137702 154908 137708
rect 156880 137692 156932 137698
rect 156880 137634 156932 137640
rect 153752 137216 153804 137222
rect 153752 137158 153804 137164
rect 153476 136740 153528 136746
rect 153476 136682 153528 136688
rect 153764 134980 153792 137158
rect 155316 136740 155368 136746
rect 155316 136682 155368 136688
rect 155328 134980 155356 136682
rect 156892 134980 156920 137634
rect 158456 134980 158484 172858
rect 159468 151814 159496 172994
rect 162504 151814 162532 174490
rect 162860 172984 162912 172990
rect 162860 172926 162912 172932
rect 162872 169726 162900 172926
rect 162860 169720 162912 169726
rect 162860 169662 162912 169668
rect 159468 151786 159680 151814
rect 162504 151786 162808 151814
rect 159652 134994 159680 151786
rect 162124 148368 162176 148374
rect 162124 148310 162176 148316
rect 161570 138816 161626 138825
rect 161570 138751 161626 138760
rect 159652 134966 160034 134994
rect 161584 134980 161612 138751
rect 162136 136542 162164 148310
rect 162780 137034 162808 151786
rect 163516 137698 163544 175100
rect 163504 137692 163556 137698
rect 163504 137634 163556 137640
rect 162780 137006 162900 137034
rect 162124 136536 162176 136542
rect 162124 136478 162176 136484
rect 162872 134994 162900 137006
rect 163608 136814 163636 173196
rect 164528 173182 164634 173210
rect 164528 137970 164556 173182
rect 164976 169720 165028 169726
rect 164976 169662 165028 169668
rect 164988 166326 165016 169662
rect 164976 166320 165028 166326
rect 164976 166262 165028 166268
rect 166552 161474 166580 179590
rect 167644 166320 167696 166326
rect 167644 166262 167696 166268
rect 166460 161446 166580 161474
rect 164516 137964 164568 137970
rect 164516 137906 164568 137912
rect 164700 137760 164752 137766
rect 164700 137702 164752 137708
rect 163596 136808 163648 136814
rect 163596 136750 163648 136756
rect 162872 134966 163162 134994
rect 164712 134980 164740 137702
rect 166460 134994 166488 161446
rect 167656 160138 167684 166262
rect 175372 162920 175424 162926
rect 175372 162862 175424 162868
rect 167644 160132 167696 160138
rect 167644 160074 167696 160080
rect 169024 160132 169076 160138
rect 169024 160074 169076 160080
rect 169036 149734 169064 160074
rect 175384 151814 175412 162862
rect 175384 151786 175504 151814
rect 169024 149728 169076 149734
rect 169024 149670 169076 149676
rect 170128 149728 170180 149734
rect 170128 149670 170180 149676
rect 170140 147626 170168 149670
rect 170128 147620 170180 147626
rect 170128 147562 170180 147568
rect 172428 147620 172480 147626
rect 172428 147562 172480 147568
rect 172440 142154 172468 147562
rect 172440 142126 172560 142154
rect 172532 138446 172560 142126
rect 172520 138440 172572 138446
rect 172520 138382 172572 138388
rect 174360 138440 174412 138446
rect 174360 138382 174412 138388
rect 172520 137964 172572 137970
rect 172520 137906 172572 137912
rect 167826 137592 167882 137601
rect 167826 137527 167882 137536
rect 166290 134966 166488 134994
rect 167840 134980 167868 137527
rect 169390 137456 169446 137465
rect 169390 137391 169446 137400
rect 169404 134980 169432 137391
rect 170956 136808 171008 136814
rect 170956 136750 171008 136756
rect 170968 134980 170996 136750
rect 172532 134980 172560 137906
rect 174084 137692 174136 137698
rect 174084 137634 174136 137640
rect 174096 134980 174124 137634
rect 174372 136610 174400 138382
rect 174360 136604 174412 136610
rect 174360 136546 174412 136552
rect 127624 134836 127676 134842
rect 127624 134778 127676 134784
rect 175372 133952 175424 133958
rect 175372 133894 175424 133900
rect 175384 130121 175412 133894
rect 175476 132494 175504 151786
rect 176016 136604 176068 136610
rect 176016 136546 176068 136552
rect 175924 136536 175976 136542
rect 175924 136478 175976 136484
rect 175476 132466 175596 132494
rect 175462 132424 175518 132433
rect 175462 132359 175518 132368
rect 175370 130112 175426 130121
rect 175370 130047 175426 130056
rect 175476 122834 175504 132359
rect 175568 128353 175596 132466
rect 175554 128344 175610 128353
rect 175554 128279 175610 128288
rect 175292 122806 175504 122834
rect 116584 84244 116636 84250
rect 116584 84186 116636 84192
rect 115846 83260 115902 83269
rect 115846 83195 115902 83204
rect 115204 74316 115256 74322
rect 115204 74258 115256 74264
rect 116596 73914 116624 84186
rect 118608 75676 118660 75682
rect 118608 75618 118660 75624
rect 170680 75676 170732 75682
rect 170680 75618 170732 75624
rect 116584 73908 116636 73914
rect 116584 73850 116636 73856
rect 118620 73166 118648 75618
rect 170404 75268 170456 75274
rect 170404 75210 170456 75216
rect 118608 73160 118660 73166
rect 118608 73102 118660 73108
rect 120080 73160 120132 73166
rect 120080 73102 120132 73108
rect 120908 73160 120960 73166
rect 120908 73102 120960 73108
rect 116584 72412 116636 72418
rect 116584 72354 116636 72360
rect 114468 22772 114520 22778
rect 114468 22714 114520 22720
rect 106292 16546 106504 16574
rect 113192 16546 114048 16574
rect 102140 10940 102192 10946
rect 102140 10882 102192 10888
rect 95792 10872 95844 10878
rect 95792 10814 95844 10820
rect 92480 10804 92532 10810
rect 92480 10746 92532 10752
rect 89166 10432 89222 10441
rect 89166 10367 89222 10376
rect 87970 7712 88026 7721
rect 87970 7647 88026 7656
rect 86224 6656 86276 6662
rect 86224 6598 86276 6604
rect 85672 5364 85724 5370
rect 85672 5306 85724 5312
rect 85684 480 85712 5306
rect 86868 5296 86920 5302
rect 86868 5238 86920 5244
rect 86880 480 86908 5238
rect 87984 480 88012 7647
rect 89180 480 89208 10367
rect 91558 7848 91614 7857
rect 91558 7783 91614 7792
rect 90362 4992 90418 5001
rect 90362 4927 90418 4936
rect 90376 480 90404 4927
rect 91572 480 91600 7783
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92492 354 92520 10746
rect 95148 8220 95200 8226
rect 95148 8162 95200 8168
rect 93952 5432 94004 5438
rect 93952 5374 94004 5380
rect 93964 480 93992 5374
rect 95160 480 95188 8162
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 95804 354 95832 10814
rect 98644 8288 98696 8294
rect 98644 8230 98696 8236
rect 97448 5500 97500 5506
rect 97448 5442 97500 5448
rect 97460 480 97488 5442
rect 98656 480 98684 8230
rect 99840 6792 99892 6798
rect 99840 6734 99892 6740
rect 99852 480 99880 6734
rect 101036 4140 101088 4146
rect 101036 4082 101088 4088
rect 101048 480 101076 4082
rect 102152 3398 102180 10882
rect 105726 9344 105782 9353
rect 105726 9279 105782 9288
rect 102232 7540 102284 7546
rect 102232 7482 102284 7488
rect 102140 3392 102192 3398
rect 102140 3334 102192 3340
rect 102244 480 102272 7482
rect 104532 6656 104584 6662
rect 104532 6598 104584 6604
rect 103336 3392 103388 3398
rect 103336 3334 103388 3340
rect 103348 480 103376 3334
rect 104544 480 104572 6598
rect 105740 480 105768 9279
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 110512 11008 110564 11014
rect 110512 10950 110564 10956
rect 109314 9480 109370 9489
rect 109314 9415 109370 9424
rect 108118 6624 108174 6633
rect 108118 6559 108174 6568
rect 108132 480 108160 6559
rect 109328 480 109356 9415
rect 110524 480 110552 10950
rect 112812 9580 112864 9586
rect 112812 9522 112864 9528
rect 111616 4752 111668 4758
rect 111616 4694 111668 4700
rect 111628 480 111656 4694
rect 112824 480 112852 9522
rect 114020 480 114048 16546
rect 116400 9648 116452 9654
rect 116400 9590 116452 9596
rect 115204 6860 115256 6866
rect 115204 6802 115256 6808
rect 115216 480 115244 6802
rect 116412 480 116440 9590
rect 116596 9382 116624 72354
rect 118148 72344 118200 72350
rect 118148 72286 118200 72292
rect 117964 72208 118016 72214
rect 117964 72150 118016 72156
rect 117320 10260 117372 10266
rect 117320 10202 117372 10208
rect 116584 9376 116636 9382
rect 116584 9318 116636 9324
rect 117228 4684 117280 4690
rect 117228 4626 117280 4632
rect 117240 4146 117268 4626
rect 117228 4140 117280 4146
rect 117228 4082 117280 4088
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117332 354 117360 10202
rect 117976 4962 118004 72150
rect 118056 72140 118108 72146
rect 118056 72082 118108 72088
rect 118068 7682 118096 72082
rect 118160 18630 118188 72286
rect 119344 71868 119396 71874
rect 119344 71810 119396 71816
rect 119356 54534 119384 71810
rect 120092 71398 120120 73102
rect 120724 73024 120776 73030
rect 120724 72966 120776 72972
rect 120080 71392 120132 71398
rect 120080 71334 120132 71340
rect 119344 54528 119396 54534
rect 119344 54470 119396 54476
rect 118148 18624 118200 18630
rect 118148 18566 118200 18572
rect 120632 10192 120684 10198
rect 120632 10134 120684 10140
rect 118056 7676 118108 7682
rect 118056 7618 118108 7624
rect 119896 7676 119948 7682
rect 119896 7618 119948 7624
rect 117964 4956 118016 4962
rect 117964 4898 118016 4904
rect 118792 4956 118844 4962
rect 118792 4898 118844 4904
rect 118804 480 118832 4898
rect 119908 480 119936 7618
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 10134
rect 120736 5370 120764 72966
rect 120816 72956 120868 72962
rect 120816 72898 120868 72904
rect 120828 6798 120856 72898
rect 120920 25566 120948 73102
rect 121092 72888 121144 72894
rect 121092 72830 121144 72836
rect 121000 72752 121052 72758
rect 121000 72694 121052 72700
rect 121012 43450 121040 72694
rect 121104 51134 121132 72830
rect 121368 72684 121420 72690
rect 121368 72626 121420 72632
rect 121092 51128 121144 51134
rect 121092 51070 121144 51076
rect 121000 43444 121052 43450
rect 121000 43386 121052 43392
rect 120908 25560 120960 25566
rect 120908 25502 120960 25508
rect 120816 6792 120868 6798
rect 120816 6734 120868 6740
rect 120724 5364 120776 5370
rect 120724 5306 120776 5312
rect 121380 4146 121408 72626
rect 121564 71913 121592 75140
rect 121656 72049 121684 75140
rect 121642 72040 121698 72049
rect 121642 71975 121698 71984
rect 121550 71904 121606 71913
rect 121550 71839 121606 71848
rect 121552 70032 121604 70038
rect 121748 69986 121776 75140
rect 121552 69974 121604 69980
rect 121460 69896 121512 69902
rect 121460 69838 121512 69844
rect 121472 66910 121500 69838
rect 121460 66904 121512 66910
rect 121460 66846 121512 66852
rect 121564 64874 121592 69974
rect 121656 69958 121776 69986
rect 121656 68270 121684 69958
rect 121736 69828 121788 69834
rect 121736 69770 121788 69776
rect 121748 69578 121776 69770
rect 121840 69714 121868 75140
rect 121932 72593 121960 75140
rect 121918 72584 121974 72593
rect 121918 72519 121974 72528
rect 122024 69902 122052 75140
rect 122116 69902 122144 75140
rect 122012 69896 122064 69902
rect 122012 69838 122064 69844
rect 122104 69896 122156 69902
rect 122104 69838 122156 69844
rect 122208 69834 122236 75140
rect 122196 69828 122248 69834
rect 122196 69770 122248 69776
rect 122300 69714 122328 75140
rect 122392 72282 122420 75140
rect 122380 72276 122432 72282
rect 122380 72218 122432 72224
rect 122380 71800 122432 71806
rect 122380 71742 122432 71748
rect 121840 69686 121960 69714
rect 121748 69550 121868 69578
rect 121644 68264 121696 68270
rect 121644 68206 121696 68212
rect 121564 64846 121776 64874
rect 121748 6322 121776 64846
rect 121736 6316 121788 6322
rect 121736 6258 121788 6264
rect 121840 6254 121868 69550
rect 121828 6248 121880 6254
rect 121828 6190 121880 6196
rect 121932 6186 121960 69686
rect 122024 69686 122328 69714
rect 122024 8974 122052 69686
rect 122104 69624 122156 69630
rect 122104 69566 122156 69572
rect 122116 13122 122144 69566
rect 122392 68354 122420 71742
rect 122208 68326 122420 68354
rect 122104 13116 122156 13122
rect 122104 13058 122156 13064
rect 122208 10742 122236 68326
rect 122288 68264 122340 68270
rect 122288 68206 122340 68212
rect 122196 10736 122248 10742
rect 122196 10678 122248 10684
rect 122012 8968 122064 8974
rect 122012 8910 122064 8916
rect 122300 6914 122328 68206
rect 122208 6886 122328 6914
rect 121920 6180 121972 6186
rect 121920 6122 121972 6128
rect 121368 4140 121420 4146
rect 121368 4082 121420 4088
rect 122208 3466 122236 6886
rect 122484 3602 122512 75140
rect 122576 70038 122604 75140
rect 122564 70032 122616 70038
rect 122564 69974 122616 69980
rect 122564 69896 122616 69902
rect 122564 69838 122616 69844
rect 122472 3596 122524 3602
rect 122472 3538 122524 3544
rect 122576 3534 122604 69838
rect 122668 69630 122696 75140
rect 122760 71874 122788 75140
rect 122852 72049 122880 75140
rect 122838 72040 122894 72049
rect 122838 71975 122894 71984
rect 122944 71913 122972 75140
rect 123036 72146 123064 75140
rect 123128 72486 123156 75140
rect 123116 72480 123168 72486
rect 123116 72422 123168 72428
rect 123024 72140 123076 72146
rect 123024 72082 123076 72088
rect 122930 71904 122986 71913
rect 122748 71868 122800 71874
rect 122930 71839 122986 71848
rect 122748 71810 122800 71816
rect 123220 70122 123248 75140
rect 122932 70100 122984 70106
rect 122932 70042 122984 70048
rect 123128 70094 123248 70122
rect 122656 69624 122708 69630
rect 122656 69566 122708 69572
rect 122944 64874 122972 70042
rect 123024 70032 123076 70038
rect 123024 69974 123076 69980
rect 123036 69442 123064 69974
rect 123128 69562 123156 70094
rect 123208 69964 123260 69970
rect 123208 69906 123260 69912
rect 123116 69556 123168 69562
rect 123116 69498 123168 69504
rect 123036 69414 123156 69442
rect 122944 64846 123064 64874
rect 123036 5030 123064 64846
rect 123128 6390 123156 69414
rect 123220 7750 123248 69906
rect 123208 7744 123260 7750
rect 123208 7686 123260 7692
rect 123312 7614 123340 75140
rect 123404 9042 123432 75140
rect 123496 69714 123524 75140
rect 123588 69902 123616 75140
rect 123680 69970 123708 75140
rect 123772 72214 123800 75140
rect 123760 72208 123812 72214
rect 123760 72150 123812 72156
rect 123864 70038 123892 75140
rect 123852 70032 123904 70038
rect 123852 69974 123904 69980
rect 123668 69964 123720 69970
rect 123668 69906 123720 69912
rect 123576 69896 123628 69902
rect 123576 69838 123628 69844
rect 123956 69834 123984 75140
rect 123944 69828 123996 69834
rect 123944 69770 123996 69776
rect 124048 69714 124076 75140
rect 124140 70106 124168 75140
rect 124232 72185 124260 75140
rect 124324 72350 124352 75140
rect 124312 72344 124364 72350
rect 124312 72286 124364 72292
rect 124218 72176 124274 72185
rect 124218 72111 124274 72120
rect 124416 72049 124444 75140
rect 124402 72040 124458 72049
rect 124402 71975 124458 71984
rect 124508 71913 124536 75140
rect 124494 71904 124550 71913
rect 124494 71839 124550 71848
rect 124128 70100 124180 70106
rect 124128 70042 124180 70048
rect 124312 70032 124364 70038
rect 124312 69974 124364 69980
rect 124128 69896 124180 69902
rect 124128 69838 124180 69844
rect 123496 69686 123616 69714
rect 123484 69624 123536 69630
rect 123484 69566 123536 69572
rect 123496 9110 123524 69566
rect 123588 10334 123616 69686
rect 123680 69686 124076 69714
rect 123680 10402 123708 69686
rect 123760 69556 123812 69562
rect 123760 69498 123812 69504
rect 123668 10396 123720 10402
rect 123668 10338 123720 10344
rect 123576 10328 123628 10334
rect 123576 10270 123628 10276
rect 123484 9104 123536 9110
rect 123484 9046 123536 9052
rect 123392 9036 123444 9042
rect 123392 8978 123444 8984
rect 123300 7608 123352 7614
rect 123300 7550 123352 7556
rect 123116 6384 123168 6390
rect 123116 6326 123168 6332
rect 123024 5024 123076 5030
rect 123024 4966 123076 4972
rect 123772 4826 123800 69498
rect 124140 4894 124168 69838
rect 124128 4888 124180 4894
rect 124128 4830 124180 4836
rect 123760 4820 123812 4826
rect 123760 4762 123812 4768
rect 124324 3738 124352 69974
rect 124600 69902 124628 75140
rect 124588 69896 124640 69902
rect 124588 69838 124640 69844
rect 124496 69828 124548 69834
rect 124496 69770 124548 69776
rect 124508 6526 124536 69770
rect 124692 69714 124720 75140
rect 124600 69686 124720 69714
rect 124496 6520 124548 6526
rect 124496 6462 124548 6468
rect 124600 6458 124628 69686
rect 124784 69578 124812 75140
rect 124876 72418 124904 75140
rect 124864 72412 124916 72418
rect 124864 72354 124916 72360
rect 124968 69834 124996 75140
rect 124956 69828 125008 69834
rect 124956 69770 125008 69776
rect 124784 69550 124996 69578
rect 124864 69488 124916 69494
rect 124864 69430 124916 69436
rect 124680 67380 124732 67386
rect 124680 67322 124732 67328
rect 124692 6594 124720 67322
rect 124772 65952 124824 65958
rect 124772 65894 124824 65900
rect 124784 9246 124812 65894
rect 124876 9314 124904 69430
rect 124864 9308 124916 9314
rect 124864 9250 124916 9256
rect 124772 9240 124824 9246
rect 124772 9182 124824 9188
rect 124968 9178 124996 69550
rect 125060 65958 125088 75140
rect 125048 65952 125100 65958
rect 125048 65894 125100 65900
rect 125152 64874 125180 75140
rect 125244 70038 125272 75140
rect 125232 70032 125284 70038
rect 125232 69974 125284 69980
rect 125232 69896 125284 69902
rect 125232 69838 125284 69844
rect 125060 64846 125180 64874
rect 125060 10470 125088 64846
rect 125048 10464 125100 10470
rect 125048 10406 125100 10412
rect 124956 9172 125008 9178
rect 124956 9114 125008 9120
rect 124680 6588 124732 6594
rect 124680 6530 124732 6536
rect 124588 6452 124640 6458
rect 124588 6394 124640 6400
rect 124312 3732 124364 3738
rect 124312 3674 124364 3680
rect 125244 3670 125272 69838
rect 125336 67386 125364 75140
rect 125428 69494 125456 75140
rect 125416 69488 125468 69494
rect 125416 69430 125468 69436
rect 125324 67380 125376 67386
rect 125324 67322 125376 67328
rect 125520 3806 125548 75140
rect 125612 72185 125640 75140
rect 125704 72321 125732 75140
rect 125690 72312 125746 72321
rect 125690 72247 125746 72256
rect 125598 72176 125654 72185
rect 125598 72111 125654 72120
rect 125796 72049 125824 75140
rect 125782 72040 125838 72049
rect 125782 71975 125838 71984
rect 125888 71913 125916 75140
rect 125874 71904 125930 71913
rect 125874 71839 125930 71848
rect 125692 69760 125744 69766
rect 125692 69702 125744 69708
rect 125704 64874 125732 69702
rect 125784 69692 125836 69698
rect 125784 69634 125836 69640
rect 125796 67590 125824 69634
rect 125980 67862 126008 75140
rect 126072 69222 126100 75140
rect 126060 69216 126112 69222
rect 126060 69158 126112 69164
rect 126164 68082 126192 75140
rect 126072 68054 126192 68082
rect 125968 67856 126020 67862
rect 125968 67798 126020 67804
rect 126072 67674 126100 68054
rect 126256 67946 126284 75140
rect 126348 72554 126376 75140
rect 126336 72548 126388 72554
rect 126336 72490 126388 72496
rect 126440 69698 126468 75140
rect 126428 69692 126480 69698
rect 126428 69634 126480 69640
rect 126532 69442 126560 75140
rect 126624 69766 126652 75140
rect 126612 69760 126664 69766
rect 126612 69702 126664 69708
rect 125888 67646 126100 67674
rect 126164 67918 126284 67946
rect 126348 69414 126560 69442
rect 125784 67584 125836 67590
rect 125784 67526 125836 67532
rect 125704 64846 125824 64874
rect 125796 5098 125824 64846
rect 125888 6730 125916 67646
rect 125968 67584 126020 67590
rect 125968 67526 126020 67532
rect 126060 67584 126112 67590
rect 126060 67526 126112 67532
rect 125980 7818 126008 67526
rect 126072 7886 126100 67526
rect 126164 9518 126192 67918
rect 126244 67856 126296 67862
rect 126244 67798 126296 67804
rect 126152 9512 126204 9518
rect 126152 9454 126204 9460
rect 126256 9450 126284 67798
rect 126348 10538 126376 69414
rect 126428 69352 126480 69358
rect 126428 69294 126480 69300
rect 126440 10606 126468 69294
rect 126520 69216 126572 69222
rect 126520 69158 126572 69164
rect 126428 10600 126480 10606
rect 126428 10542 126480 10548
rect 126336 10532 126388 10538
rect 126336 10474 126388 10480
rect 126244 9444 126296 9450
rect 126244 9386 126296 9392
rect 126060 7880 126112 7886
rect 126060 7822 126112 7828
rect 125968 7812 126020 7818
rect 125968 7754 126020 7760
rect 125876 6724 125928 6730
rect 125876 6666 125928 6672
rect 125784 5092 125836 5098
rect 125784 5034 125836 5040
rect 126532 3874 126560 69158
rect 126716 67590 126744 75140
rect 126808 69358 126836 75140
rect 126796 69352 126848 69358
rect 126796 69294 126848 69300
rect 126704 67584 126756 67590
rect 126704 67526 126756 67532
rect 126900 3942 126928 75140
rect 126992 71913 127020 75140
rect 127084 72049 127112 75140
rect 127070 72040 127126 72049
rect 127070 71975 127126 71984
rect 126978 71904 127034 71913
rect 126978 71839 127034 71848
rect 127072 69828 127124 69834
rect 127072 69770 127124 69776
rect 127084 4010 127112 69770
rect 127176 69714 127204 75140
rect 127268 69850 127296 75140
rect 127360 71806 127388 75140
rect 127348 71800 127400 71806
rect 127348 71742 127400 71748
rect 127268 69822 127388 69850
rect 127176 69686 127296 69714
rect 127164 69624 127216 69630
rect 127164 69566 127216 69572
rect 127176 5234 127204 69566
rect 127164 5228 127216 5234
rect 127164 5170 127216 5176
rect 127268 5166 127296 69686
rect 127360 69562 127388 69822
rect 127452 69630 127480 75140
rect 127440 69624 127492 69630
rect 127440 69566 127492 69572
rect 127348 69556 127400 69562
rect 127348 69498 127400 69504
rect 127440 69352 127492 69358
rect 127440 69294 127492 69300
rect 127348 69284 127400 69290
rect 127348 69226 127400 69232
rect 127360 5302 127388 69226
rect 127452 8090 127480 69294
rect 127440 8084 127492 8090
rect 127440 8026 127492 8032
rect 127544 8022 127572 75140
rect 127636 69714 127664 75140
rect 127728 69834 127756 75140
rect 127820 69850 127848 75140
rect 127912 73166 127940 75140
rect 127900 73160 127952 73166
rect 127900 73102 127952 73108
rect 127716 69828 127768 69834
rect 127820 69822 127940 69850
rect 127716 69770 127768 69776
rect 127636 69686 127848 69714
rect 127624 69556 127676 69562
rect 127624 69498 127676 69504
rect 127532 8016 127584 8022
rect 127532 7958 127584 7964
rect 127636 7954 127664 69498
rect 127716 69148 127768 69154
rect 127716 69090 127768 69096
rect 127728 8158 127756 69090
rect 127820 10674 127848 69686
rect 127912 69358 127940 69822
rect 127900 69352 127952 69358
rect 127900 69294 127952 69300
rect 127808 10668 127860 10674
rect 127808 10610 127860 10616
rect 127716 8152 127768 8158
rect 127716 8094 127768 8100
rect 127624 7948 127676 7954
rect 127624 7890 127676 7896
rect 127348 5296 127400 5302
rect 127348 5238 127400 5244
rect 127256 5160 127308 5166
rect 127256 5102 127308 5108
rect 128004 4078 128032 75140
rect 128096 69154 128124 75140
rect 128188 73030 128216 75140
rect 128176 73024 128228 73030
rect 128176 72966 128228 72972
rect 128280 69290 128308 75140
rect 128372 72049 128400 75140
rect 128464 72185 128492 75140
rect 128556 73137 128584 75140
rect 128542 73128 128598 73137
rect 128542 73063 128598 73072
rect 128450 72176 128506 72185
rect 128450 72111 128506 72120
rect 128358 72040 128414 72049
rect 128358 71975 128414 71984
rect 128648 71913 128676 75140
rect 128634 71904 128690 71913
rect 128634 71839 128690 71848
rect 128544 70032 128596 70038
rect 128544 69974 128596 69980
rect 128268 69284 128320 69290
rect 128268 69226 128320 69232
rect 128084 69148 128136 69154
rect 128084 69090 128136 69096
rect 128556 4690 128584 69974
rect 128740 69714 128768 75140
rect 128648 69686 128768 69714
rect 128648 65482 128676 69686
rect 128832 69630 128860 75140
rect 128820 69624 128872 69630
rect 128820 69566 128872 69572
rect 128924 65770 128952 75140
rect 128740 65742 128952 65770
rect 128636 65476 128688 65482
rect 128636 65418 128688 65424
rect 128636 65340 128688 65346
rect 128636 65282 128688 65288
rect 128648 6662 128676 65282
rect 128740 8226 128768 65742
rect 128820 65680 128872 65686
rect 128820 65622 128872 65628
rect 128728 8220 128780 8226
rect 128728 8162 128780 8168
rect 128832 7546 128860 65622
rect 128912 65612 128964 65618
rect 128912 65554 128964 65560
rect 128924 8294 128952 65554
rect 129016 10878 129044 75140
rect 129108 69850 129136 75140
rect 129200 69970 129228 75140
rect 129292 72962 129320 75140
rect 129280 72956 129332 72962
rect 129280 72898 129332 72904
rect 129384 70038 129412 75140
rect 129372 70032 129424 70038
rect 129372 69974 129424 69980
rect 129188 69964 129240 69970
rect 129188 69906 129240 69912
rect 129108 69822 129320 69850
rect 129292 69714 129320 69822
rect 129188 69692 129240 69698
rect 129292 69686 129412 69714
rect 129188 69634 129240 69640
rect 129200 65618 129228 69634
rect 129280 69624 129332 69630
rect 129280 69566 129332 69572
rect 129188 65612 129240 65618
rect 129188 65554 129240 65560
rect 129096 65544 129148 65550
rect 129096 65486 129148 65492
rect 129108 10946 129136 65486
rect 129188 65476 129240 65482
rect 129188 65418 129240 65424
rect 129096 10940 129148 10946
rect 129096 10882 129148 10888
rect 129004 10872 129056 10878
rect 129004 10814 129056 10820
rect 129200 10810 129228 65418
rect 129188 10804 129240 10810
rect 129188 10746 129240 10752
rect 128912 8288 128964 8294
rect 128912 8230 128964 8236
rect 128820 7540 128872 7546
rect 128820 7482 128872 7488
rect 128636 6656 128688 6662
rect 128636 6598 128688 6604
rect 129292 5438 129320 69566
rect 129384 5506 129412 69686
rect 129476 65686 129504 75140
rect 129464 65680 129516 65686
rect 129464 65622 129516 65628
rect 129568 65550 129596 75140
rect 129556 65544 129608 65550
rect 129556 65486 129608 65492
rect 129660 65346 129688 75140
rect 129752 72185 129780 75140
rect 129844 72758 129872 75140
rect 129832 72752 129884 72758
rect 129832 72694 129884 72700
rect 129738 72176 129794 72185
rect 129738 72111 129794 72120
rect 129936 71913 129964 75140
rect 130028 72049 130056 75140
rect 130014 72040 130070 72049
rect 130014 71975 130070 71984
rect 129922 71904 129978 71913
rect 129922 71839 129978 71848
rect 130120 69970 130148 75140
rect 130108 69964 130160 69970
rect 130108 69906 130160 69912
rect 130212 69850 130240 75140
rect 129844 69822 130240 69850
rect 129648 65340 129700 65346
rect 129648 65282 129700 65288
rect 129372 5500 129424 5506
rect 129372 5442 129424 5448
rect 129280 5432 129332 5438
rect 129280 5374 129332 5380
rect 129844 4758 129872 69822
rect 130016 69760 130068 69766
rect 130016 69702 130068 69708
rect 129924 67652 129976 67658
rect 129924 67594 129976 67600
rect 129936 4962 129964 67594
rect 130028 6866 130056 69702
rect 130200 69624 130252 69630
rect 130200 69566 130252 69572
rect 130108 69556 130160 69562
rect 130108 69498 130160 69504
rect 130120 7682 130148 69498
rect 130212 9654 130240 69566
rect 130200 9648 130252 9654
rect 130200 9590 130252 9596
rect 130304 9586 130332 75140
rect 130396 72894 130424 75140
rect 130384 72888 130436 72894
rect 130384 72830 130436 72836
rect 130384 69964 130436 69970
rect 130384 69906 130436 69912
rect 130396 11014 130424 69906
rect 130488 69834 130516 75140
rect 130476 69828 130528 69834
rect 130476 69770 130528 69776
rect 130476 69692 130528 69698
rect 130476 69634 130528 69640
rect 130384 11008 130436 11014
rect 130384 10950 130436 10956
rect 130488 10198 130516 69634
rect 130580 69630 130608 75140
rect 130568 69624 130620 69630
rect 130568 69566 130620 69572
rect 130672 64874 130700 75140
rect 130764 67658 130792 75140
rect 130856 69562 130884 75140
rect 130948 69698 130976 75140
rect 130936 69692 130988 69698
rect 130936 69634 130988 69640
rect 130844 69556 130896 69562
rect 130844 69498 130896 69504
rect 130752 67652 130804 67658
rect 130752 67594 130804 67600
rect 130580 64846 130700 64874
rect 130580 10266 130608 64846
rect 130568 10260 130620 10266
rect 130568 10202 130620 10208
rect 130476 10192 130528 10198
rect 130476 10134 130528 10140
rect 130292 9580 130344 9586
rect 130292 9522 130344 9528
rect 130108 7676 130160 7682
rect 130108 7618 130160 7624
rect 130016 6860 130068 6866
rect 130016 6802 130068 6808
rect 129924 4956 129976 4962
rect 129924 4898 129976 4904
rect 129832 4752 129884 4758
rect 129832 4694 129884 4700
rect 128544 4684 128596 4690
rect 128544 4626 128596 4632
rect 127992 4072 128044 4078
rect 127992 4014 128044 4020
rect 127072 4004 127124 4010
rect 127072 3946 127124 3952
rect 126888 3936 126940 3942
rect 126888 3878 126940 3884
rect 126520 3868 126572 3874
rect 126520 3810 126572 3816
rect 125508 3800 125560 3806
rect 125508 3742 125560 3748
rect 125232 3664 125284 3670
rect 123482 3632 123538 3641
rect 125232 3606 125284 3612
rect 123482 3567 123538 3576
rect 125876 3596 125928 3602
rect 122564 3528 122616 3534
rect 122564 3470 122616 3476
rect 122196 3460 122248 3466
rect 122196 3402 122248 3408
rect 122288 3392 122340 3398
rect 122288 3334 122340 3340
rect 122300 480 122328 3334
rect 123496 480 123524 3567
rect 125876 3538 125928 3544
rect 124678 3496 124734 3505
rect 124678 3431 124734 3440
rect 124692 480 124720 3431
rect 125888 480 125916 3538
rect 129372 3528 129424 3534
rect 129372 3470 129424 3476
rect 126980 3460 127032 3466
rect 126980 3402 127032 3408
rect 126992 480 127020 3402
rect 128176 3188 128228 3194
rect 128176 3130 128228 3136
rect 128188 480 128216 3130
rect 129384 480 129412 3470
rect 131040 3398 131068 75140
rect 131132 71913 131160 75140
rect 131224 72049 131252 75140
rect 131210 72040 131266 72049
rect 131210 71975 131266 71984
rect 131118 71904 131174 71913
rect 131118 71839 131174 71848
rect 131212 70100 131264 70106
rect 131212 70042 131264 70048
rect 131120 69692 131172 69698
rect 131120 69634 131172 69640
rect 131132 11694 131160 69634
rect 131120 11688 131172 11694
rect 131120 11630 131172 11636
rect 131120 11552 131172 11558
rect 131120 11494 131172 11500
rect 131132 3602 131160 11494
rect 131120 3596 131172 3602
rect 131120 3538 131172 3544
rect 131224 3534 131252 70042
rect 131316 69562 131344 75140
rect 131408 69714 131436 75140
rect 131500 69986 131528 75140
rect 131592 70106 131620 75140
rect 131580 70100 131632 70106
rect 131580 70042 131632 70048
rect 131500 69958 131620 69986
rect 131408 69686 131528 69714
rect 131304 69556 131356 69562
rect 131304 69498 131356 69504
rect 131500 69442 131528 69686
rect 131316 69414 131528 69442
rect 131592 69426 131620 69958
rect 131580 69420 131632 69426
rect 131316 11778 131344 69414
rect 131580 69362 131632 69368
rect 131396 69352 131448 69358
rect 131684 69306 131712 75140
rect 131776 69698 131804 75140
rect 131764 69692 131816 69698
rect 131764 69634 131816 69640
rect 131396 69294 131448 69300
rect 131408 11898 131436 69294
rect 131500 69278 131712 69306
rect 131396 11892 131448 11898
rect 131396 11834 131448 11840
rect 131316 11750 131436 11778
rect 131304 11688 131356 11694
rect 131304 11630 131356 11636
rect 131212 3528 131264 3534
rect 131212 3470 131264 3476
rect 131028 3392 131080 3398
rect 131028 3334 131080 3340
rect 130568 3324 130620 3330
rect 130568 3266 130620 3272
rect 130580 480 130608 3266
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131316 354 131344 11630
rect 131408 3466 131436 11750
rect 131396 3460 131448 3466
rect 131396 3402 131448 3408
rect 131500 3330 131528 69278
rect 131580 69216 131632 69222
rect 131580 69158 131632 69164
rect 131488 3324 131540 3330
rect 131488 3266 131540 3272
rect 131592 3194 131620 69158
rect 131868 4078 131896 75140
rect 131856 4072 131908 4078
rect 131856 4014 131908 4020
rect 131960 3398 131988 75140
rect 132052 3942 132080 75140
rect 132040 3936 132092 3942
rect 132040 3878 132092 3884
rect 131948 3392 132000 3398
rect 131948 3334 132000 3340
rect 132144 3330 132172 75140
rect 132236 72049 132264 75140
rect 132328 72622 132356 75140
rect 132316 72616 132368 72622
rect 132316 72558 132368 72564
rect 132222 72040 132278 72049
rect 132222 71975 132278 71984
rect 132420 71913 132448 75140
rect 132406 71904 132462 71913
rect 132512 71874 132540 75140
rect 132406 71839 132462 71848
rect 132500 71868 132552 71874
rect 132500 71810 132552 71816
rect 132604 5438 132632 75140
rect 132696 72690 132724 75140
rect 132684 72684 132736 72690
rect 132684 72626 132736 72632
rect 132592 5432 132644 5438
rect 132592 5374 132644 5380
rect 132788 5370 132816 75140
rect 132776 5364 132828 5370
rect 132776 5306 132828 5312
rect 132880 4010 132908 75140
rect 132972 4978 133000 75140
rect 133064 5166 133092 75140
rect 133052 5160 133104 5166
rect 133052 5102 133104 5108
rect 133156 5098 133184 75140
rect 133144 5092 133196 5098
rect 133144 5034 133196 5040
rect 132972 4950 133092 4978
rect 132960 4072 133012 4078
rect 132960 4014 133012 4020
rect 132868 4004 132920 4010
rect 132868 3946 132920 3952
rect 132132 3324 132184 3330
rect 132132 3266 132184 3272
rect 131580 3188 131632 3194
rect 131580 3130 131632 3136
rect 132972 480 133000 4014
rect 133064 3602 133092 4950
rect 133052 3596 133104 3602
rect 133052 3538 133104 3544
rect 133248 3534 133276 75140
rect 133340 4962 133368 75140
rect 133432 5030 133460 75140
rect 133420 5024 133472 5030
rect 133420 4966 133472 4972
rect 133328 4956 133380 4962
rect 133328 4898 133380 4904
rect 133236 3528 133288 3534
rect 133236 3470 133288 3476
rect 133524 3466 133552 75140
rect 133616 72049 133644 75140
rect 133708 72185 133736 75140
rect 133694 72176 133750 72185
rect 133694 72111 133750 72120
rect 133602 72040 133658 72049
rect 133602 71975 133658 71984
rect 133800 71913 133828 75140
rect 133786 71904 133842 71913
rect 133786 71839 133842 71848
rect 133892 4894 133920 75140
rect 133984 71806 134012 75140
rect 133972 71800 134024 71806
rect 133972 71742 134024 71748
rect 133880 4888 133932 4894
rect 133880 4830 133932 4836
rect 134076 4010 134104 75140
rect 134064 4004 134116 4010
rect 134064 3946 134116 3952
rect 134168 3874 134196 75140
rect 134260 4826 134288 75140
rect 134248 4820 134300 4826
rect 134248 4762 134300 4768
rect 134156 3868 134208 3874
rect 134156 3810 134208 3816
rect 134352 3806 134380 75140
rect 134340 3800 134392 3806
rect 134340 3742 134392 3748
rect 134444 3738 134472 75140
rect 134536 5302 134564 75140
rect 134524 5296 134576 5302
rect 134524 5238 134576 5244
rect 134432 3732 134484 3738
rect 134432 3674 134484 3680
rect 134628 3670 134656 75140
rect 134720 72554 134748 75140
rect 134708 72548 134760 72554
rect 134708 72490 134760 72496
rect 134812 10878 134840 75140
rect 134800 10872 134852 10878
rect 134800 10814 134852 10820
rect 134904 9654 134932 75140
rect 134996 72049 135024 75140
rect 135088 72185 135116 75140
rect 135074 72176 135130 72185
rect 135074 72111 135130 72120
rect 134982 72040 135038 72049
rect 134982 71975 135038 71984
rect 135180 71913 135208 75140
rect 135166 71904 135222 71913
rect 135166 71839 135222 71848
rect 135272 25498 135300 75140
rect 135364 32978 135392 75140
rect 135352 32972 135404 32978
rect 135352 32914 135404 32920
rect 135260 25492 135312 25498
rect 135260 25434 135312 25440
rect 134892 9648 134944 9654
rect 134892 9590 134944 9596
rect 135456 9586 135484 75140
rect 135548 26246 135576 75140
rect 135640 32910 135668 75140
rect 135732 72486 135760 75140
rect 135720 72480 135772 72486
rect 135720 72422 135772 72428
rect 135628 32904 135680 32910
rect 135628 32846 135680 32852
rect 135536 26240 135588 26246
rect 135536 26182 135588 26188
rect 135824 26178 135852 75140
rect 135916 32842 135944 75140
rect 135904 32836 135956 32842
rect 135904 32778 135956 32784
rect 135812 26172 135864 26178
rect 135812 26114 135864 26120
rect 135444 9580 135496 9586
rect 135444 9522 135496 9528
rect 136008 9518 136036 75140
rect 136100 27538 136128 75140
rect 136192 71913 136220 75140
rect 136284 73030 136312 75140
rect 136272 73024 136324 73030
rect 136272 72966 136324 72972
rect 136376 72049 136404 75140
rect 136468 72185 136496 75140
rect 136454 72176 136510 72185
rect 136454 72111 136510 72120
rect 136362 72040 136418 72049
rect 136362 71975 136418 71984
rect 136560 71913 136588 75140
rect 136178 71904 136234 71913
rect 136546 71904 136602 71913
rect 136178 71839 136234 71848
rect 136272 71868 136324 71874
rect 136652 71874 136680 75140
rect 136546 71839 136602 71848
rect 136640 71868 136692 71874
rect 136272 71810 136324 71816
rect 136640 71810 136692 71816
rect 136284 64874 136312 71810
rect 136192 64846 136312 64874
rect 136088 27532 136140 27538
rect 136088 27474 136140 27480
rect 135996 9512 136048 9518
rect 135996 9454 136048 9460
rect 135260 3936 135312 3942
rect 135260 3878 135312 3884
rect 134616 3664 134668 3670
rect 134616 3606 134668 3612
rect 133512 3460 133564 3466
rect 133512 3402 133564 3408
rect 134156 3392 134208 3398
rect 134156 3334 134208 3340
rect 134168 480 134196 3334
rect 135272 480 135300 3878
rect 136192 2990 136220 64846
rect 136744 32774 136772 75140
rect 136836 73166 136864 75140
rect 136824 73160 136876 73166
rect 136824 73102 136876 73108
rect 136732 32768 136784 32774
rect 136732 32710 136784 32716
rect 136928 27470 136956 75140
rect 137020 32706 137048 75140
rect 137008 32700 137060 32706
rect 137008 32642 137060 32648
rect 136916 27464 136968 27470
rect 136916 27406 136968 27412
rect 137112 10810 137140 75140
rect 137204 27334 137232 75140
rect 137192 27328 137244 27334
rect 137192 27270 137244 27276
rect 137100 10804 137152 10810
rect 137100 10746 137152 10752
rect 137296 5234 137324 75140
rect 137388 10742 137416 75140
rect 137480 27266 137508 75140
rect 137572 32638 137600 75140
rect 137664 73098 137692 75140
rect 137652 73092 137704 73098
rect 137652 73034 137704 73040
rect 137756 72978 137784 75140
rect 137664 72950 137784 72978
rect 137664 72418 137692 72950
rect 137744 72616 137796 72622
rect 137744 72558 137796 72564
rect 137652 72412 137704 72418
rect 137652 72354 137704 72360
rect 137652 71800 137704 71806
rect 137652 71742 137704 71748
rect 137560 32632 137612 32638
rect 137560 32574 137612 32580
rect 137468 27260 137520 27266
rect 137468 27202 137520 27208
rect 137664 16574 137692 71742
rect 137756 69578 137784 72558
rect 137848 72049 137876 75140
rect 137834 72040 137890 72049
rect 137834 71975 137890 71984
rect 137940 71913 137968 75140
rect 137926 71904 137982 71913
rect 137926 71839 137982 71848
rect 138032 69714 138060 75140
rect 138124 69834 138152 75140
rect 138112 69828 138164 69834
rect 138112 69770 138164 69776
rect 138032 69686 138152 69714
rect 137756 69550 138060 69578
rect 137664 16546 137784 16574
rect 137376 10736 137428 10742
rect 137376 10678 137428 10684
rect 137284 5228 137336 5234
rect 137284 5170 137336 5176
rect 137650 3632 137706 3641
rect 137650 3567 137706 3576
rect 136456 3324 136508 3330
rect 136456 3266 136508 3272
rect 136180 2984 136232 2990
rect 136180 2926 136232 2932
rect 136468 480 136496 3266
rect 137664 480 137692 3567
rect 137756 3398 137784 16546
rect 138032 6914 138060 69550
rect 138124 28150 138152 69686
rect 138112 28144 138164 28150
rect 138112 28086 138164 28092
rect 138216 12238 138244 75140
rect 138308 28218 138336 75140
rect 138400 34406 138428 75140
rect 138388 34400 138440 34406
rect 138388 34342 138440 34348
rect 138296 28212 138348 28218
rect 138296 28154 138348 28160
rect 138204 12232 138256 12238
rect 138204 12174 138256 12180
rect 138492 12170 138520 75140
rect 138584 27198 138612 75140
rect 138676 34338 138704 75140
rect 138664 34332 138716 34338
rect 138664 34274 138716 34280
rect 138572 27192 138624 27198
rect 138572 27134 138624 27140
rect 138480 12164 138532 12170
rect 138480 12106 138532 12112
rect 138768 12102 138796 75140
rect 138860 72690 138888 75140
rect 138848 72684 138900 72690
rect 138848 72626 138900 72632
rect 138952 71913 138980 75140
rect 139044 72049 139072 75140
rect 139030 72040 139086 72049
rect 139030 71975 139086 71984
rect 139136 71913 139164 75140
rect 139228 72622 139256 75140
rect 139216 72616 139268 72622
rect 139216 72558 139268 72564
rect 139320 72185 139348 75140
rect 139306 72176 139362 72185
rect 139306 72111 139362 72120
rect 138938 71904 138994 71913
rect 138938 71839 138994 71848
rect 139122 71904 139178 71913
rect 139122 71839 139178 71848
rect 138848 69828 138900 69834
rect 138848 69770 138900 69776
rect 138860 34474 138888 69770
rect 138848 34468 138900 34474
rect 138848 34410 138900 34416
rect 139412 28966 139440 75140
rect 139400 28960 139452 28966
rect 139400 28902 139452 28908
rect 139504 20466 139532 75140
rect 139492 20460 139544 20466
rect 139492 20402 139544 20408
rect 139596 13462 139624 75140
rect 139688 27130 139716 75140
rect 139780 34270 139808 75140
rect 139768 34264 139820 34270
rect 139768 34206 139820 34212
rect 139676 27124 139728 27130
rect 139676 27066 139728 27072
rect 139584 13456 139636 13462
rect 139584 13398 139636 13404
rect 138756 12096 138808 12102
rect 138756 12038 138808 12044
rect 138032 6886 138888 6914
rect 137744 3392 137796 3398
rect 137744 3334 137796 3340
rect 138860 480 138888 6886
rect 139872 6798 139900 75140
rect 139964 26110 139992 75140
rect 139952 26104 140004 26110
rect 139952 26046 140004 26052
rect 140056 20398 140084 75140
rect 140044 20392 140096 20398
rect 140044 20334 140096 20340
rect 140148 13394 140176 75140
rect 140240 28830 140268 75140
rect 140332 72185 140360 75140
rect 140318 72176 140374 72185
rect 140318 72111 140374 72120
rect 140424 71913 140452 75140
rect 140516 72758 140544 75140
rect 140504 72752 140556 72758
rect 140504 72694 140556 72700
rect 140608 72049 140636 75140
rect 140594 72040 140650 72049
rect 140594 71975 140650 71984
rect 140700 71913 140728 75140
rect 140410 71904 140466 71913
rect 140410 71839 140466 71848
rect 140686 71904 140742 71913
rect 140686 71839 140742 71848
rect 140228 28824 140280 28830
rect 140228 28766 140280 28772
rect 140792 28762 140820 75140
rect 140884 34202 140912 75140
rect 140976 74254 141004 75140
rect 140964 74248 141016 74254
rect 140964 74190 141016 74196
rect 140872 34196 140924 34202
rect 140872 34138 140924 34144
rect 140780 28756 140832 28762
rect 140780 28698 140832 28704
rect 141068 28626 141096 75140
rect 141056 28620 141108 28626
rect 141056 28562 141108 28568
rect 141160 19106 141188 75140
rect 141148 19100 141200 19106
rect 141148 19042 141200 19048
rect 141252 14890 141280 75140
rect 141344 24818 141372 75140
rect 141436 34134 141464 75140
rect 141424 34128 141476 34134
rect 141424 34070 141476 34076
rect 141332 24812 141384 24818
rect 141332 24754 141384 24760
rect 141240 14884 141292 14890
rect 141240 14826 141292 14832
rect 141528 14822 141556 75140
rect 141620 72962 141648 75140
rect 141608 72956 141660 72962
rect 141608 72898 141660 72904
rect 141712 20330 141740 75140
rect 141804 74934 141832 75140
rect 141792 74928 141844 74934
rect 141792 74870 141844 74876
rect 141896 26042 141924 75140
rect 141988 72049 142016 75140
rect 141974 72040 142030 72049
rect 141974 71975 142030 71984
rect 142080 71913 142108 75140
rect 142172 72894 142200 75140
rect 142160 72888 142212 72894
rect 142160 72830 142212 72836
rect 142066 71904 142122 71913
rect 142066 71839 142122 71848
rect 142264 32570 142292 75140
rect 142252 32564 142304 32570
rect 142252 32506 142304 32512
rect 141884 26036 141936 26042
rect 141884 25978 141936 25984
rect 141700 20324 141752 20330
rect 141700 20266 141752 20272
rect 141516 14816 141568 14822
rect 141516 14758 141568 14764
rect 142356 14754 142384 75140
rect 142344 14748 142396 14754
rect 142344 14690 142396 14696
rect 140136 13388 140188 13394
rect 140136 13330 140188 13336
rect 142448 7954 142476 75140
rect 142540 34066 142568 75140
rect 142528 34060 142580 34066
rect 142528 34002 142580 34008
rect 142632 14686 142660 75140
rect 142724 72146 142752 75140
rect 142712 72140 142764 72146
rect 142712 72082 142764 72088
rect 142816 17678 142844 75140
rect 142804 17672 142856 17678
rect 142804 17614 142856 17620
rect 142908 16386 142936 75140
rect 142896 16380 142948 16386
rect 142896 16322 142948 16328
rect 142620 14680 142672 14686
rect 142620 14622 142672 14628
rect 143000 10674 143028 75140
rect 143092 33998 143120 75140
rect 143184 71913 143212 75140
rect 143276 72185 143304 75140
rect 143262 72176 143318 72185
rect 143262 72111 143318 72120
rect 143368 72049 143396 75140
rect 143354 72040 143410 72049
rect 143354 71975 143410 71984
rect 143460 71913 143488 75140
rect 143170 71904 143226 71913
rect 143170 71839 143226 71848
rect 143446 71904 143502 71913
rect 143446 71839 143502 71848
rect 143172 71800 143224 71806
rect 143172 71742 143224 71748
rect 143080 33992 143132 33998
rect 143080 33934 143132 33940
rect 143184 27606 143212 71742
rect 143172 27600 143224 27606
rect 143172 27542 143224 27548
rect 143552 24750 143580 75140
rect 143644 33930 143672 75140
rect 143736 74186 143764 75140
rect 143724 74180 143776 74186
rect 143724 74122 143776 74128
rect 143632 33924 143684 33930
rect 143632 33866 143684 33872
rect 143540 24744 143592 24750
rect 143540 24686 143592 24692
rect 142988 10668 143040 10674
rect 142988 10610 143040 10616
rect 142436 7948 142488 7954
rect 142436 7890 142488 7896
rect 139860 6792 139912 6798
rect 139860 6734 139912 6740
rect 143828 6730 143856 75140
rect 143920 16318 143948 75140
rect 143908 16312 143960 16318
rect 143908 16254 143960 16260
rect 144012 16250 144040 75140
rect 144000 16244 144052 16250
rect 144000 16186 144052 16192
rect 144104 7886 144132 75140
rect 144196 33862 144224 75140
rect 144184 33856 144236 33862
rect 144184 33798 144236 33804
rect 144288 16182 144316 75140
rect 144380 25974 144408 75140
rect 144368 25968 144420 25974
rect 144368 25910 144420 25916
rect 144276 16176 144328 16182
rect 144276 16118 144328 16124
rect 144472 10606 144500 75140
rect 144564 71913 144592 75140
rect 144656 72049 144684 75140
rect 144748 72185 144776 75140
rect 144734 72176 144790 72185
rect 144734 72111 144790 72120
rect 144642 72040 144698 72049
rect 144642 71975 144698 71984
rect 144840 71913 144868 75140
rect 144550 71904 144606 71913
rect 144550 71839 144606 71848
rect 144826 71904 144882 71913
rect 144826 71839 144882 71848
rect 144932 30258 144960 75140
rect 145024 33794 145052 75140
rect 145116 74866 145144 75140
rect 145104 74860 145156 74866
rect 145104 74802 145156 74808
rect 145012 33788 145064 33794
rect 145012 33730 145064 33736
rect 144920 30252 144972 30258
rect 144920 30194 144972 30200
rect 145208 30190 145236 75140
rect 145300 35154 145328 75140
rect 145288 35148 145340 35154
rect 145288 35090 145340 35096
rect 145196 30184 145248 30190
rect 145196 30126 145248 30132
rect 144460 10600 144512 10606
rect 144460 10542 144512 10548
rect 145392 9450 145420 75140
rect 145484 72282 145512 75140
rect 145472 72276 145524 72282
rect 145472 72218 145524 72224
rect 145576 35902 145604 75140
rect 145564 35896 145616 35902
rect 145564 35838 145616 35844
rect 145380 9444 145432 9450
rect 145380 9386 145432 9392
rect 145668 9382 145696 75140
rect 145656 9376 145708 9382
rect 145656 9318 145708 9324
rect 145760 9314 145788 75140
rect 145852 71806 145880 75140
rect 145840 71800 145892 71806
rect 145840 71742 145892 71748
rect 145944 10538 145972 75140
rect 146036 72185 146064 75140
rect 146022 72176 146078 72185
rect 146022 72111 146078 72120
rect 146024 72072 146076 72078
rect 146024 72014 146076 72020
rect 146036 27402 146064 72014
rect 146128 71913 146156 75140
rect 146220 72049 146248 75140
rect 146206 72040 146262 72049
rect 146206 71975 146262 71984
rect 146114 71904 146170 71913
rect 146114 71839 146170 71848
rect 146024 27396 146076 27402
rect 146024 27338 146076 27344
rect 145932 10532 145984 10538
rect 145932 10474 145984 10480
rect 146312 10470 146340 75140
rect 146404 35766 146432 75140
rect 146496 74118 146524 75140
rect 146484 74112 146536 74118
rect 146484 74054 146536 74060
rect 146484 72684 146536 72690
rect 146484 72626 146536 72632
rect 146496 72214 146524 72626
rect 146484 72208 146536 72214
rect 146484 72150 146536 72156
rect 146392 35760 146444 35766
rect 146392 35702 146444 35708
rect 146588 12034 146616 75140
rect 146680 35698 146708 75140
rect 146772 74730 146800 75140
rect 146760 74724 146812 74730
rect 146760 74666 146812 74672
rect 146760 72956 146812 72962
rect 146760 72898 146812 72904
rect 146772 71942 146800 72898
rect 146760 71936 146812 71942
rect 146760 71878 146812 71884
rect 146668 35692 146720 35698
rect 146668 35634 146720 35640
rect 146864 13326 146892 75140
rect 146956 35630 146984 75140
rect 146944 35624 146996 35630
rect 146944 35566 146996 35572
rect 147048 17610 147076 75140
rect 147036 17604 147088 17610
rect 147036 17546 147088 17552
rect 146852 13320 146904 13326
rect 146852 13262 146904 13268
rect 147140 13258 147168 75140
rect 147232 20262 147260 75140
rect 147324 71913 147352 75140
rect 147416 72185 147444 75140
rect 147508 72321 147536 75140
rect 147494 72312 147550 72321
rect 147494 72247 147550 72256
rect 147402 72176 147458 72185
rect 147402 72111 147458 72120
rect 147600 72049 147628 75140
rect 147586 72040 147642 72049
rect 147586 71975 147642 71984
rect 147310 71904 147366 71913
rect 147310 71839 147366 71848
rect 147312 71800 147364 71806
rect 147312 71742 147364 71748
rect 147324 35834 147352 71742
rect 147312 35828 147364 35834
rect 147312 35770 147364 35776
rect 147220 20256 147272 20262
rect 147220 20198 147272 20204
rect 147128 13252 147180 13258
rect 147128 13194 147180 13200
rect 146576 12028 146628 12034
rect 146576 11970 146628 11976
rect 146300 10464 146352 10470
rect 146300 10406 146352 10412
rect 145748 9308 145800 9314
rect 145748 9250 145800 9256
rect 144092 7880 144144 7886
rect 144092 7822 144144 7828
rect 147692 7818 147720 75140
rect 147784 35562 147812 75140
rect 147876 74050 147904 75140
rect 147864 74044 147916 74050
rect 147864 73986 147916 73992
rect 147772 35556 147824 35562
rect 147772 35498 147824 35504
rect 147968 9246 147996 75140
rect 148060 22098 148088 75140
rect 148048 22092 148100 22098
rect 148048 22034 148100 22040
rect 147956 9240 148008 9246
rect 147956 9182 148008 9188
rect 148152 9178 148180 75140
rect 148244 11966 148272 75140
rect 148336 27062 148364 75140
rect 148324 27056 148376 27062
rect 148324 26998 148376 27004
rect 148232 11960 148284 11966
rect 148232 11902 148284 11908
rect 148428 11898 148456 75140
rect 148520 16114 148548 75140
rect 148612 35494 148640 75140
rect 148704 72729 148732 75140
rect 148690 72720 148746 72729
rect 148690 72655 148746 72664
rect 148796 72457 148824 75140
rect 148888 72865 148916 75140
rect 148874 72856 148930 72865
rect 148874 72791 148930 72800
rect 148980 72729 149008 75140
rect 148966 72720 149022 72729
rect 148966 72655 149022 72664
rect 148782 72448 148838 72457
rect 148782 72383 148838 72392
rect 148600 35488 148652 35494
rect 148600 35430 148652 35436
rect 148508 16108 148560 16114
rect 148508 16050 148560 16056
rect 149072 16046 149100 75140
rect 149164 72826 149192 75140
rect 149152 72820 149204 72826
rect 149152 72762 149204 72768
rect 149152 72548 149204 72554
rect 149152 72490 149204 72496
rect 149060 16040 149112 16046
rect 149060 15982 149112 15988
rect 148416 11892 148468 11898
rect 148416 11834 148468 11840
rect 148140 9172 148192 9178
rect 148140 9114 148192 9120
rect 147680 7812 147732 7818
rect 147680 7754 147732 7760
rect 143816 6724 143868 6730
rect 143816 6666 143868 6672
rect 142436 5432 142488 5438
rect 142436 5374 142488 5380
rect 140042 3496 140098 3505
rect 140042 3431 140098 3440
rect 140056 480 140084 3431
rect 141240 2984 141292 2990
rect 141240 2926 141292 2932
rect 141252 480 141280 2926
rect 142448 480 142476 5374
rect 144736 5364 144788 5370
rect 144736 5306 144788 5312
rect 143540 4140 143592 4146
rect 143540 4082 143592 4088
rect 143552 480 143580 4082
rect 144748 480 144776 5306
rect 148324 5160 148376 5166
rect 148324 5102 148376 5108
rect 146944 4072 146996 4078
rect 146944 4014 146996 4020
rect 145932 4004 145984 4010
rect 145932 3946 145984 3952
rect 145944 480 145972 3946
rect 146956 3398 146984 4014
rect 147128 3596 147180 3602
rect 147128 3538 147180 3544
rect 146944 3392 146996 3398
rect 146944 3334 146996 3340
rect 147140 480 147168 3538
rect 148336 480 148364 5102
rect 149164 3330 149192 72490
rect 149256 11830 149284 75140
rect 149348 25906 149376 75140
rect 149440 35358 149468 75140
rect 149428 35352 149480 35358
rect 149428 35294 149480 35300
rect 149336 25900 149388 25906
rect 149336 25842 149388 25848
rect 149532 18970 149560 75140
rect 149520 18964 149572 18970
rect 149520 18906 149572 18912
rect 149624 14618 149652 75140
rect 149716 71806 149744 75140
rect 149704 71800 149756 71806
rect 149704 71742 149756 71748
rect 149612 14612 149664 14618
rect 149612 14554 149664 14560
rect 149808 13190 149836 75140
rect 149796 13184 149848 13190
rect 149796 13126 149848 13132
rect 149244 11824 149296 11830
rect 149244 11766 149296 11772
rect 149900 5166 149928 75140
rect 149992 72729 150020 75140
rect 149978 72720 150034 72729
rect 149978 72655 150034 72664
rect 150084 72457 150112 75140
rect 150176 72593 150204 75140
rect 150268 72690 150296 75140
rect 150360 72865 150388 75140
rect 150346 72856 150402 72865
rect 150346 72791 150402 72800
rect 150256 72684 150308 72690
rect 150256 72626 150308 72632
rect 150162 72584 150218 72593
rect 150162 72519 150218 72528
rect 150070 72448 150126 72457
rect 150070 72383 150126 72392
rect 150164 72208 150216 72214
rect 150164 72150 150216 72156
rect 150176 28082 150204 72150
rect 150452 28422 150480 75140
rect 150440 28416 150492 28422
rect 150440 28358 150492 28364
rect 150164 28076 150216 28082
rect 150164 28018 150216 28024
rect 150544 25838 150572 75140
rect 150636 74934 150664 75140
rect 150624 74928 150676 74934
rect 150624 74870 150676 74876
rect 150728 30122 150756 75140
rect 150820 72418 150848 75140
rect 150808 72412 150860 72418
rect 150808 72354 150860 72360
rect 150716 30116 150768 30122
rect 150716 30058 150768 30064
rect 150532 25832 150584 25838
rect 150532 25774 150584 25780
rect 150912 18902 150940 75140
rect 150900 18896 150952 18902
rect 150900 18838 150952 18844
rect 151004 13122 151032 75140
rect 150992 13116 151044 13122
rect 150992 13058 151044 13064
rect 151096 6662 151124 75140
rect 151188 18834 151216 75140
rect 151280 72622 151308 75140
rect 151268 72616 151320 72622
rect 151268 72558 151320 72564
rect 151372 71874 151400 75140
rect 151360 71868 151412 71874
rect 151360 71810 151412 71816
rect 151176 18828 151228 18834
rect 151176 18770 151228 18776
rect 151464 14550 151492 75140
rect 151556 72729 151584 75140
rect 151648 72865 151676 75140
rect 151634 72856 151690 72865
rect 151634 72791 151690 72800
rect 151636 72752 151688 72758
rect 151542 72720 151598 72729
rect 151636 72694 151688 72700
rect 151542 72655 151598 72664
rect 151544 71936 151596 71942
rect 151544 71878 151596 71884
rect 151556 28694 151584 71878
rect 151648 28898 151676 72694
rect 151740 72457 151768 75140
rect 151726 72448 151782 72457
rect 151726 72383 151782 72392
rect 151832 71942 151860 75140
rect 151924 72010 151952 75140
rect 152016 73982 152044 75140
rect 152004 73976 152056 73982
rect 152004 73918 152056 73924
rect 152004 73364 152056 73370
rect 152004 73306 152056 73312
rect 152016 72758 152044 73306
rect 152004 72752 152056 72758
rect 152004 72694 152056 72700
rect 151912 72004 151964 72010
rect 151912 71946 151964 71952
rect 151820 71936 151872 71942
rect 151820 71878 151872 71884
rect 151636 28892 151688 28898
rect 151636 28834 151688 28840
rect 151544 28688 151596 28694
rect 151544 28630 151596 28636
rect 151452 14544 151504 14550
rect 151452 14486 151504 14492
rect 152108 9110 152136 75140
rect 152200 73370 152228 75140
rect 152188 73364 152240 73370
rect 152188 73306 152240 73312
rect 152188 73228 152240 73234
rect 152188 73170 152240 73176
rect 152200 72350 152228 73170
rect 152188 72344 152240 72350
rect 152188 72286 152240 72292
rect 152292 20194 152320 75140
rect 152280 20188 152332 20194
rect 152280 20130 152332 20136
rect 152096 9104 152148 9110
rect 152096 9046 152148 9052
rect 151084 6656 151136 6662
rect 151084 6598 151136 6604
rect 152384 6594 152412 75140
rect 152476 36582 152504 75140
rect 152464 36576 152516 36582
rect 152464 36518 152516 36524
rect 152568 20126 152596 75140
rect 152556 20120 152608 20126
rect 152556 20062 152608 20068
rect 152660 10402 152688 75140
rect 152752 73234 152780 75140
rect 152740 73228 152792 73234
rect 152740 73170 152792 73176
rect 152740 72888 152792 72894
rect 152740 72830 152792 72836
rect 152752 64874 152780 72830
rect 152844 72593 152872 75140
rect 152936 72865 152964 75140
rect 152922 72856 152978 72865
rect 152922 72791 152978 72800
rect 153028 72729 153056 75140
rect 153120 73001 153148 75140
rect 153106 72992 153162 73001
rect 153106 72927 153162 72936
rect 153014 72720 153070 72729
rect 153014 72655 153070 72664
rect 152830 72584 152886 72593
rect 152830 72519 152886 72528
rect 153108 72548 153160 72554
rect 153108 72490 153160 72496
rect 152924 72412 152976 72418
rect 152924 72354 152976 72360
rect 152752 64846 152872 64874
rect 152844 28558 152872 64846
rect 152832 28552 152884 28558
rect 152832 28494 152884 28500
rect 152936 28354 152964 72354
rect 153016 72072 153068 72078
rect 153016 72014 153068 72020
rect 153028 28490 153056 72014
rect 153120 40730 153148 72490
rect 153108 40724 153160 40730
rect 153108 40666 153160 40672
rect 153016 28484 153068 28490
rect 153016 28426 153068 28432
rect 152924 28348 152976 28354
rect 152924 28290 152976 28296
rect 153212 24682 153240 75140
rect 153304 72078 153332 75140
rect 153396 74458 153424 75140
rect 153384 74452 153436 74458
rect 153384 74394 153436 74400
rect 153292 72072 153344 72078
rect 153292 72014 153344 72020
rect 153200 24676 153252 24682
rect 153200 24618 153252 24624
rect 152648 10396 152700 10402
rect 152648 10338 152700 10344
rect 153488 9042 153516 75140
rect 153476 9036 153528 9042
rect 153476 8978 153528 8984
rect 153580 8974 153608 75140
rect 153672 20058 153700 75140
rect 153764 25770 153792 75140
rect 153856 72282 153884 75140
rect 153844 72276 153896 72282
rect 153844 72218 153896 72224
rect 153752 25764 153804 25770
rect 153752 25706 153804 25712
rect 153660 20052 153712 20058
rect 153660 19994 153712 20000
rect 153948 15978 153976 75140
rect 153936 15972 153988 15978
rect 153936 15914 153988 15920
rect 153568 8968 153620 8974
rect 153568 8910 153620 8916
rect 154040 7750 154068 75140
rect 154132 72865 154160 75140
rect 154118 72856 154174 72865
rect 154118 72791 154174 72800
rect 154224 72729 154252 75140
rect 154210 72720 154266 72729
rect 154210 72655 154266 72664
rect 154212 72616 154264 72622
rect 154212 72558 154264 72564
rect 154224 30054 154252 72558
rect 154316 72457 154344 75140
rect 154408 72962 154436 75140
rect 154396 72956 154448 72962
rect 154396 72898 154448 72904
rect 154396 72820 154448 72826
rect 154396 72762 154448 72768
rect 154302 72448 154358 72457
rect 154408 72434 154436 72762
rect 154500 72593 154528 75140
rect 154486 72584 154542 72593
rect 154486 72519 154542 72528
rect 154408 72406 154528 72434
rect 154302 72383 154358 72392
rect 154396 72208 154448 72214
rect 154396 72150 154448 72156
rect 154408 64874 154436 72150
rect 154316 64846 154436 64874
rect 154316 30326 154344 64846
rect 154500 35426 154528 72406
rect 154488 35420 154540 35426
rect 154488 35362 154540 35368
rect 154304 30320 154356 30326
rect 154304 30262 154356 30268
rect 154212 30048 154264 30054
rect 154212 29990 154264 29996
rect 154592 26994 154620 75140
rect 154580 26988 154632 26994
rect 154580 26930 154632 26936
rect 154684 21962 154712 75140
rect 154776 74497 154804 75140
rect 154762 74488 154818 74497
rect 154762 74423 154818 74432
rect 154672 21956 154724 21962
rect 154672 21898 154724 21904
rect 154868 17542 154896 75140
rect 154960 72146 154988 75140
rect 154948 72140 155000 72146
rect 154948 72082 155000 72088
rect 155052 21894 155080 75140
rect 155144 29918 155172 75140
rect 155132 29912 155184 29918
rect 155132 29854 155184 29860
rect 155040 21888 155092 21894
rect 155040 21830 155092 21836
rect 155236 21826 155264 75140
rect 155224 21820 155276 21826
rect 155224 21762 155276 21768
rect 154856 17536 154908 17542
rect 154856 17478 154908 17484
rect 155328 17474 155356 75140
rect 155316 17468 155368 17474
rect 155316 17410 155368 17416
rect 155420 17406 155448 75140
rect 155512 73001 155540 75140
rect 155498 72992 155554 73001
rect 155498 72927 155554 72936
rect 155408 17400 155460 17406
rect 155408 17342 155460 17348
rect 155604 17338 155632 75140
rect 155696 72321 155724 75140
rect 155788 72457 155816 75140
rect 155880 72729 155908 75140
rect 155866 72720 155922 72729
rect 155866 72655 155922 72664
rect 155774 72448 155830 72457
rect 155774 72383 155830 72392
rect 155682 72312 155738 72321
rect 155682 72247 155738 72256
rect 155776 72004 155828 72010
rect 155776 71946 155828 71952
rect 155788 36650 155816 71946
rect 155776 36644 155828 36650
rect 155776 36586 155828 36592
rect 155972 29782 156000 75140
rect 156064 72894 156092 75140
rect 156156 74633 156184 75140
rect 156142 74624 156198 74633
rect 156142 74559 156198 74568
rect 156052 72888 156104 72894
rect 156052 72830 156104 72836
rect 155960 29776 156012 29782
rect 155960 29718 156012 29724
rect 156248 29714 156276 75140
rect 156236 29708 156288 29714
rect 156236 29650 156288 29656
rect 156340 21758 156368 75140
rect 156328 21752 156380 21758
rect 156328 21694 156380 21700
rect 156432 21690 156460 75140
rect 156420 21684 156472 21690
rect 156420 21626 156472 21632
rect 155592 17332 155644 17338
rect 155592 17274 155644 17280
rect 156524 10334 156552 75140
rect 156616 72826 156644 75140
rect 156604 72820 156656 72826
rect 156604 72762 156656 72768
rect 156708 18766 156736 75140
rect 156800 29646 156828 75140
rect 156892 72729 156920 75140
rect 156984 72865 157012 75140
rect 156970 72856 157026 72865
rect 156970 72791 157026 72800
rect 156878 72720 156934 72729
rect 156878 72655 156934 72664
rect 157076 72593 157104 75140
rect 157062 72584 157118 72593
rect 157062 72519 157118 72528
rect 157062 72312 157118 72321
rect 157062 72247 157118 72256
rect 156972 71800 157024 71806
rect 156972 71742 157024 71748
rect 156788 29640 156840 29646
rect 156788 29582 156840 29588
rect 156984 22030 157012 71742
rect 157076 29850 157104 72247
rect 157168 72049 157196 75140
rect 157260 72729 157288 75140
rect 157246 72720 157302 72729
rect 157246 72655 157302 72664
rect 157154 72040 157210 72049
rect 157154 71975 157210 71984
rect 157156 71936 157208 71942
rect 157156 71878 157208 71884
rect 157168 64874 157196 71878
rect 157168 64846 157288 64874
rect 157260 29986 157288 64846
rect 157248 29980 157300 29986
rect 157248 29922 157300 29928
rect 157064 29844 157116 29850
rect 157064 29786 157116 29792
rect 157352 23458 157380 75140
rect 157444 72758 157472 75140
rect 157536 74390 157564 75140
rect 157524 74384 157576 74390
rect 157524 74326 157576 74332
rect 157432 72752 157484 72758
rect 157432 72694 157484 72700
rect 157524 72480 157576 72486
rect 157524 72422 157576 72428
rect 157536 71942 157564 72422
rect 157524 71936 157576 71942
rect 157524 71878 157576 71884
rect 157628 31754 157656 75140
rect 157616 31748 157668 31754
rect 157616 31690 157668 31696
rect 157340 23452 157392 23458
rect 157340 23394 157392 23400
rect 156972 22024 157024 22030
rect 156972 21966 157024 21972
rect 156696 18760 156748 18766
rect 156696 18702 156748 18708
rect 157720 12306 157748 75140
rect 157812 73846 157840 75140
rect 157800 73840 157852 73846
rect 157800 73782 157852 73788
rect 157798 72040 157854 72049
rect 157798 71975 157854 71984
rect 157812 35222 157840 71975
rect 157800 35216 157852 35222
rect 157800 35158 157852 35164
rect 157904 14482 157932 75140
rect 157996 26926 158024 75140
rect 157984 26920 158036 26926
rect 157984 26862 158036 26868
rect 158088 19990 158116 75140
rect 158180 31686 158208 75140
rect 158272 72690 158300 75140
rect 158364 72865 158392 75140
rect 158350 72856 158406 72865
rect 158350 72791 158406 72800
rect 158260 72684 158312 72690
rect 158260 72626 158312 72632
rect 158260 72548 158312 72554
rect 158260 72490 158312 72496
rect 158272 64874 158300 72490
rect 158456 72457 158484 75140
rect 158548 72729 158576 75140
rect 158534 72720 158590 72729
rect 158534 72655 158590 72664
rect 158640 72593 158668 75140
rect 158626 72584 158682 72593
rect 158626 72519 158682 72528
rect 158442 72448 158498 72457
rect 158442 72383 158498 72392
rect 158444 71868 158496 71874
rect 158444 71810 158496 71816
rect 158272 64846 158392 64874
rect 158364 35290 158392 64846
rect 158456 36718 158484 71810
rect 158444 36712 158496 36718
rect 158444 36654 158496 36660
rect 158352 35284 158404 35290
rect 158352 35226 158404 35232
rect 158168 31680 158220 31686
rect 158168 31622 158220 31628
rect 158732 31618 158760 75140
rect 158824 73137 158852 75140
rect 158810 73128 158866 73137
rect 158810 73063 158866 73072
rect 158812 72752 158864 72758
rect 158812 72694 158864 72700
rect 158824 72554 158852 72694
rect 158812 72548 158864 72554
rect 158812 72490 158864 72496
rect 158916 72185 158944 75140
rect 158902 72176 158958 72185
rect 158902 72111 158958 72120
rect 158720 31612 158772 31618
rect 158720 31554 158772 31560
rect 159008 21622 159036 75140
rect 159100 31550 159128 75140
rect 159088 31544 159140 31550
rect 159088 31486 159140 31492
rect 158996 21616 159048 21622
rect 158996 21558 159048 21564
rect 158076 19984 158128 19990
rect 158076 19926 158128 19932
rect 157892 14476 157944 14482
rect 157892 14418 157944 14424
rect 157708 12300 157760 12306
rect 157708 12242 157760 12248
rect 156512 10328 156564 10334
rect 156512 10270 156564 10276
rect 154028 7744 154080 7750
rect 154028 7686 154080 7692
rect 152372 6588 152424 6594
rect 152372 6530 152424 6536
rect 149888 5160 149940 5166
rect 149888 5102 149940 5108
rect 149520 5092 149572 5098
rect 149520 5034 149572 5040
rect 149152 3324 149204 3330
rect 149152 3266 149204 3272
rect 149532 480 149560 5034
rect 153016 5024 153068 5030
rect 153016 4966 153068 4972
rect 155406 4992 155462 5001
rect 151820 4956 151872 4962
rect 151820 4898 151872 4904
rect 150624 3528 150676 3534
rect 150624 3470 150676 3476
rect 150636 480 150664 3470
rect 151832 480 151860 4898
rect 153028 480 153056 4966
rect 155406 4927 155462 4936
rect 154212 3460 154264 3466
rect 154212 3402 154264 3408
rect 154224 480 154252 3402
rect 155420 480 155448 4927
rect 158904 4888 158956 4894
rect 156602 4856 156658 4865
rect 158904 4830 158956 4836
rect 156602 4791 156658 4800
rect 156616 480 156644 4791
rect 157798 3360 157854 3369
rect 157798 3295 157854 3304
rect 157812 480 157840 3295
rect 158916 480 158944 4830
rect 159192 3602 159220 75140
rect 159284 21554 159312 75140
rect 159272 21548 159324 21554
rect 159272 21490 159324 21496
rect 159376 11762 159404 75140
rect 159364 11756 159416 11762
rect 159364 11698 159416 11704
rect 159180 3596 159232 3602
rect 159180 3538 159232 3544
rect 159468 3534 159496 75140
rect 159560 21486 159588 75140
rect 159652 72457 159680 75140
rect 159638 72448 159694 72457
rect 159638 72383 159694 72392
rect 159548 21480 159600 21486
rect 159548 21422 159600 21428
rect 159456 3528 159508 3534
rect 159456 3470 159508 3476
rect 159744 3466 159772 75140
rect 159836 21418 159864 75140
rect 159928 72865 159956 75140
rect 159914 72856 159970 72865
rect 159914 72791 159970 72800
rect 160020 72729 160048 75140
rect 160006 72720 160062 72729
rect 160006 72655 160062 72664
rect 160112 23390 160140 75140
rect 160204 31414 160232 75140
rect 160296 72321 160324 75140
rect 160282 72312 160338 72321
rect 160282 72247 160338 72256
rect 160192 31408 160244 31414
rect 160192 31350 160244 31356
rect 160100 23384 160152 23390
rect 160100 23326 160152 23332
rect 160388 23322 160416 75140
rect 160376 23316 160428 23322
rect 160376 23258 160428 23264
rect 159824 21412 159876 21418
rect 159824 21354 159876 21360
rect 160480 5098 160508 75140
rect 160468 5092 160520 5098
rect 160468 5034 160520 5040
rect 160572 5030 160600 75140
rect 160664 23254 160692 75140
rect 160756 31346 160784 75140
rect 160744 31340 160796 31346
rect 160744 31282 160796 31288
rect 160652 23248 160704 23254
rect 160652 23190 160704 23196
rect 160560 5024 160612 5030
rect 160560 4966 160612 4972
rect 160100 4072 160152 4078
rect 160100 4014 160152 4020
rect 159732 3460 159784 3466
rect 159732 3402 159784 3408
rect 160112 480 160140 4014
rect 160848 3777 160876 75140
rect 160940 23186 160968 75140
rect 161032 72865 161060 75140
rect 161018 72856 161074 72865
rect 161018 72791 161074 72800
rect 161124 72729 161152 75140
rect 161110 72720 161166 72729
rect 161110 72655 161166 72664
rect 161216 72593 161244 75140
rect 161308 73137 161336 75140
rect 161294 73128 161350 73137
rect 161294 73063 161350 73072
rect 161400 72729 161428 75140
rect 161386 72720 161442 72729
rect 161386 72655 161442 72664
rect 161202 72584 161258 72593
rect 161202 72519 161258 72528
rect 161294 72448 161350 72457
rect 161294 72383 161350 72392
rect 161308 64874 161336 72383
rect 161124 64846 161336 64874
rect 161124 31482 161152 64846
rect 161112 31476 161164 31482
rect 161112 31418 161164 31424
rect 160928 23180 160980 23186
rect 160928 23122 160980 23128
rect 161492 23118 161520 75140
rect 161480 23112 161532 23118
rect 161480 23054 161532 23060
rect 161584 6458 161612 75140
rect 161676 74769 161704 75140
rect 161662 74760 161718 74769
rect 161662 74695 161718 74704
rect 161664 74520 161716 74526
rect 161662 74488 161664 74497
rect 161716 74488 161718 74497
rect 161662 74423 161718 74432
rect 161662 74216 161718 74225
rect 161662 74151 161718 74160
rect 161676 73846 161704 74151
rect 161664 73840 161716 73846
rect 161664 73782 161716 73788
rect 161664 73568 161716 73574
rect 161664 73510 161716 73516
rect 161676 73166 161704 73510
rect 161664 73160 161716 73166
rect 161664 73102 161716 73108
rect 161768 23050 161796 75140
rect 161860 31210 161888 75140
rect 161848 31204 161900 31210
rect 161848 31146 161900 31152
rect 161756 23044 161808 23050
rect 161756 22986 161808 22992
rect 161572 6452 161624 6458
rect 161572 6394 161624 6400
rect 161952 4962 161980 75140
rect 162044 22982 162072 75140
rect 162136 31074 162164 75140
rect 162124 31068 162176 31074
rect 162124 31010 162176 31016
rect 162032 22976 162084 22982
rect 162032 22918 162084 22924
rect 161940 4956 161992 4962
rect 161940 4898 161992 4904
rect 162228 4894 162256 75140
rect 162320 22914 162348 75140
rect 162412 73302 162440 75140
rect 162400 73296 162452 73302
rect 162400 73238 162452 73244
rect 162398 73128 162454 73137
rect 162398 73063 162454 73072
rect 162412 64874 162440 73063
rect 162504 72729 162532 75140
rect 162490 72720 162546 72729
rect 162490 72655 162546 72664
rect 162492 72616 162544 72622
rect 162490 72584 162492 72593
rect 162544 72584 162546 72593
rect 162490 72519 162546 72528
rect 162596 72457 162624 75140
rect 162688 72865 162716 75140
rect 162674 72856 162730 72865
rect 162674 72791 162730 72800
rect 162780 72729 162808 75140
rect 162766 72720 162822 72729
rect 162766 72655 162822 72664
rect 162582 72448 162638 72457
rect 162582 72383 162638 72392
rect 162412 64846 162624 64874
rect 162596 31278 162624 64846
rect 162584 31272 162636 31278
rect 162584 31214 162636 31220
rect 162872 24614 162900 75140
rect 162860 24608 162912 24614
rect 162860 24550 162912 24556
rect 162308 22908 162360 22914
rect 162308 22850 162360 22856
rect 162964 15910 162992 75140
rect 163056 73137 163084 75140
rect 163042 73128 163098 73137
rect 163042 73063 163098 73072
rect 163148 24546 163176 75140
rect 163136 24540 163188 24546
rect 163136 24482 163188 24488
rect 163240 18698 163268 75140
rect 163332 72321 163360 75140
rect 163318 72312 163374 72321
rect 163318 72247 163374 72256
rect 163424 24478 163452 75140
rect 163516 58682 163544 75140
rect 163504 58676 163556 58682
rect 163504 58618 163556 58624
rect 163412 24472 163464 24478
rect 163412 24414 163464 24420
rect 163228 18692 163280 18698
rect 163228 18634 163280 18640
rect 162952 15904 163004 15910
rect 162952 15846 163004 15852
rect 163608 6390 163636 75140
rect 163700 24410 163728 75140
rect 163688 24404 163740 24410
rect 163688 24346 163740 24352
rect 163792 19038 163820 75140
rect 163780 19032 163832 19038
rect 163780 18974 163832 18980
rect 163596 6384 163648 6390
rect 163596 6326 163648 6332
rect 163884 6322 163912 75140
rect 163976 72865 164004 75140
rect 163962 72856 164018 72865
rect 163962 72791 164018 72800
rect 164068 72593 164096 75140
rect 164160 72729 164188 75140
rect 164252 74769 164280 75140
rect 164238 74760 164294 74769
rect 164238 74695 164294 74704
rect 164238 74488 164294 74497
rect 164238 74423 164294 74432
rect 164146 72720 164202 72729
rect 164146 72655 164202 72664
rect 164054 72584 164110 72593
rect 164054 72519 164110 72528
rect 164252 24342 164280 74423
rect 164344 32502 164372 75140
rect 164436 74934 164464 75140
rect 164424 74928 164476 74934
rect 164424 74870 164476 74876
rect 164424 74588 164476 74594
rect 164424 74530 164476 74536
rect 164436 74390 164464 74530
rect 164424 74384 164476 74390
rect 164424 74326 164476 74332
rect 164422 74216 164478 74225
rect 164422 74151 164478 74160
rect 164436 73846 164464 74151
rect 164424 73840 164476 73846
rect 164424 73782 164476 73788
rect 164424 73160 164476 73166
rect 164424 73102 164476 73108
rect 164436 72758 164464 73102
rect 164424 72752 164476 72758
rect 164424 72694 164476 72700
rect 164332 32496 164384 32502
rect 164332 32438 164384 32444
rect 164240 24336 164292 24342
rect 164240 24278 164292 24284
rect 164528 24274 164556 75140
rect 164516 24268 164568 24274
rect 164516 24210 164568 24216
rect 164620 18630 164648 75140
rect 164712 74769 164740 75140
rect 164698 74760 164754 74769
rect 164698 74695 164754 74704
rect 164804 74610 164832 75140
rect 164712 74582 164832 74610
rect 164712 71448 164740 74582
rect 164896 74225 164924 75140
rect 164882 74216 164938 74225
rect 164882 74151 164938 74160
rect 164882 72856 164938 72865
rect 164882 72791 164938 72800
rect 164712 71420 164832 71448
rect 164698 71360 164754 71369
rect 164698 71295 164754 71304
rect 164608 18624 164660 18630
rect 164608 18566 164660 18572
rect 164712 7682 164740 71295
rect 164804 25702 164832 71420
rect 164792 25696 164844 25702
rect 164792 25638 164844 25644
rect 164896 17270 164924 72791
rect 164884 17264 164936 17270
rect 164884 17206 164936 17212
rect 164700 7676 164752 7682
rect 164700 7618 164752 7624
rect 164988 7614 165016 75140
rect 165080 74934 165108 75140
rect 165068 74928 165120 74934
rect 165068 74870 165120 74876
rect 165068 73092 165120 73098
rect 165068 73034 165120 73040
rect 165080 72554 165108 73034
rect 165068 72548 165120 72554
rect 165068 72490 165120 72496
rect 165172 22846 165200 75140
rect 165264 72729 165292 75140
rect 165356 72865 165384 75140
rect 165342 72856 165398 72865
rect 165342 72791 165398 72800
rect 165250 72720 165306 72729
rect 165250 72655 165306 72664
rect 165448 72593 165476 75140
rect 165540 72729 165568 75140
rect 165526 72720 165582 72729
rect 165526 72655 165582 72664
rect 165434 72584 165490 72593
rect 165434 72519 165490 72528
rect 165526 72312 165582 72321
rect 165526 72247 165582 72256
rect 165252 71936 165304 71942
rect 165252 71878 165304 71884
rect 165160 22840 165212 22846
rect 165160 22782 165212 22788
rect 164976 7608 165028 7614
rect 164976 7550 165028 7556
rect 163872 6316 163924 6322
rect 163872 6258 163924 6264
rect 162216 4888 162268 4894
rect 162216 4830 162268 4836
rect 163688 4820 163740 4826
rect 163688 4762 163740 4768
rect 161296 3936 161348 3942
rect 161296 3878 161348 3884
rect 160834 3768 160890 3777
rect 160834 3703 160890 3712
rect 161308 480 161336 3878
rect 162492 3868 162544 3874
rect 162492 3810 162544 3816
rect 162504 480 162532 3810
rect 163700 480 163728 4762
rect 164884 3800 164936 3806
rect 164884 3742 164936 3748
rect 164896 480 164924 3742
rect 165264 3262 165292 71878
rect 165540 70145 165568 72247
rect 165526 70136 165582 70145
rect 165526 70071 165582 70080
rect 165632 25634 165660 75140
rect 165620 25628 165672 25634
rect 165620 25570 165672 25576
rect 165724 24206 165752 75140
rect 165712 24200 165764 24206
rect 165712 24142 165764 24148
rect 165816 6254 165844 75140
rect 165908 24138 165936 75140
rect 166000 28286 166028 75140
rect 165988 28280 166040 28286
rect 165988 28222 166040 28228
rect 165896 24132 165948 24138
rect 165896 24074 165948 24080
rect 165804 6248 165856 6254
rect 165804 6190 165856 6196
rect 166092 6186 166120 75140
rect 166184 25566 166212 75140
rect 166276 32434 166304 75140
rect 166368 72865 166396 75140
rect 166354 72856 166410 72865
rect 166354 72791 166410 72800
rect 166356 72752 166408 72758
rect 166356 72694 166408 72700
rect 166264 32428 166316 32434
rect 166264 32370 166316 32376
rect 166368 31142 166396 72694
rect 166460 64874 166488 75140
rect 166552 72729 166580 75140
rect 166538 72720 166594 72729
rect 166538 72655 166594 72664
rect 166644 72486 166672 75140
rect 166736 73166 166764 75140
rect 166828 73409 166856 75140
rect 166814 73400 166870 73409
rect 166814 73335 166870 73344
rect 166724 73160 166776 73166
rect 166724 73102 166776 73108
rect 166632 72480 166684 72486
rect 166632 72422 166684 72428
rect 166920 71058 166948 75140
rect 167012 72026 167040 75140
rect 167104 74458 167132 75140
rect 167092 74452 167144 74458
rect 167092 74394 167144 74400
rect 167196 74390 167224 75140
rect 167288 74497 167316 75140
rect 167274 74488 167330 74497
rect 167274 74423 167330 74432
rect 167184 74384 167236 74390
rect 167380 74361 167408 75140
rect 167184 74326 167236 74332
rect 167366 74352 167422 74361
rect 167366 74287 167422 74296
rect 167472 74225 167500 75140
rect 167458 74216 167514 74225
rect 167458 74151 167514 74160
rect 167458 74080 167514 74089
rect 167458 74015 167514 74024
rect 167472 73574 167500 74015
rect 167564 73574 167592 75140
rect 167656 74644 167684 75140
rect 167748 74905 167776 75140
rect 167734 74896 167790 74905
rect 167734 74831 167790 74840
rect 167656 74616 167776 74644
rect 167644 74520 167696 74526
rect 167644 74462 167696 74468
rect 167460 73568 167512 73574
rect 167460 73510 167512 73516
rect 167552 73568 167604 73574
rect 167552 73510 167604 73516
rect 167274 72856 167330 72865
rect 167274 72791 167330 72800
rect 167012 72010 167132 72026
rect 167012 72004 167144 72010
rect 167012 71998 167092 72004
rect 167092 71946 167144 71952
rect 166908 71052 166960 71058
rect 166908 70994 166960 71000
rect 166460 64846 166856 64874
rect 166356 31136 166408 31142
rect 166356 31078 166408 31084
rect 166172 25560 166224 25566
rect 166172 25502 166224 25508
rect 166080 6180 166132 6186
rect 166080 6122 166132 6128
rect 166828 4826 166856 64846
rect 167288 6526 167316 72791
rect 167368 72412 167420 72418
rect 167368 72354 167420 72360
rect 167276 6520 167328 6526
rect 167276 6462 167328 6468
rect 167184 5296 167236 5302
rect 167184 5238 167236 5244
rect 166816 4820 166868 4826
rect 166816 4762 166868 4768
rect 166080 3732 166132 3738
rect 166080 3674 166132 3680
rect 165252 3256 165304 3262
rect 165252 3198 165304 3204
rect 166092 480 166120 3674
rect 167196 480 167224 5238
rect 167380 3398 167408 72354
rect 167460 72344 167512 72350
rect 167460 72286 167512 72292
rect 167472 4078 167500 72286
rect 167552 72140 167604 72146
rect 167552 72082 167604 72088
rect 167460 4072 167512 4078
rect 167460 4014 167512 4020
rect 167564 4010 167592 72082
rect 167552 4004 167604 4010
rect 167552 3946 167604 3952
rect 167656 3806 167684 74462
rect 167748 73642 167776 74616
rect 167736 73636 167788 73642
rect 167736 73578 167788 73584
rect 167840 73098 167868 75140
rect 167736 73092 167788 73098
rect 167736 73034 167788 73040
rect 167828 73092 167880 73098
rect 167828 73034 167880 73040
rect 167748 72758 167776 73034
rect 167736 72752 167788 72758
rect 167736 72694 167788 72700
rect 167932 72418 167960 75140
rect 168024 73137 168052 75140
rect 168116 74798 168144 75140
rect 168104 74792 168156 74798
rect 168104 74734 168156 74740
rect 168104 74656 168156 74662
rect 168208 74633 168236 75140
rect 168300 74905 168328 75140
rect 168286 74896 168342 74905
rect 168286 74831 168342 74840
rect 168104 74598 168156 74604
rect 168194 74624 168250 74633
rect 168116 73154 168144 74598
rect 168194 74559 168250 74568
rect 168392 73914 168420 75140
rect 168380 73908 168432 73914
rect 168380 73850 168432 73856
rect 168010 73128 168066 73137
rect 168116 73126 168236 73154
rect 168010 73063 168066 73072
rect 168104 73024 168156 73030
rect 168104 72966 168156 72972
rect 167920 72412 167972 72418
rect 167920 72354 167972 72360
rect 167736 72208 167788 72214
rect 167736 72150 167788 72156
rect 167644 3800 167696 3806
rect 167644 3742 167696 3748
rect 167748 3738 167776 72150
rect 168116 4146 168144 72966
rect 168104 4140 168156 4146
rect 168104 4082 168156 4088
rect 168208 3942 168236 73126
rect 168484 73030 168512 75140
rect 168576 74526 168604 75140
rect 168564 74520 168616 74526
rect 168564 74462 168616 74468
rect 168472 73024 168524 73030
rect 168472 72966 168524 72972
rect 168562 72720 168618 72729
rect 168562 72655 168618 72664
rect 168288 72276 168340 72282
rect 168288 72218 168340 72224
rect 168196 3936 168248 3942
rect 168196 3878 168248 3884
rect 168300 3874 168328 72218
rect 168576 72185 168604 72655
rect 168562 72176 168618 72185
rect 168562 72111 168618 72120
rect 168668 71602 168696 75140
rect 168656 71596 168708 71602
rect 168656 71538 168708 71544
rect 168760 71466 168788 75140
rect 168748 71460 168800 71466
rect 168748 71402 168800 71408
rect 168852 71398 168880 75140
rect 168944 71534 168972 75140
rect 169036 71670 169064 75140
rect 169128 73817 169156 75140
rect 169114 73808 169170 73817
rect 169114 73743 169170 73752
rect 169220 73681 169248 75140
rect 169206 73672 169262 73681
rect 169206 73607 169262 73616
rect 169312 73545 169340 75140
rect 169404 74769 169432 75140
rect 169390 74760 169446 74769
rect 169390 74695 169446 74704
rect 169392 74656 169444 74662
rect 169392 74598 169444 74604
rect 169404 73817 169432 74598
rect 169496 73953 169524 75140
rect 169588 74769 169616 75140
rect 169574 74760 169630 74769
rect 169574 74695 169630 74704
rect 169482 73944 169538 73953
rect 169482 73879 169538 73888
rect 169390 73808 169446 73817
rect 169390 73743 169446 73752
rect 169298 73536 169354 73545
rect 169680 73506 169708 75140
rect 169772 74934 169800 75140
rect 169760 74928 169812 74934
rect 169760 74870 169812 74876
rect 169298 73471 169354 73480
rect 169668 73500 169720 73506
rect 169668 73442 169720 73448
rect 169864 73438 169892 75140
rect 169956 73710 169984 75140
rect 170048 74322 170076 75140
rect 170036 74316 170088 74322
rect 170036 74258 170088 74264
rect 170140 73778 170168 75140
rect 170128 73772 170180 73778
rect 170128 73714 170180 73720
rect 169944 73704 169996 73710
rect 169944 73646 169996 73652
rect 169852 73432 169904 73438
rect 169852 73374 169904 73380
rect 169024 71664 169076 71670
rect 169024 71606 169076 71612
rect 168932 71528 168984 71534
rect 168932 71470 168984 71476
rect 168840 71392 168892 71398
rect 168840 71334 168892 71340
rect 170232 45558 170260 75140
rect 170220 45552 170272 45558
rect 170220 45494 170272 45500
rect 170324 22710 170352 75140
rect 170416 75002 170444 75210
rect 170496 75200 170548 75206
rect 170496 75142 170548 75148
rect 170404 74996 170456 75002
rect 170404 74938 170456 74944
rect 170404 74724 170456 74730
rect 170404 74666 170456 74672
rect 170416 74594 170444 74666
rect 170508 74594 170536 75142
rect 170588 75132 170640 75138
rect 170588 75074 170640 75080
rect 170404 74588 170456 74594
rect 170404 74530 170456 74536
rect 170496 74588 170548 74594
rect 170496 74530 170548 74536
rect 170600 72554 170628 75074
rect 170692 74866 170720 75618
rect 172244 75336 172296 75342
rect 172244 75278 172296 75284
rect 170864 75064 170916 75070
rect 170864 75006 170916 75012
rect 170772 74928 170824 74934
rect 170772 74870 170824 74876
rect 170680 74860 170732 74866
rect 170680 74802 170732 74808
rect 170784 74746 170812 74870
rect 170692 74718 170812 74746
rect 170692 74662 170720 74718
rect 170680 74656 170732 74662
rect 170680 74598 170732 74604
rect 170876 74089 170904 75006
rect 172256 74866 172284 75278
rect 172794 75168 172850 75177
rect 172794 75103 172850 75112
rect 172610 74896 172666 74905
rect 172244 74860 172296 74866
rect 172610 74831 172666 74840
rect 172244 74802 172296 74808
rect 172152 74792 172204 74798
rect 172152 74734 172204 74740
rect 172334 74760 172390 74769
rect 172060 74724 172112 74730
rect 172060 74666 172112 74672
rect 170862 74080 170918 74089
rect 170862 74015 170918 74024
rect 172072 73574 172100 74666
rect 172164 73642 172192 74734
rect 172334 74695 172390 74704
rect 172348 73817 172376 74695
rect 172624 74633 172652 74831
rect 172808 74633 172836 75103
rect 172610 74624 172666 74633
rect 172610 74559 172666 74568
rect 172794 74624 172850 74633
rect 172794 74559 172850 74568
rect 172334 73808 172390 73817
rect 172334 73743 172390 73752
rect 172152 73636 172204 73642
rect 172152 73578 172204 73584
rect 172060 73568 172112 73574
rect 172060 73510 172112 73516
rect 172888 73160 172940 73166
rect 172888 73102 172940 73108
rect 170588 72548 170640 72554
rect 170588 72490 170640 72496
rect 172900 72457 172928 73102
rect 172886 72448 172942 72457
rect 172886 72383 172942 72392
rect 175292 33114 175320 122806
rect 175936 109041 175964 136478
rect 176028 117298 176056 136546
rect 176672 119785 176700 226986
rect 176752 213988 176804 213994
rect 176752 213930 176804 213936
rect 176764 126993 176792 213930
rect 188344 205692 188396 205698
rect 188344 205634 188396 205640
rect 185584 165640 185636 165646
rect 185584 165582 185636 165588
rect 176844 136468 176896 136474
rect 176844 136410 176896 136416
rect 176750 126984 176806 126993
rect 176750 126919 176806 126928
rect 176658 119776 176714 119785
rect 176658 119711 176714 119720
rect 176016 117292 176068 117298
rect 176016 117234 176068 117240
rect 176660 117292 176712 117298
rect 176660 117234 176712 117240
rect 176672 110401 176700 117234
rect 176856 111761 176884 136410
rect 178132 136400 178184 136406
rect 178132 136342 178184 136348
rect 178040 136128 178092 136134
rect 178040 136070 178092 136076
rect 177304 134768 177356 134774
rect 177304 134710 177356 134716
rect 177316 118590 177344 134710
rect 178052 125497 178080 136070
rect 178038 125488 178094 125497
rect 178038 125423 178094 125432
rect 178144 122505 178172 136342
rect 178592 136332 178644 136338
rect 178592 136274 178644 136280
rect 178408 136264 178460 136270
rect 178408 136206 178460 136212
rect 178316 134700 178368 134706
rect 178316 134642 178368 134648
rect 178130 122496 178186 122505
rect 178130 122431 178186 122440
rect 177304 118584 177356 118590
rect 177304 118526 177356 118532
rect 178224 118584 178276 118590
rect 178224 118526 178276 118532
rect 176842 111752 176898 111761
rect 176842 111687 176898 111696
rect 176658 110392 176714 110401
rect 176658 110327 176714 110336
rect 175922 109032 175978 109041
rect 175922 108967 175978 108976
rect 178236 107545 178264 118526
rect 178328 115297 178356 134642
rect 178420 121281 178448 136206
rect 178500 136060 178552 136066
rect 178500 136002 178552 136008
rect 178512 124137 178540 136002
rect 178498 124128 178554 124137
rect 178498 124063 178554 124072
rect 178406 121272 178462 121281
rect 178406 121207 178462 121216
rect 178604 118289 178632 136274
rect 178776 136196 178828 136202
rect 178776 136138 178828 136144
rect 178684 134632 178736 134638
rect 178684 134574 178736 134580
rect 178590 118280 178646 118289
rect 178590 118215 178646 118224
rect 178314 115288 178370 115297
rect 178314 115223 178370 115232
rect 178696 113121 178724 134574
rect 178788 116793 178816 136138
rect 178866 131200 178922 131209
rect 178866 131135 178922 131144
rect 178774 116784 178830 116793
rect 178774 116719 178830 116728
rect 178682 113112 178738 113121
rect 178682 113047 178738 113056
rect 178222 107536 178278 107545
rect 178222 107471 178278 107480
rect 178040 106276 178092 106282
rect 178040 106218 178092 106224
rect 178052 106049 178080 106218
rect 178038 106040 178094 106049
rect 178038 105975 178094 105984
rect 178040 104848 178092 104854
rect 178040 104790 178092 104796
rect 178052 104553 178080 104790
rect 178038 104544 178094 104553
rect 178038 104479 178094 104488
rect 178040 103488 178092 103494
rect 178040 103430 178092 103436
rect 178052 103057 178080 103430
rect 178038 103048 178094 103057
rect 178038 102983 178094 102992
rect 178040 102128 178092 102134
rect 178040 102070 178092 102076
rect 178052 101697 178080 102070
rect 178038 101688 178094 101697
rect 178038 101623 178094 101632
rect 178040 100700 178092 100706
rect 178040 100642 178092 100648
rect 178052 100201 178080 100642
rect 178038 100192 178094 100201
rect 178038 100127 178094 100136
rect 175924 99408 175976 99414
rect 175924 99350 175976 99356
rect 175936 75750 175964 99350
rect 178040 99340 178092 99346
rect 178040 99282 178092 99288
rect 178052 98841 178080 99282
rect 178038 98832 178094 98841
rect 178038 98767 178094 98776
rect 178040 97980 178092 97986
rect 178040 97922 178092 97928
rect 178052 97345 178080 97922
rect 178038 97336 178094 97345
rect 178038 97271 178094 97280
rect 178040 95192 178092 95198
rect 178038 95160 178040 95169
rect 178092 95160 178094 95169
rect 178038 95095 178094 95104
rect 178040 93832 178092 93838
rect 178038 93800 178040 93809
rect 178092 93800 178094 93809
rect 178038 93735 178094 93744
rect 178040 92472 178092 92478
rect 178040 92414 178092 92420
rect 178052 92313 178080 92414
rect 178038 92304 178094 92313
rect 178038 92239 178094 92248
rect 178040 91044 178092 91050
rect 178040 90986 178092 90992
rect 178052 90953 178080 90986
rect 178038 90944 178094 90953
rect 178038 90879 178094 90888
rect 178040 89684 178092 89690
rect 178040 89626 178092 89632
rect 178052 89457 178080 89626
rect 178038 89448 178094 89457
rect 178038 89383 178094 89392
rect 178040 88324 178092 88330
rect 178040 88266 178092 88272
rect 178052 88097 178080 88266
rect 178038 88088 178094 88097
rect 178038 88023 178094 88032
rect 178040 86964 178092 86970
rect 178040 86906 178092 86912
rect 178052 86601 178080 86906
rect 178038 86592 178094 86601
rect 178038 86527 178094 86536
rect 178040 85536 178092 85542
rect 178040 85478 178092 85484
rect 178052 85105 178080 85478
rect 178038 85096 178094 85105
rect 178038 85031 178094 85040
rect 178040 84176 178092 84182
rect 178040 84118 178092 84124
rect 178052 83745 178080 84118
rect 178038 83736 178094 83745
rect 178038 83671 178094 83680
rect 178040 82816 178092 82822
rect 178040 82758 178092 82764
rect 178052 82249 178080 82758
rect 178038 82240 178094 82249
rect 178038 82175 178094 82184
rect 178682 78704 178738 78713
rect 178682 78639 178738 78648
rect 178038 76664 178094 76673
rect 178038 76599 178094 76608
rect 178052 75954 178080 76599
rect 178040 75948 178092 75954
rect 178040 75890 178092 75896
rect 175924 75744 175976 75750
rect 175924 75686 175976 75692
rect 175372 75200 175424 75206
rect 175372 75142 175424 75148
rect 175384 74526 175412 75142
rect 175372 74520 175424 74526
rect 175372 74462 175424 74468
rect 178696 46918 178724 78639
rect 178880 72078 178908 131135
rect 184204 125656 184256 125662
rect 184204 125598 184256 125604
rect 179236 85604 179288 85610
rect 179236 85546 179288 85552
rect 179248 80889 179276 85546
rect 184216 82822 184244 125598
rect 185596 84182 185624 165582
rect 188356 85542 188384 205634
rect 207032 198014 207060 230588
rect 236012 230574 236578 230602
rect 207020 198008 207072 198014
rect 207020 197950 207072 197956
rect 236012 196654 236040 230574
rect 266556 228478 266584 230588
rect 266544 228472 266596 228478
rect 266544 228414 266596 228420
rect 236644 228404 236696 228410
rect 236644 228346 236696 228352
rect 236656 196722 236684 228346
rect 296732 199442 296760 230588
rect 327092 228478 327120 230588
rect 356072 230574 356546 230602
rect 297364 228472 297416 228478
rect 297364 228414 297416 228420
rect 327080 228472 327132 228478
rect 327080 228414 327132 228420
rect 296720 199436 296772 199442
rect 296720 199378 296772 199384
rect 236644 196716 236696 196722
rect 236644 196658 236696 196664
rect 236000 196648 236052 196654
rect 236000 196590 236052 196596
rect 297376 195906 297404 228414
rect 355324 197396 355376 197402
rect 355324 197338 355376 197344
rect 297364 195900 297416 195906
rect 297364 195842 297416 195848
rect 217324 193860 217376 193866
rect 217324 193802 217376 193808
rect 188344 85536 188396 85542
rect 188344 85478 188396 85484
rect 185584 84176 185636 84182
rect 185584 84118 185636 84124
rect 184204 82816 184256 82822
rect 184204 82758 184256 82764
rect 179234 80880 179290 80889
rect 179234 80815 179290 80824
rect 195980 75064 196032 75070
rect 195980 75006 196032 75012
rect 178868 72072 178920 72078
rect 178868 72014 178920 72020
rect 178684 46912 178736 46918
rect 178684 46854 178736 46860
rect 175280 33108 175332 33114
rect 175280 33050 175332 33056
rect 176660 32972 176712 32978
rect 176660 32914 176712 32920
rect 173898 32736 173954 32745
rect 173898 32671 173954 32680
rect 172518 25664 172574 25673
rect 172518 25599 172574 25608
rect 170312 22704 170364 22710
rect 170312 22646 170364 22652
rect 172532 16574 172560 25599
rect 172532 16546 172744 16574
rect 169024 12300 169076 12306
rect 169024 12242 169076 12248
rect 168288 3868 168340 3874
rect 168288 3810 168340 3816
rect 167736 3732 167788 3738
rect 167736 3674 167788 3680
rect 169036 3670 169064 12242
rect 170312 10872 170364 10878
rect 170312 10814 170364 10820
rect 169666 8120 169722 8129
rect 169666 8055 169722 8064
rect 168380 3664 168432 3670
rect 168380 3606 168432 3612
rect 169024 3664 169076 3670
rect 169024 3606 169076 3612
rect 167368 3392 167420 3398
rect 167368 3334 167420 3340
rect 168392 480 168420 3606
rect 169680 3330 169708 8055
rect 169576 3324 169628 3330
rect 169576 3266 169628 3272
rect 169668 3324 169720 3330
rect 169668 3266 169720 3272
rect 169588 480 169616 3266
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 10814
rect 171968 9648 172020 9654
rect 171968 9590 172020 9596
rect 171980 480 172008 9590
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 32671
rect 176672 11694 176700 32914
rect 180800 32904 180852 32910
rect 180800 32846 180852 32852
rect 179420 26240 179472 26246
rect 179420 26182 179472 26188
rect 176752 25492 176804 25498
rect 176752 25434 176804 25440
rect 176660 11688 176712 11694
rect 176660 11630 176712 11636
rect 176764 6914 176792 25434
rect 179432 16574 179460 26182
rect 180812 16574 180840 32846
rect 184940 32836 184992 32842
rect 184940 32778 184992 32784
rect 183560 26172 183612 26178
rect 183560 26114 183612 26120
rect 183572 16574 183600 26114
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 183572 16546 183784 16574
rect 177856 11688 177908 11694
rect 177856 11630 177908 11636
rect 176672 6886 176792 6914
rect 175464 3324 175516 3330
rect 175464 3266 175516 3272
rect 175476 480 175504 3266
rect 176672 480 176700 6886
rect 177868 480 177896 11630
rect 179052 9580 179104 9586
rect 179052 9522 179104 9528
rect 179064 480 179092 9522
rect 180260 480 180288 16546
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 182548 3256 182600 3262
rect 182548 3198 182600 3204
rect 182560 480 182588 3198
rect 183756 480 183784 16546
rect 184952 480 184980 32778
rect 194600 32768 194652 32774
rect 194600 32710 194652 32716
rect 187698 32600 187754 32609
rect 187698 32535 187754 32544
rect 186320 27532 186372 27538
rect 186320 27474 186372 27480
rect 186332 16574 186360 27474
rect 187712 16574 187740 32535
rect 191838 32464 191894 32473
rect 191838 32399 191894 32408
rect 190458 27160 190514 27169
rect 190458 27095 190514 27104
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 186136 9512 186188 9518
rect 186136 9454 186188 9460
rect 186148 480 186176 9454
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 181414 -960 181526 326
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 189724 4140 189776 4146
rect 189724 4082 189776 4088
rect 189736 480 189764 4082
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190472 354 190500 27095
rect 191852 16574 191880 32399
rect 193220 27600 193272 27606
rect 193220 27542 193272 27548
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 3330 193260 27542
rect 194612 16574 194640 32710
rect 195992 16574 196020 75006
rect 207020 73228 207072 73234
rect 207020 73170 207072 73176
rect 198740 32700 198792 32706
rect 198740 32642 198792 32648
rect 197360 27464 197412 27470
rect 197360 27406 197412 27412
rect 197372 16574 197400 27406
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 193310 4720 193366 4729
rect 193310 4655 193366 4664
rect 193220 3324 193272 3330
rect 193220 3266 193272 3272
rect 193324 2394 193352 4655
rect 194416 3324 194468 3330
rect 194416 3266 194468 3272
rect 193232 2366 193352 2394
rect 193232 480 193260 2366
rect 194428 480 194456 3266
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 32642
rect 205640 32632 205692 32638
rect 205640 32574 205692 32580
rect 201500 27328 201552 27334
rect 201500 27270 201552 27276
rect 200304 10804 200356 10810
rect 200304 10746 200356 10752
rect 200316 480 200344 10746
rect 201512 480 201540 27270
rect 204260 27260 204312 27266
rect 204260 27202 204312 27208
rect 204272 16574 204300 27202
rect 205652 16574 205680 32574
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 203432 10736 203484 10742
rect 203432 10678 203484 10684
rect 202696 5228 202748 5234
rect 202696 5170 202748 5176
rect 202708 480 202736 5170
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 10678
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 73170
rect 217336 72418 217364 193802
rect 355336 189786 355364 197338
rect 356072 195974 356100 230574
rect 380176 228478 380204 231095
rect 366364 228472 366416 228478
rect 366364 228414 366416 228420
rect 380164 228472 380216 228478
rect 380164 228414 380216 228420
rect 364984 205760 365036 205766
rect 364984 205702 365036 205708
rect 362960 201544 363012 201550
rect 362960 201486 363012 201492
rect 362224 198076 362276 198082
rect 362224 198018 362276 198024
rect 356060 195968 356112 195974
rect 356060 195910 356112 195916
rect 341524 189780 341576 189786
rect 341524 189722 341576 189728
rect 355324 189780 355376 189786
rect 355324 189722 355376 189728
rect 341536 179450 341564 189722
rect 362236 189106 362264 198018
rect 362972 197402 363000 201486
rect 364996 198082 365024 205702
rect 366376 201550 366404 228414
rect 386524 228410 386552 230588
rect 390836 230512 390888 230518
rect 390836 230454 390888 230460
rect 386512 228404 386564 228410
rect 386512 228346 386564 228352
rect 387064 227792 387116 227798
rect 387064 227734 387116 227740
rect 384948 226296 385000 226302
rect 384948 226238 385000 226244
rect 384960 223650 384988 226238
rect 384948 223644 385000 223650
rect 384948 223586 385000 223592
rect 380900 223576 380952 223582
rect 380900 223518 380952 223524
rect 380912 221474 380940 223518
rect 372620 221468 372672 221474
rect 372620 221410 372672 221416
rect 380900 221468 380952 221474
rect 380900 221410 380952 221416
rect 372632 220454 372660 221410
rect 369860 220448 369912 220454
rect 369860 220390 369912 220396
rect 372620 220448 372672 220454
rect 372620 220390 372672 220396
rect 369872 216714 369900 220390
rect 387076 218754 387104 227734
rect 390848 226370 390876 230454
rect 392596 227798 392624 232319
rect 396552 232150 396580 238682
rect 394700 232144 394752 232150
rect 394700 232086 394752 232092
rect 396540 232144 396592 232150
rect 396540 232086 396592 232092
rect 394712 230518 394740 232086
rect 394700 230512 394752 230518
rect 394700 230454 394752 230460
rect 392584 227792 392636 227798
rect 392584 227734 392636 227740
rect 390836 226364 390888 226370
rect 390836 226306 390888 226312
rect 379520 218748 379572 218754
rect 379520 218690 379572 218696
rect 387064 218748 387116 218754
rect 387064 218690 387116 218696
rect 379532 216730 379560 218690
rect 369860 216708 369912 216714
rect 369860 216650 369912 216656
rect 379440 216702 379560 216730
rect 366456 216640 366508 216646
rect 366456 216582 366508 216588
rect 366468 205766 366496 216582
rect 379440 211954 379468 216702
rect 375288 211948 375340 211954
rect 375288 211890 375340 211896
rect 379428 211948 379480 211954
rect 379428 211890 379480 211896
rect 375300 209846 375328 211890
rect 371148 209840 371200 209846
rect 371148 209782 371200 209788
rect 375288 209840 375340 209846
rect 375288 209782 375340 209788
rect 366456 205760 366508 205766
rect 366456 205702 366508 205708
rect 371160 204814 371188 209782
rect 382924 209092 382976 209098
rect 382924 209034 382976 209040
rect 367744 204808 367796 204814
rect 367744 204750 367796 204756
rect 371148 204808 371200 204814
rect 371148 204750 371200 204756
rect 366364 201544 366416 201550
rect 366364 201486 366416 201492
rect 364984 198076 365036 198082
rect 364984 198018 365036 198024
rect 362960 197396 363012 197402
rect 362960 197338 363012 197344
rect 359464 189100 359516 189106
rect 359464 189042 359516 189048
rect 362224 189100 362276 189106
rect 362224 189042 362276 189048
rect 336556 179444 336608 179450
rect 336556 179386 336608 179392
rect 341524 179444 341576 179450
rect 341524 179386 341576 179392
rect 336568 174690 336596 179386
rect 329104 174684 329156 174690
rect 329104 174626 329156 174632
rect 336556 174684 336608 174690
rect 336556 174626 336608 174632
rect 329116 163538 329144 174626
rect 359372 166320 359424 166326
rect 359372 166262 359424 166268
rect 314660 163532 314712 163538
rect 314660 163474 314712 163480
rect 329104 163532 329156 163538
rect 329104 163474 329156 163480
rect 314672 156602 314700 163474
rect 359384 162178 359412 166262
rect 338764 162172 338816 162178
rect 338764 162114 338816 162120
rect 359372 162172 359424 162178
rect 359372 162114 359424 162120
rect 309784 156596 309836 156602
rect 309784 156538 309836 156544
rect 314660 156596 314712 156602
rect 314660 156538 314712 156544
rect 309796 149122 309824 156538
rect 307668 149116 307720 149122
rect 307668 149058 307720 149064
rect 309784 149116 309836 149122
rect 309784 149058 309836 149064
rect 307680 143614 307708 149058
rect 303620 143608 303672 143614
rect 303620 143550 303672 143556
rect 307668 143608 307720 143614
rect 307668 143550 307720 143556
rect 303632 138106 303660 143550
rect 300860 138100 300912 138106
rect 300860 138042 300912 138048
rect 303620 138100 303672 138106
rect 303620 138042 303672 138048
rect 300872 136066 300900 138042
rect 295340 136060 295392 136066
rect 295340 136002 295392 136008
rect 300860 136060 300912 136066
rect 300860 136002 300912 136008
rect 295352 134570 295380 136002
rect 295340 134564 295392 134570
rect 295340 134506 295392 134512
rect 333980 112464 334032 112470
rect 333980 112406 334032 112412
rect 333992 111110 334020 112406
rect 324320 111104 324372 111110
rect 324320 111046 324372 111052
rect 333980 111104 334032 111110
rect 333980 111046 334032 111052
rect 324332 107658 324360 111046
rect 324240 107630 324360 107658
rect 324240 104854 324268 107630
rect 324228 104848 324280 104854
rect 324228 104790 324280 104796
rect 338776 91798 338804 162114
rect 359476 155990 359504 189042
rect 367756 187746 367784 204750
rect 382936 198762 382964 209034
rect 377404 198756 377456 198762
rect 377404 198698 377456 198704
rect 382924 198756 382976 198762
rect 382924 198698 382976 198704
rect 366364 187740 366416 187746
rect 366364 187682 366416 187688
rect 367744 187740 367796 187746
rect 367744 187682 367796 187688
rect 364984 174684 365036 174690
rect 364984 174626 365036 174632
rect 362224 168564 362276 168570
rect 362224 168506 362276 168512
rect 362236 160138 362264 168506
rect 364996 166326 365024 174626
rect 366376 168570 366404 187682
rect 377416 184210 377444 198698
rect 371884 184204 371936 184210
rect 371884 184146 371936 184152
rect 377404 184204 377456 184210
rect 377404 184146 377456 184152
rect 371896 176730 371924 184146
rect 368480 176724 368532 176730
rect 368480 176666 368532 176672
rect 371884 176724 371936 176730
rect 371884 176666 371936 176672
rect 368492 174690 368520 176666
rect 368480 174684 368532 174690
rect 368480 174626 368532 174632
rect 366364 168564 366416 168570
rect 366364 168506 366416 168512
rect 364984 166320 365036 166326
rect 364984 166262 365036 166268
rect 360200 160132 360252 160138
rect 360200 160074 360252 160080
rect 362224 160132 362276 160138
rect 362224 160074 362276 160080
rect 359464 155984 359516 155990
rect 359464 155926 359516 155932
rect 356704 155916 356756 155922
rect 356704 155858 356756 155864
rect 351920 145580 351972 145586
rect 351920 145522 351972 145528
rect 351932 143614 351960 145522
rect 351920 143608 351972 143614
rect 351920 143550 351972 143556
rect 347044 143540 347096 143546
rect 347044 143482 347096 143488
rect 347056 121514 347084 143482
rect 356716 124234 356744 155858
rect 360212 154222 360240 160074
rect 357992 154216 358044 154222
rect 357992 154158 358044 154164
rect 360200 154216 360252 154222
rect 360200 154158 360252 154164
rect 358004 145586 358032 154158
rect 357992 145580 358044 145586
rect 357992 145522 358044 145528
rect 350724 124228 350776 124234
rect 350724 124170 350776 124176
rect 356704 124228 356756 124234
rect 356704 124170 356756 124176
rect 350736 121514 350764 124170
rect 345756 121508 345808 121514
rect 345756 121450 345808 121456
rect 347044 121508 347096 121514
rect 347044 121450 347096 121456
rect 347872 121508 347924 121514
rect 347872 121450 347924 121456
rect 350724 121508 350776 121514
rect 350724 121450 350776 121456
rect 345768 118250 345796 121450
rect 342260 118244 342312 118250
rect 342260 118186 342312 118192
rect 345756 118244 345808 118250
rect 345756 118186 345808 118192
rect 342272 114578 342300 118186
rect 347884 117978 347912 121450
rect 343640 117972 343692 117978
rect 343640 117914 343692 117920
rect 347872 117972 347924 117978
rect 347872 117914 347924 117920
rect 342260 114572 342312 114578
rect 342260 114514 342312 114520
rect 340420 114504 340472 114510
rect 340420 114446 340472 114452
rect 340432 112470 340460 114446
rect 343652 113762 343680 117914
rect 341524 113756 341576 113762
rect 341524 113698 341576 113704
rect 343640 113756 343692 113762
rect 343640 113698 343692 113704
rect 340420 112464 340472 112470
rect 340420 112406 340472 112412
rect 341536 106282 341564 113698
rect 341524 106276 341576 106282
rect 341524 106218 341576 106224
rect 320824 91792 320876 91798
rect 320824 91734 320876 91740
rect 338764 91792 338816 91798
rect 338764 91734 338816 91740
rect 320836 84862 320864 91734
rect 307760 84856 307812 84862
rect 307760 84798 307812 84804
rect 320824 84856 320876 84862
rect 320824 84798 320876 84804
rect 307772 77994 307800 84798
rect 299388 77988 299440 77994
rect 299388 77930 299440 77936
rect 307760 77988 307812 77994
rect 307760 77930 307812 77936
rect 299400 75206 299428 77930
rect 299388 75200 299440 75206
rect 299388 75142 299440 75148
rect 259460 75132 259512 75138
rect 259460 75074 259512 75080
rect 249800 74248 249852 74254
rect 249800 74190 249852 74196
rect 217324 72412 217376 72418
rect 217324 72354 217376 72360
rect 226340 40724 226392 40730
rect 226340 40666 226392 40672
rect 212540 34468 212592 34474
rect 212540 34410 212592 34416
rect 209778 34096 209834 34105
rect 209778 34031 209834 34040
rect 208400 27396 208452 27402
rect 208400 27338 208452 27344
rect 208412 16574 208440 27338
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209792 480 209820 34031
rect 211160 28144 211212 28150
rect 211160 28086 211212 28092
rect 211172 16574 211200 28086
rect 212552 16574 212580 34410
rect 216680 34400 216732 34406
rect 216680 34342 216732 34348
rect 215300 28212 215352 28218
rect 215300 28154 215352 28160
rect 211172 16546 211752 16574
rect 212552 16546 213408 16574
rect 210974 12200 211030 12209
rect 210974 12135 211030 12144
rect 210988 480 211016 12135
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213380 480 213408 16546
rect 214472 12232 214524 12238
rect 214472 12174 214524 12180
rect 214484 480 214512 12174
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 28154
rect 216692 16574 216720 34342
rect 219440 34332 219492 34338
rect 219440 34274 219492 34280
rect 218060 27192 218112 27198
rect 218060 27134 218112 27140
rect 216692 16546 216904 16574
rect 216876 480 216904 16546
rect 218072 11694 218100 27134
rect 219452 16574 219480 34274
rect 222200 28076 222252 28082
rect 222200 28018 222252 28024
rect 222212 16574 222240 28018
rect 223578 20224 223634 20233
rect 223578 20159 223634 20168
rect 219452 16546 220032 16574
rect 222212 16546 222792 16574
rect 218152 12164 218204 12170
rect 218152 12106 218204 12112
rect 218060 11688 218112 11694
rect 218060 11630 218112 11636
rect 218164 6914 218192 12106
rect 219256 11688 219308 11694
rect 219256 11630 219308 11636
rect 218072 6886 218192 6914
rect 218072 480 218100 6886
rect 219268 480 219296 11630
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 221096 12096 221148 12102
rect 221096 12038 221148 12044
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 12038
rect 222764 480 222792 16546
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 20159
rect 225142 12880 225198 12889
rect 225142 12815 225198 12824
rect 225156 480 225184 12815
rect 226352 3330 226380 40666
rect 234620 34264 234672 34270
rect 234620 34206 234672 34212
rect 229100 28960 229152 28966
rect 229100 28902 229152 28908
rect 229112 16574 229140 28902
rect 233240 27124 233292 27130
rect 233240 27066 233292 27072
rect 230480 20460 230532 20466
rect 230480 20402 230532 20408
rect 230492 16574 230520 20402
rect 233252 16574 233280 27066
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 233252 16546 233464 16574
rect 228730 6896 228786 6905
rect 228730 6831 228786 6840
rect 226430 6080 226486 6089
rect 226430 6015 226486 6024
rect 226340 3324 226392 3330
rect 226340 3266 226392 3272
rect 226444 3074 226472 6015
rect 227536 3324 227588 3330
rect 227536 3266 227588 3272
rect 226352 3046 226472 3074
rect 226352 480 226380 3046
rect 227548 480 227576 3266
rect 228744 480 228772 6831
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 231860 13456 231912 13462
rect 231860 13398 231912 13404
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 13398
rect 233436 480 233464 16546
rect 234632 480 234660 34206
rect 248420 34196 248472 34202
rect 248420 34138 248472 34144
rect 241518 33960 241574 33969
rect 241518 33895 241574 33904
rect 240140 28824 240192 28830
rect 240140 28766 240192 28772
rect 236000 26104 236052 26110
rect 236000 26046 236052 26052
rect 236012 16574 236040 26046
rect 237380 20392 237432 20398
rect 237380 20334 237432 20340
rect 237392 16574 237420 20334
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 235816 6792 235868 6798
rect 235816 6734 235868 6740
rect 235828 480 235856 6734
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239312 13388 239364 13394
rect 239312 13330 239364 13336
rect 239324 480 239352 13330
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 28766
rect 241532 16574 241560 33895
rect 242900 28892 242952 28898
rect 242900 28834 242952 28840
rect 241532 16546 241744 16574
rect 241716 480 241744 16546
rect 242912 11694 242940 28834
rect 247040 28756 247092 28762
rect 247040 28698 247092 28704
rect 244278 20088 244334 20097
rect 244278 20023 244334 20032
rect 244292 16574 244320 20023
rect 247052 16574 247080 28698
rect 244292 16546 245240 16574
rect 247052 16546 247632 16574
rect 242990 13696 243046 13705
rect 242990 13631 243046 13640
rect 242900 11688 242952 11694
rect 242900 11630 242952 11636
rect 243004 6914 243032 13631
rect 244096 11688 244148 11694
rect 244096 11630 244148 11636
rect 242912 6886 243032 6914
rect 242912 480 242940 6886
rect 244108 480 244136 11630
rect 245212 480 245240 16546
rect 246394 6760 246450 6769
rect 246394 6695 246450 6704
rect 246408 480 246436 6695
rect 247604 480 247632 16546
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 354 248460 34138
rect 249812 16574 249840 74190
rect 255320 34128 255372 34134
rect 255320 34070 255372 34076
rect 251180 28620 251232 28626
rect 251180 28562 251232 28568
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 480 251220 28562
rect 253940 24812 253992 24818
rect 253940 24754 253992 24760
rect 251272 19100 251324 19106
rect 251272 19042 251324 19048
rect 251284 16574 251312 19042
rect 253952 16574 253980 24754
rect 255332 16574 255360 34070
rect 258080 28688 258132 28694
rect 258080 28630 258132 28636
rect 258092 16574 258120 28630
rect 251284 16546 252416 16574
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 258092 16546 258304 16574
rect 252388 480 252416 16546
rect 253480 14884 253532 14890
rect 253480 14826 253532 14832
rect 253492 480 253520 14826
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 256700 14816 256752 14822
rect 256700 14758 256752 14764
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 14758
rect 258276 480 258304 16546
rect 259472 11694 259500 75074
rect 302240 74996 302292 75002
rect 302240 74938 302292 74944
rect 284300 74180 284352 74186
rect 284300 74122 284352 74128
rect 269120 34060 269172 34066
rect 269120 34002 269172 34008
rect 262218 33824 262274 33833
rect 262218 33759 262274 33768
rect 260840 26036 260892 26042
rect 260840 25978 260892 25984
rect 259552 20324 259604 20330
rect 259552 20266 259604 20272
rect 259460 11688 259512 11694
rect 259460 11630 259512 11636
rect 259564 6914 259592 20266
rect 260852 16574 260880 25978
rect 262232 16574 262260 33759
rect 266360 32564 266412 32570
rect 266360 32506 266412 32512
rect 264980 28552 265032 28558
rect 264980 28494 265032 28500
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 260656 11688 260708 11694
rect 260656 11630 260708 11636
rect 259472 6886 259592 6914
rect 259472 480 259500 6886
rect 260668 480 260696 11630
rect 261772 480 261800 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264150 15192 264206 15201
rect 264150 15127 264206 15136
rect 264164 480 264192 15127
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 28494
rect 266372 16574 266400 32506
rect 269132 16574 269160 34002
rect 276020 33992 276072 33998
rect 276020 33934 276072 33940
rect 271880 28484 271932 28490
rect 271880 28426 271932 28432
rect 271892 16574 271920 28426
rect 273260 17672 273312 17678
rect 273260 17614 273312 17620
rect 266372 16546 266584 16574
rect 269132 16546 270080 16574
rect 271892 16546 272472 16574
rect 266556 480 266584 16546
rect 267740 14748 267792 14754
rect 267740 14690 267792 14696
rect 267752 480 267780 14690
rect 268844 7948 268896 7954
rect 268844 7890 268896 7896
rect 268856 480 268884 7890
rect 270052 480 270080 16546
rect 270776 14680 270828 14686
rect 270776 14622 270828 14628
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 354 270816 14622
rect 272444 480 272472 16546
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 17614
rect 274824 16380 274876 16386
rect 274824 16322 274876 16328
rect 274836 480 274864 16322
rect 276032 4146 276060 33934
rect 278778 27024 278834 27033
rect 278778 26959 278834 26968
rect 278792 16574 278820 26959
rect 282920 24744 282972 24750
rect 282920 24686 282972 24692
rect 282932 16574 282960 24686
rect 278792 16546 279096 16574
rect 282932 16546 283144 16574
rect 276112 10668 276164 10674
rect 276112 10610 276164 10616
rect 276020 4140 276072 4146
rect 276020 4082 276072 4088
rect 276124 3482 276152 10610
rect 278318 7984 278374 7993
rect 278318 7919 278374 7928
rect 276756 4140 276808 4146
rect 276756 4082 276808 4088
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276768 354 276796 4082
rect 278332 480 278360 7919
rect 277094 354 277206 480
rect 276768 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280710 13560 280766 13569
rect 280710 13495 280766 13504
rect 280724 480 280752 13495
rect 281906 7848 281962 7857
rect 281906 7783 281962 7792
rect 281920 480 281948 7783
rect 283116 480 283144 16546
rect 284312 4146 284340 74122
rect 298098 35320 298154 35329
rect 298098 35255 298154 35264
rect 284392 33924 284444 33930
rect 284392 33866 284444 33872
rect 284300 4140 284352 4146
rect 284300 4082 284352 4088
rect 284404 3482 284432 33866
rect 291200 33856 291252 33862
rect 291200 33798 291252 33804
rect 291212 16574 291240 33798
rect 292580 25968 292632 25974
rect 292580 25910 292632 25916
rect 291212 16546 291424 16574
rect 287336 16312 287388 16318
rect 287336 16254 287388 16260
rect 286600 6724 286652 6730
rect 286600 6666 286652 6672
rect 285036 4140 285088 4146
rect 285036 4082 285088 4088
rect 284312 3454 284432 3482
rect 284312 480 284340 3454
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285048 354 285076 4082
rect 286612 480 286640 6666
rect 285374 354 285486 480
rect 285048 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16254
rect 288992 16244 289044 16250
rect 288992 16186 289044 16192
rect 289004 480 289032 16186
rect 290188 7880 290240 7886
rect 290188 7822 290240 7828
rect 290200 480 290228 7822
rect 291396 480 291424 16546
rect 292592 4146 292620 25910
rect 295614 16280 295670 16289
rect 295614 16215 295670 16224
rect 292672 16176 292724 16182
rect 292672 16118 292724 16124
rect 292580 4140 292632 4146
rect 292580 4082 292632 4088
rect 292684 3482 292712 16118
rect 294880 10600 294932 10606
rect 294880 10542 294932 10548
rect 293316 4140 293368 4146
rect 293316 4082 293368 4088
rect 292592 3454 292712 3482
rect 292592 480 292620 3454
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293328 354 293356 4082
rect 294892 480 294920 10542
rect 293654 354 293766 480
rect 293328 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16215
rect 297270 15056 297326 15065
rect 297270 14991 297326 15000
rect 297284 480 297312 14991
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298112 354 298140 35255
rect 300860 33788 300912 33794
rect 300860 33730 300912 33736
rect 299480 30252 299532 30258
rect 299480 30194 299532 30200
rect 299492 3330 299520 30194
rect 300872 16574 300900 33730
rect 302252 16574 302280 74938
rect 324320 74928 324372 74934
rect 324320 74870 324372 74876
rect 320180 74112 320232 74118
rect 320180 74054 320232 74060
rect 307760 35896 307812 35902
rect 307760 35838 307812 35844
rect 305000 35148 305052 35154
rect 305000 35090 305052 35096
rect 303620 30184 303672 30190
rect 303620 30126 303672 30132
rect 303632 16574 303660 30126
rect 305012 16574 305040 35090
rect 300872 16546 301544 16574
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 299662 9072 299718 9081
rect 299662 9007 299718 9016
rect 299480 3324 299532 3330
rect 299480 3266 299532 3272
rect 299676 480 299704 9007
rect 300768 3324 300820 3330
rect 300768 3266 300820 3272
rect 300780 480 300808 3266
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303172 480 303200 16546
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 306748 9444 306800 9450
rect 306748 9386 306800 9392
rect 306760 480 306788 9386
rect 307772 3330 307800 35838
rect 311900 35828 311952 35834
rect 311900 35770 311952 35776
rect 307852 30320 307904 30326
rect 307852 30262 307904 30268
rect 307864 16574 307892 30262
rect 311912 16574 311940 35770
rect 318800 35760 318852 35766
rect 318800 35702 318852 35708
rect 314658 29608 314714 29617
rect 314658 29543 314714 29552
rect 312544 19032 312596 19038
rect 312544 18974 312596 18980
rect 307864 16546 307984 16574
rect 311912 16546 312216 16574
rect 307760 3324 307812 3330
rect 307760 3266 307812 3272
rect 307956 480 307984 16546
rect 310244 9376 310296 9382
rect 310244 9318 310296 9324
rect 309048 3324 309100 3330
rect 309048 3266 309100 3272
rect 309060 480 309088 3266
rect 310256 480 310284 9318
rect 311440 9308 311492 9314
rect 311440 9250 311492 9256
rect 311452 480 311480 9250
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 312556 4146 312584 18974
rect 313832 10532 313884 10538
rect 313832 10474 313884 10480
rect 312544 4140 312596 4146
rect 312544 4082 312596 4088
rect 313844 480 313872 10474
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 29543
rect 316038 17640 316094 17649
rect 316038 17575 316094 17584
rect 316052 3330 316080 17575
rect 318812 16574 318840 35702
rect 320192 16574 320220 74054
rect 322940 35692 322992 35698
rect 322940 35634 322992 35640
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 316222 14920 316278 14929
rect 316222 14855 316278 14864
rect 316040 3324 316092 3330
rect 316040 3266 316092 3272
rect 316236 480 316264 14855
rect 318064 10464 318116 10470
rect 318064 10406 318116 10412
rect 317328 3324 317380 3330
rect 317328 3266 317380 3272
rect 317340 480 317368 3266
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 10406
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322112 12028 322164 12034
rect 322112 11970 322164 11976
rect 322124 480 322152 11970
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 35634
rect 324332 3210 324360 74870
rect 374000 74860 374052 74866
rect 374000 74802 374052 74808
rect 338120 74044 338172 74050
rect 338120 73986 338172 73992
rect 326344 58676 326396 58682
rect 326344 58618 326396 58624
rect 325700 35624 325752 35630
rect 325700 35566 325752 35572
rect 324412 13320 324464 13326
rect 324412 13262 324464 13268
rect 324424 3330 324452 13262
rect 325712 6914 325740 35566
rect 326356 16574 326384 58618
rect 336740 35556 336792 35562
rect 336740 35498 336792 35504
rect 332598 35184 332654 35193
rect 332598 35119 332654 35128
rect 329840 20256 329892 20262
rect 329840 20198 329892 20204
rect 327080 17604 327132 17610
rect 327080 17546 327132 17552
rect 327092 16574 327120 17546
rect 329852 16574 329880 20198
rect 326356 16546 326476 16574
rect 327092 16546 328040 16574
rect 329852 16546 330432 16574
rect 325712 6886 326384 6914
rect 324412 3324 324464 3330
rect 324412 3266 324464 3272
rect 325608 3324 325660 3330
rect 325608 3266 325660 3272
rect 324332 3182 324452 3210
rect 324424 480 324452 3182
rect 325620 480 325648 3266
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 6886
rect 326448 3262 326476 16546
rect 326436 3256 326488 3262
rect 326436 3198 326488 3204
rect 328012 480 328040 16546
rect 328736 13252 328788 13258
rect 328736 13194 328788 13200
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 13194
rect 330404 480 330432 16546
rect 331218 10432 331274 10441
rect 331218 10367 331274 10376
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 10367
rect 332612 3330 332640 35119
rect 336752 16574 336780 35498
rect 338132 16574 338160 73986
rect 347780 35488 347832 35494
rect 347780 35430 347832 35436
rect 343640 27056 343692 27062
rect 343640 26998 343692 27004
rect 340880 22092 340932 22098
rect 340880 22034 340932 22040
rect 340892 16574 340920 22034
rect 343652 16574 343680 26998
rect 347792 16574 347820 35430
rect 354680 35420 354732 35426
rect 354680 35362 354732 35368
rect 350538 21448 350594 21457
rect 350538 21383 350594 21392
rect 350552 16574 350580 21383
rect 354692 16574 354720 35362
rect 357440 35352 357492 35358
rect 357440 35294 357492 35300
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 340892 16546 341012 16574
rect 343652 16546 344600 16574
rect 347792 16546 348096 16574
rect 350552 16546 351224 16574
rect 354692 16546 355272 16574
rect 332690 14784 332746 14793
rect 332690 14719 332746 14728
rect 332600 3324 332652 3330
rect 332600 3266 332652 3272
rect 332704 480 332732 14719
rect 334622 10296 334678 10305
rect 334622 10231 334678 10240
rect 333888 3324 333940 3330
rect 333888 3266 333940 3272
rect 333900 480 333928 3266
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 10231
rect 336280 7812 336332 7818
rect 336280 7754 336332 7760
rect 336292 480 336320 7754
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 339868 9240 339920 9246
rect 339868 9182 339920 9188
rect 339880 480 339908 9182
rect 340984 480 341012 16546
rect 342904 11960 342956 11966
rect 342904 11902 342956 11908
rect 342168 9172 342220 9178
rect 342168 9114 342220 9120
rect 342180 480 342208 9114
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 11902
rect 344572 480 344600 16546
rect 346952 16108 347004 16114
rect 346952 16050 347004 16056
rect 345296 11892 345348 11898
rect 345296 11834 345348 11840
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 11834
rect 346964 480 346992 16050
rect 348068 480 348096 16546
rect 349158 16144 349214 16153
rect 349158 16079 349214 16088
rect 349172 3262 349200 16079
rect 349250 12064 349306 12073
rect 349250 11999 349306 12008
rect 349160 3256 349212 3262
rect 349160 3198 349212 3204
rect 349264 480 349292 11999
rect 350448 3256 350500 3262
rect 350448 3198 350500 3204
rect 350460 480 350488 3198
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 353576 16040 353628 16046
rect 353576 15982 353628 15988
rect 352838 11928 352894 11937
rect 352838 11863 352894 11872
rect 352852 480 352880 11863
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 15982
rect 355244 480 355272 16546
rect 356336 11824 356388 11830
rect 356336 11766 356388 11772
rect 356348 480 356376 11766
rect 357452 3262 357480 35294
rect 368480 35284 368532 35290
rect 368480 35226 368532 35232
rect 367098 26888 367154 26897
rect 367098 26823 367154 26832
rect 357532 25900 357584 25906
rect 357532 25842 357584 25848
rect 357440 3256 357492 3262
rect 357440 3198 357492 3204
rect 357544 480 357572 25842
rect 361580 22024 361632 22030
rect 361580 21966 361632 21972
rect 358820 18964 358872 18970
rect 358820 18906 358872 18912
rect 358832 16574 358860 18906
rect 361592 16574 361620 21966
rect 367112 16574 367140 26823
rect 368492 16574 368520 35226
rect 371240 28416 371292 28422
rect 371240 28358 371292 28364
rect 358832 16546 359504 16574
rect 361592 16546 361896 16574
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 358728 3256 358780 3262
rect 358728 3198 358780 3204
rect 358740 480 358768 3198
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 361120 14612 361172 14618
rect 361120 14554 361172 14560
rect 361132 480 361160 14554
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 365718 13424 365774 13433
rect 365718 13359 365774 13368
rect 363512 13184 363564 13190
rect 363512 13126 363564 13132
rect 363524 480 363552 13126
rect 364616 5160 364668 5166
rect 364616 5102 364668 5108
rect 364628 480 364656 5102
rect 365732 3262 365760 13359
rect 365810 11792 365866 11801
rect 365810 11727 365866 11736
rect 365720 3256 365772 3262
rect 365720 3198 365772 3204
rect 365824 480 365852 11727
rect 367008 3256 367060 3262
rect 367008 3198 367060 3204
rect 367020 480 367048 3198
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 370134 13288 370190 13297
rect 370134 13223 370190 13232
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 13223
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 28358
rect 372620 25832 372672 25838
rect 372620 25774 372672 25780
rect 372632 16574 372660 25774
rect 372632 16546 372936 16574
rect 372908 480 372936 16546
rect 374012 3074 374040 74802
rect 396736 74798 396764 378150
rect 396908 364404 396960 364410
rect 396908 364346 396960 364352
rect 396816 324352 396868 324358
rect 396816 324294 396868 324300
rect 396724 74792 396776 74798
rect 396724 74734 396776 74740
rect 396828 74730 396856 324294
rect 396920 137630 396948 364346
rect 397092 311908 397144 311914
rect 397092 311850 397144 311856
rect 397000 271924 397052 271930
rect 397000 271866 397052 271872
rect 396908 137624 396960 137630
rect 396908 137566 396960 137572
rect 396816 74724 396868 74730
rect 396816 74666 396868 74672
rect 397012 74225 397040 271866
rect 397104 137562 397132 311850
rect 397184 258120 397236 258126
rect 397184 258062 397236 258068
rect 397092 137556 397144 137562
rect 397092 137498 397144 137504
rect 397196 137494 397224 258062
rect 397184 137488 397236 137494
rect 397184 137430 397236 137436
rect 396998 74216 397054 74225
rect 396998 74151 397054 74160
rect 390560 73976 390612 73982
rect 390560 73918 390612 73924
rect 382280 36712 382332 36718
rect 382280 36654 382332 36660
rect 374092 30116 374144 30122
rect 374092 30058 374144 30064
rect 374104 3262 374132 30058
rect 375380 28348 375432 28354
rect 375380 28290 375432 28296
rect 375392 16574 375420 28290
rect 376760 18896 376812 18902
rect 376760 18838 376812 18844
rect 376772 16574 376800 18838
rect 380900 18828 380952 18834
rect 380900 18770 380952 18776
rect 380912 16574 380940 18770
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 380912 16546 381216 16574
rect 374092 3256 374144 3262
rect 374092 3198 374144 3204
rect 375288 3256 375340 3262
rect 375288 3198 375340 3204
rect 374012 3046 374132 3074
rect 374104 480 374132 3046
rect 375300 480 375328 3198
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 378416 13116 378468 13122
rect 378416 13058 378468 13064
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 13058
rect 379980 6656 380032 6662
rect 379980 6598 380032 6604
rect 379992 480 380020 6598
rect 381188 480 381216 16546
rect 382292 3262 382320 36654
rect 382372 30048 382424 30054
rect 382372 29990 382424 29996
rect 382280 3256 382332 3262
rect 382280 3198 382332 3204
rect 382384 480 382412 29990
rect 389180 29980 389232 29986
rect 389180 29922 389232 29928
rect 386418 24440 386474 24449
rect 386418 24375 386474 24384
rect 386432 16574 386460 24375
rect 389192 16574 389220 29922
rect 386432 16546 386736 16574
rect 389192 16546 389496 16574
rect 384304 14544 384356 14550
rect 384304 14486 384356 14492
rect 383568 3256 383620 3262
rect 383568 3198 383620 3204
rect 383580 480 383608 3198
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 14486
rect 385958 6624 386014 6633
rect 385958 6559 386014 6568
rect 385972 480 386000 6559
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387798 14648 387854 14657
rect 387798 14583 387854 14592
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 14583
rect 389468 480 389496 16546
rect 390572 3262 390600 73918
rect 397472 73030 397500 703520
rect 410524 700460 410576 700466
rect 410524 700402 410576 700408
rect 409144 700392 409196 700398
rect 409144 700334 409196 700340
rect 407764 700324 407816 700330
rect 407764 700266 407816 700272
rect 406384 616888 406436 616894
rect 406384 616830 406436 616836
rect 397552 599616 397604 599622
rect 397552 599558 397604 599564
rect 397564 209098 397592 599558
rect 405004 563100 405056 563106
rect 405004 563042 405056 563048
rect 403624 510672 403676 510678
rect 403624 510614 403676 510620
rect 400864 456816 400916 456822
rect 400864 456758 400916 456764
rect 399484 444440 399536 444446
rect 399484 444382 399536 444388
rect 397552 209092 397604 209098
rect 397552 209034 397604 209040
rect 399496 187678 399524 444382
rect 399484 187672 399536 187678
rect 399484 187614 399536 187620
rect 400876 92478 400904 456758
rect 403636 93838 403664 510614
rect 405016 95198 405044 563042
rect 406396 97986 406424 616830
rect 407776 100706 407804 700266
rect 409156 102134 409184 700334
rect 410536 103494 410564 700402
rect 412652 137426 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 700466 429884 703520
rect 429844 700460 429896 700466
rect 429844 700402 429896 700408
rect 417424 404388 417476 404394
rect 417424 404330 417476 404336
rect 414664 351960 414716 351966
rect 414664 351902 414716 351908
rect 413284 244316 413336 244322
rect 413284 244258 413336 244264
rect 412640 137420 412692 137426
rect 412640 137362 412692 137368
rect 410524 103488 410576 103494
rect 410524 103430 410576 103436
rect 409144 102128 409196 102134
rect 409144 102070 409196 102076
rect 407764 100700 407816 100706
rect 407764 100642 407816 100648
rect 406384 97980 406436 97986
rect 406384 97922 406436 97928
rect 405004 95192 405056 95198
rect 405004 95134 405056 95140
rect 403624 93832 403676 93838
rect 403624 93774 403676 93780
rect 400864 92472 400916 92478
rect 400864 92414 400916 92420
rect 413296 86970 413324 244258
rect 414676 89690 414704 351902
rect 417436 91050 417464 404330
rect 417424 91044 417476 91050
rect 417424 90986 417476 90992
rect 414664 89684 414716 89690
rect 414664 89626 414716 89632
rect 413284 86964 413336 86970
rect 413284 86906 413336 86912
rect 462332 73914 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 477512 137358 477540 702406
rect 494808 700398 494836 703520
rect 494796 700392 494848 700398
rect 494796 700334 494848 700340
rect 520924 231872 520976 231878
rect 520924 231814 520976 231820
rect 477500 137352 477552 137358
rect 477500 137294 477552 137300
rect 462412 74656 462464 74662
rect 462412 74598 462464 74604
rect 462320 73908 462372 73914
rect 462320 73850 462372 73856
rect 397460 73024 397512 73030
rect 397460 72966 397512 72972
rect 422300 72956 422352 72962
rect 422300 72898 422352 72904
rect 390652 36644 390704 36650
rect 390652 36586 390704 36592
rect 390560 3256 390612 3262
rect 390560 3198 390612 3204
rect 390664 480 390692 36586
rect 397460 36576 397512 36582
rect 397460 36518 397512 36524
rect 394700 20188 394752 20194
rect 394700 20130 394752 20136
rect 394712 16574 394740 20130
rect 397472 16574 397500 36518
rect 414020 25764 414072 25770
rect 414020 25706 414072 25712
rect 407212 24676 407264 24682
rect 407212 24618 407264 24624
rect 398840 20120 398892 20126
rect 398840 20062 398892 20068
rect 394712 16546 395384 16574
rect 397472 16546 397776 16574
rect 393044 9104 393096 9110
rect 393044 9046 393096 9052
rect 391848 3256 391900 3262
rect 391848 3198 391900 3204
rect 391860 480 391888 3198
rect 393056 480 393084 9046
rect 394240 3392 394292 3398
rect 394240 3334 394292 3340
rect 394252 480 394280 3334
rect 395356 480 395384 16546
rect 396540 6588 396592 6594
rect 396540 6530 396592 6536
rect 396552 480 396580 6530
rect 397748 480 397776 16546
rect 398852 3210 398880 20062
rect 406014 16008 406070 16017
rect 406014 15943 406070 15952
rect 402518 14512 402574 14521
rect 402518 14447 402574 14456
rect 398932 10396 398984 10402
rect 398932 10338 398984 10344
rect 398944 3398 398972 10338
rect 401324 4072 401376 4078
rect 401324 4014 401376 4020
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 398852 3182 398972 3210
rect 398944 480 398972 3182
rect 400140 480 400168 3334
rect 401336 480 401364 4014
rect 402532 480 402560 14447
rect 403622 11656 403678 11665
rect 403622 11591 403678 11600
rect 403636 480 403664 11591
rect 404818 5536 404874 5545
rect 404818 5471 404874 5480
rect 404832 480 404860 5471
rect 406028 480 406056 15943
rect 407224 480 407252 24618
rect 412640 20052 412692 20058
rect 412640 19994 412692 20000
rect 410800 9036 410852 9042
rect 410800 8978 410852 8984
rect 408408 4004 408460 4010
rect 408408 3946 408460 3952
rect 408420 480 408448 3946
rect 409604 3936 409656 3942
rect 409604 3878 409656 3884
rect 409616 480 409644 3878
rect 410812 480 410840 8978
rect 411904 8968 411956 8974
rect 411904 8910 411956 8916
rect 411916 480 411944 8910
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 19994
rect 414032 16574 414060 25706
rect 420918 17504 420974 17513
rect 420918 17439 420974 17448
rect 414032 16546 414336 16574
rect 414308 480 414336 16546
rect 415492 15972 415544 15978
rect 415492 15914 415544 15920
rect 415400 3868 415452 3874
rect 415400 3810 415452 3816
rect 415412 1986 415440 3810
rect 415504 3398 415532 15914
rect 420182 15872 420238 15881
rect 420182 15807 420238 15816
rect 418526 13152 418582 13161
rect 418526 13087 418582 13096
rect 417884 7744 417936 7750
rect 417884 7686 417936 7692
rect 415492 3392 415544 3398
rect 415492 3334 415544 3340
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 415412 1958 415532 1986
rect 415504 480 415532 1958
rect 416700 480 416728 3334
rect 417896 480 417924 7686
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418540 354 418568 13087
rect 420196 480 420224 15807
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 17439
rect 422312 16574 422340 72898
rect 443000 72888 443052 72894
rect 443000 72830 443052 72836
rect 431960 29912 432012 29918
rect 431960 29854 432012 29860
rect 423680 26988 423732 26994
rect 423680 26930 423732 26936
rect 422312 16546 422616 16574
rect 422588 480 422616 16546
rect 423692 1290 423720 26930
rect 425060 21956 425112 21962
rect 425060 21898 425112 21904
rect 423770 17368 423826 17377
rect 423770 17303 423826 17312
rect 423680 1284 423732 1290
rect 423680 1226 423732 1232
rect 423784 480 423812 17303
rect 425072 16574 425100 21898
rect 430580 21888 430632 21894
rect 430580 21830 430632 21836
rect 427820 17536 427872 17542
rect 427820 17478 427872 17484
rect 427832 16574 427860 17478
rect 430592 16574 430620 21830
rect 425072 16546 425744 16574
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 424968 1284 425020 1290
rect 424968 1226 425020 1232
rect 424980 480 425008 1226
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 427268 3800 427320 3806
rect 427268 3742 427320 3748
rect 427280 480 427308 3742
rect 428476 480 428504 16546
rect 429660 3732 429712 3738
rect 429660 3674 429712 3680
rect 429672 480 429700 3674
rect 430868 480 430896 16546
rect 431972 1170 432000 29854
rect 438860 29844 438912 29850
rect 438860 29786 438912 29792
rect 432052 21820 432104 21826
rect 432052 21762 432104 21768
rect 432064 3398 432092 21762
rect 433340 17468 433392 17474
rect 433340 17410 433392 17416
rect 433352 16574 433380 17410
rect 434720 17400 434772 17406
rect 434720 17342 434772 17348
rect 434732 16574 434760 17342
rect 437480 17332 437532 17338
rect 437480 17274 437532 17280
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 432052 3392 432104 3398
rect 432052 3334 432104 3340
rect 433248 3392 433300 3398
rect 433248 3334 433300 3340
rect 431972 1142 432092 1170
rect 432064 480 432092 1142
rect 433260 480 433288 3334
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426134 -960 426246 326
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436744 6520 436796 6526
rect 436744 6462 436796 6468
rect 436756 480 436784 6462
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 17274
rect 438872 16574 438900 29786
rect 441620 29776 441672 29782
rect 441620 29718 441672 29724
rect 440238 22944 440294 22953
rect 440238 22879 440294 22888
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 3210 440280 22879
rect 440330 17232 440386 17241
rect 440330 17167 440386 17176
rect 440344 3398 440372 17167
rect 441632 16574 441660 29718
rect 443012 16574 443040 72830
rect 449900 72820 449952 72826
rect 449900 72762 449952 72768
rect 445022 31240 445078 31249
rect 445022 31175 445078 31184
rect 445036 16574 445064 31175
rect 445760 29708 445812 29714
rect 445760 29650 445812 29656
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 445036 16546 445156 16574
rect 440332 3392 440384 3398
rect 440332 3334 440384 3340
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 440252 3182 440372 3210
rect 440344 480 440372 3182
rect 441540 480 441568 3334
rect 442644 480 442672 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445022 4040 445078 4049
rect 445022 3975 445078 3984
rect 445036 480 445064 3975
rect 445128 3738 445156 16546
rect 445116 3732 445168 3738
rect 445116 3674 445168 3680
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 29650
rect 447140 21752 447192 21758
rect 447140 21694 447192 21700
rect 447152 16574 447180 21694
rect 448520 21684 448572 21690
rect 448520 21626 448572 21632
rect 447152 16546 447456 16574
rect 447428 480 447456 16546
rect 448532 3210 448560 21626
rect 449912 16574 449940 72762
rect 460940 72752 460992 72758
rect 460940 72694 460992 72700
rect 456800 35216 456852 35222
rect 456800 35158 456852 35164
rect 452660 29640 452712 29646
rect 452660 29582 452712 29588
rect 451280 18760 451332 18766
rect 451280 18702 451332 18708
rect 451292 16574 451320 18702
rect 452672 16574 452700 29582
rect 454038 22808 454094 22817
rect 454038 22743 454094 22752
rect 449912 16546 450952 16574
rect 451292 16546 451688 16574
rect 452672 16546 453344 16574
rect 448612 10328 448664 10334
rect 448612 10270 448664 10276
rect 448624 3398 448652 10270
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453316 480 453344 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 22743
rect 455418 18864 455474 18873
rect 455418 18799 455474 18808
rect 455432 16574 455460 18799
rect 455432 16546 455736 16574
rect 455708 480 455736 16546
rect 456812 3398 456840 35158
rect 456890 25528 456946 25537
rect 456890 25463 456946 25472
rect 456800 3392 456852 3398
rect 456800 3334 456852 3340
rect 456904 480 456932 25463
rect 459560 23452 459612 23458
rect 459560 23394 459612 23400
rect 458178 18728 458234 18737
rect 458178 18663 458234 18672
rect 458192 16574 458220 18663
rect 459572 16574 459600 23394
rect 460952 16574 460980 72694
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462424 354 462452 74598
rect 520936 74361 520964 231814
rect 527192 75041 527220 703520
rect 543476 699825 543504 703520
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 543462 699816 543518 699825
rect 543462 699751 543518 699760
rect 580446 683904 580502 683913
rect 580446 683839 580502 683848
rect 566464 670744 566516 670750
rect 580172 670744 580224 670750
rect 566464 670686 566516 670692
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 561968 311914 562272 311930
rect 561956 311908 562284 311914
rect 562008 311902 562232 311908
rect 561956 311850 562008 311856
rect 562232 311850 562284 311856
rect 552676 298790 552704 302124
rect 556080 300898 556108 302124
rect 556172 302110 557290 302138
rect 556068 300892 556120 300898
rect 556068 300834 556120 300840
rect 552664 298784 552716 298790
rect 552664 298726 552716 298732
rect 552676 88330 552704 298726
rect 556172 285666 556200 302110
rect 556160 285660 556212 285666
rect 556160 285602 556212 285608
rect 566476 99346 566504 670686
rect 580170 670647 580226 670656
rect 580354 644056 580410 644065
rect 580354 643991 580410 644000
rect 579986 617536 580042 617545
rect 579986 617471 580042 617480
rect 580000 616894 580028 617471
rect 579988 616888 580040 616894
rect 579988 616830 580040 616836
rect 580262 591016 580318 591025
rect 580262 590951 580318 590960
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 579802 511320 579858 511329
rect 579802 511255 579858 511264
rect 579816 510678 579844 511255
rect 579804 510672 579856 510678
rect 579804 510614 579856 510620
rect 580078 471472 580134 471481
rect 580078 471407 580134 471416
rect 579986 458144 580042 458153
rect 579986 458079 580042 458088
rect 580000 456822 580028 458079
rect 579988 456816 580040 456822
rect 579988 456758 580040 456764
rect 579986 444816 580042 444825
rect 579986 444751 580042 444760
rect 580000 444446 580028 444751
rect 579988 444440 580040 444446
rect 579988 444382 580040 444388
rect 579986 404968 580042 404977
rect 579986 404903 580042 404912
rect 580000 404394 580028 404903
rect 579988 404388 580040 404394
rect 579988 404330 580040 404336
rect 579986 378448 580042 378457
rect 579986 378383 580042 378392
rect 580000 378214 580028 378383
rect 579988 378208 580040 378214
rect 579988 378150 580040 378156
rect 579986 365120 580042 365129
rect 579986 365055 580042 365064
rect 580000 364410 580028 365055
rect 579988 364404 580040 364410
rect 579988 364346 580040 364352
rect 579988 351960 580040 351966
rect 579986 351928 579988 351937
rect 580040 351928 580042 351937
rect 579986 351863 580042 351872
rect 579986 338600 580042 338609
rect 579986 338535 580042 338544
rect 580000 338162 580028 338535
rect 566556 338156 566608 338162
rect 566556 338098 566608 338104
rect 579988 338156 580040 338162
rect 579988 338098 580040 338104
rect 566568 300898 566596 338098
rect 579802 325272 579858 325281
rect 579802 325207 579858 325216
rect 579816 324358 579844 325207
rect 579804 324352 579856 324358
rect 579804 324294 579856 324300
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580000 311914 580028 312015
rect 579988 311908 580040 311914
rect 579988 311850 580040 311856
rect 566556 300892 566608 300898
rect 566556 300834 566608 300840
rect 579988 298784 580040 298790
rect 579986 298752 579988 298761
rect 580040 298752 580042 298761
rect 579986 298687 580042 298696
rect 579988 285660 580040 285666
rect 579988 285602 580040 285608
rect 580000 285433 580028 285602
rect 579986 285424 580042 285433
rect 579986 285359 580042 285368
rect 579986 272232 580042 272241
rect 579986 272167 580042 272176
rect 580000 271930 580028 272167
rect 579988 271924 580040 271930
rect 579988 271866 580040 271872
rect 579986 258904 580042 258913
rect 579986 258839 580042 258848
rect 580000 258126 580028 258839
rect 579988 258120 580040 258126
rect 579988 258062 580040 258068
rect 579986 245576 580042 245585
rect 579986 245511 580042 245520
rect 580000 244322 580028 245511
rect 579988 244316 580040 244322
rect 579988 244258 580040 244264
rect 579802 232384 579858 232393
rect 579802 232319 579858 232328
rect 579816 231878 579844 232319
rect 579804 231872 579856 231878
rect 579804 231814 579856 231820
rect 579802 219056 579858 219065
rect 579802 218991 579858 219000
rect 579816 218074 579844 218991
rect 579804 218068 579856 218074
rect 579804 218010 579856 218016
rect 579986 205728 580042 205737
rect 579986 205663 579988 205672
rect 580040 205663 580042 205672
rect 579988 205634 580040 205640
rect 579986 179208 580042 179217
rect 579986 179143 580042 179152
rect 580000 178090 580028 179143
rect 579988 178084 580040 178090
rect 579988 178026 580040 178032
rect 579802 165880 579858 165889
rect 579802 165815 579858 165824
rect 579816 165646 579844 165815
rect 579804 165640 579856 165646
rect 579804 165582 579856 165588
rect 579986 139360 580042 139369
rect 579986 139295 580042 139304
rect 580000 138038 580028 139295
rect 579988 138032 580040 138038
rect 579988 137974 580040 137980
rect 580092 135930 580120 471407
rect 580184 193866 580212 537775
rect 580172 193860 580224 193866
rect 580172 193802 580224 193808
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580080 135924 580132 135930
rect 580080 135866 580132 135872
rect 580078 126032 580134 126041
rect 580078 125967 580134 125976
rect 580092 125662 580120 125967
rect 580080 125656 580132 125662
rect 580080 125598 580132 125604
rect 580078 99512 580134 99521
rect 580078 99447 580134 99456
rect 580092 99414 580120 99447
rect 580080 99408 580132 99414
rect 580080 99350 580132 99356
rect 566464 99340 566516 99346
rect 566464 99282 566516 99288
rect 552664 88324 552716 88330
rect 552664 88266 552716 88272
rect 580078 86184 580134 86193
rect 580078 86119 580134 86128
rect 580092 85610 580120 86119
rect 580080 85604 580132 85610
rect 580080 85546 580132 85552
rect 562324 75948 562376 75954
rect 562324 75890 562376 75896
rect 527178 75032 527234 75041
rect 527178 74967 527234 74976
rect 550640 74588 550692 74594
rect 550640 74530 550692 74536
rect 520922 74352 520978 74361
rect 520922 74287 520978 74296
rect 465172 73840 465224 73846
rect 465172 73782 465224 73788
rect 463700 31748 463752 31754
rect 463700 31690 463752 31696
rect 463712 16574 463740 31690
rect 465184 16574 465212 73782
rect 478878 72856 478934 72865
rect 478878 72791 478934 72800
rect 471980 72684 472032 72690
rect 471980 72626 472032 72632
rect 470600 31680 470652 31686
rect 470600 31622 470652 31628
rect 467840 26920 467892 26926
rect 467840 26862 467892 26868
rect 467852 16574 467880 26862
rect 469220 19984 469272 19990
rect 469220 19926 469272 19932
rect 469232 16574 469260 19926
rect 463712 16546 464016 16574
rect 465184 16546 465856 16574
rect 467852 16546 468248 16574
rect 469232 16546 469904 16574
rect 463988 480 464016 16546
rect 465172 3664 465224 3670
rect 465172 3606 465224 3612
rect 465184 480 465212 3606
rect 462750 354 462862 480
rect 462424 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 467472 14476 467524 14482
rect 467472 14418 467524 14424
rect 467484 480 467512 14418
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 469876 480 469904 16546
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 31622
rect 471992 16574 472020 72626
rect 474738 65512 474794 65521
rect 474738 65447 474794 65456
rect 473358 31104 473414 31113
rect 473358 31039 473414 31048
rect 471992 16546 472296 16574
rect 472268 480 472296 16546
rect 473372 3398 473400 31039
rect 473450 19952 473506 19961
rect 473450 19887 473506 19896
rect 473360 3392 473412 3398
rect 473360 3334 473412 3340
rect 473464 480 473492 19887
rect 474752 16574 474780 65447
rect 477500 31612 477552 31618
rect 477500 31554 477552 31560
rect 476118 21312 476174 21321
rect 476118 21247 476174 21256
rect 476132 16574 476160 21247
rect 477512 16574 477540 31554
rect 474752 16546 475792 16574
rect 476132 16546 476528 16574
rect 477512 16546 478184 16574
rect 474188 3392 474240 3398
rect 474188 3334 474240 3340
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474200 354 474228 3334
rect 475764 480 475792 16546
rect 474526 354 474638 480
rect 474200 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478052 3528 478104 3534
rect 478052 3470 478104 3476
rect 478064 3398 478092 3470
rect 478052 3392 478104 3398
rect 478052 3334 478104 3340
rect 478156 480 478184 16546
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478892 354 478920 72791
rect 480258 72720 480314 72729
rect 480258 72655 480314 72664
rect 480272 16574 480300 72655
rect 514760 72616 514812 72622
rect 498198 72584 498254 72593
rect 514760 72558 514812 72564
rect 498198 72519 498254 72528
rect 481640 31544 481692 31550
rect 481640 31486 481692 31492
rect 480272 16546 480576 16574
rect 480548 480 480576 16546
rect 481652 8294 481680 31486
rect 490012 31476 490064 31482
rect 490012 31418 490064 31424
rect 481732 21616 481784 21622
rect 481732 21558 481784 21564
rect 481640 8288 481692 8294
rect 481640 8230 481692 8236
rect 481744 480 481772 21558
rect 484400 21548 484452 21554
rect 484400 21490 484452 21496
rect 484412 16574 484440 21490
rect 488540 21480 488592 21486
rect 488540 21422 488592 21428
rect 488552 16574 488580 21422
rect 484412 16546 484808 16574
rect 488552 16546 488856 16574
rect 482468 8288 482520 8294
rect 482468 8230 482520 8236
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482480 354 482508 8230
rect 484032 3596 484084 3602
rect 484032 3538 484084 3544
rect 484044 480 484072 3538
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486424 11756 486476 11762
rect 486424 11698 486476 11704
rect 486436 480 486464 11698
rect 487620 3392 487672 3398
rect 487620 3334 487672 3340
rect 487632 480 487660 3334
rect 488828 480 488856 16546
rect 490024 6914 490052 31418
rect 496820 31408 496872 31414
rect 496820 31350 496872 31356
rect 492678 30968 492734 30977
rect 492678 30903 492734 30912
rect 491300 21412 491352 21418
rect 491300 21354 491352 21360
rect 491312 16574 491340 21354
rect 492692 16574 492720 30903
rect 495440 23384 495492 23390
rect 495440 23326 495492 23332
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 489932 6886 490052 6914
rect 489932 480 489960 6886
rect 491116 3460 491168 3466
rect 491116 3402 491168 3408
rect 491128 480 491156 3402
rect 492324 480 492352 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494702 3904 494758 3913
rect 494702 3839 494758 3848
rect 494716 480 494744 3839
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 23326
rect 496832 16574 496860 31350
rect 496832 16546 497136 16574
rect 497108 480 497136 16546
rect 498212 480 498240 72519
rect 503720 31340 503772 31346
rect 503720 31282 503772 31288
rect 498292 23316 498344 23322
rect 498292 23258 498344 23264
rect 498304 16574 498332 23258
rect 502340 23248 502392 23254
rect 502340 23190 502392 23196
rect 502352 16574 502380 23190
rect 498304 16546 498976 16574
rect 502352 16546 503024 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500592 5092 500644 5098
rect 500592 5034 500644 5040
rect 500604 480 500632 5034
rect 501788 5024 501840 5030
rect 501788 4966 501840 4972
rect 501800 480 501828 4966
rect 502996 480 503024 16546
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 31282
rect 510620 31272 510672 31278
rect 510620 31214 510672 31220
rect 506480 23180 506532 23186
rect 506480 23122 506532 23128
rect 505374 3768 505430 3777
rect 505374 3703 505430 3712
rect 505388 480 505416 3703
rect 506492 480 506520 23122
rect 509238 22672 509294 22681
rect 509238 22607 509294 22616
rect 509252 16574 509280 22607
rect 510632 16574 510660 31214
rect 513380 23112 513432 23118
rect 513380 23054 513432 23060
rect 509252 16546 509648 16574
rect 510632 16546 511304 16574
rect 507214 13016 507270 13025
rect 507214 12951 507270 12960
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 12951
rect 508870 5400 508926 5409
rect 508870 5335 508926 5344
rect 508884 480 508912 5335
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511276 480 511304 16546
rect 512458 5264 512514 5273
rect 512458 5199 512514 5208
rect 512472 480 512500 5199
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513392 354 513420 23054
rect 514772 16574 514800 72558
rect 549260 32496 549312 32502
rect 549260 32438 549312 32444
rect 517520 31204 517572 31210
rect 517520 31146 517572 31152
rect 516140 23044 516192 23050
rect 516140 22986 516192 22992
rect 516152 16574 516180 22986
rect 517532 16574 517560 31146
rect 524420 31136 524472 31142
rect 524420 31078 524472 31084
rect 521660 31068 521712 31074
rect 521660 31010 521712 31016
rect 520280 22976 520332 22982
rect 520280 22918 520332 22924
rect 514772 16546 515536 16574
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 514760 6452 514812 6458
rect 514760 6394 514812 6400
rect 514772 480 514800 6394
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515508 354 515536 16546
rect 517164 480 517192 16546
rect 515926 354 516038 480
rect 515508 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519544 4956 519596 4962
rect 519544 4898 519596 4904
rect 519556 480 519584 4898
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 22918
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 31010
rect 523040 22908 523092 22914
rect 523040 22850 523092 22856
rect 523052 16574 523080 22850
rect 524432 16574 524460 31078
rect 531320 24608 531372 24614
rect 531320 24550 531372 24556
rect 527178 24304 527234 24313
rect 527178 24239 527234 24248
rect 527192 16574 527220 24239
rect 528558 18592 528614 18601
rect 528558 18527 528614 18536
rect 523052 16546 523816 16574
rect 524432 16546 525472 16574
rect 527192 16546 527864 16574
rect 523040 4888 523092 4894
rect 523040 4830 523092 4836
rect 523052 480 523080 4830
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 525444 480 525472 16546
rect 526626 6488 526682 6497
rect 526626 6423 526682 6432
rect 526640 480 526668 6423
rect 527836 480 527864 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 354 528600 18527
rect 530122 6352 530178 6361
rect 530122 6287 530178 6296
rect 530136 480 530164 6287
rect 531332 480 531360 24550
rect 534080 24540 534132 24546
rect 534080 24482 534132 24488
rect 534092 16574 534120 24482
rect 538220 24472 538272 24478
rect 538220 24414 538272 24420
rect 535460 18692 535512 18698
rect 535460 18634 535512 18640
rect 535472 16574 535500 18634
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 532056 15904 532108 15910
rect 532056 15846 532108 15852
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 528990 -960 529102 326
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532068 354 532096 15846
rect 533710 3632 533766 3641
rect 533710 3567 533766 3576
rect 533724 480 533752 3567
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537206 3496 537262 3505
rect 537206 3431 537262 3440
rect 537220 480 537248 3431
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 24414
rect 540980 24404 541032 24410
rect 540980 24346 541032 24352
rect 540992 16574 541020 24346
rect 547880 24336 547932 24342
rect 547880 24278 547932 24284
rect 545118 24168 545174 24177
rect 545118 24103 545174 24112
rect 545132 16574 545160 24103
rect 547892 16574 547920 24278
rect 549272 16574 549300 32438
rect 550652 16574 550680 74530
rect 558920 72548 558972 72554
rect 558920 72490 558972 72496
rect 556160 25696 556212 25702
rect 556160 25638 556212 25644
rect 552020 24268 552072 24274
rect 552020 24210 552072 24216
rect 552032 16574 552060 24210
rect 553400 18624 553452 18630
rect 553400 18566 553452 18572
rect 553412 16574 553440 18566
rect 540992 16546 542032 16574
rect 545132 16546 545528 16574
rect 547892 16546 548656 16574
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 540796 6384 540848 6390
rect 540796 6326 540848 6332
rect 539600 3324 539652 3330
rect 539600 3266 539652 3272
rect 539612 480 539640 3266
rect 540808 480 540836 6326
rect 542004 480 542032 16546
rect 544384 6316 544436 6322
rect 544384 6258 544436 6264
rect 543188 4140 543240 4146
rect 543188 4082 543240 4088
rect 543200 480 543228 4082
rect 544396 480 544424 6258
rect 545500 480 545528 16546
rect 547878 5128 547934 5137
rect 547878 5063 547934 5072
rect 546684 3732 546736 3738
rect 546684 3674 546736 3680
rect 546696 480 546724 3674
rect 547892 480 547920 5063
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 550284 480 550312 16546
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 554964 7676 555016 7682
rect 554964 7618 555016 7624
rect 554976 480 555004 7618
rect 556172 480 556200 25638
rect 556252 17264 556304 17270
rect 556252 17206 556304 17212
rect 556264 16574 556292 17206
rect 558932 16574 558960 72490
rect 560300 22840 560352 22846
rect 560300 22782 560352 22788
rect 560312 16574 560340 22782
rect 556264 16546 556936 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558552 7608 558604 7614
rect 558552 7550 558604 7556
rect 558564 480 558592 7550
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562046 7712 562102 7721
rect 562046 7647 562102 7656
rect 562060 480 562088 7647
rect 562336 6866 562364 75890
rect 580184 74497 580212 192471
rect 580170 74488 580226 74497
rect 580170 74423 580226 74432
rect 580276 73137 580304 590951
rect 580368 74769 580396 643991
rect 580460 174350 580488 683839
rect 580538 630864 580594 630873
rect 580538 630799 580594 630808
rect 580448 174344 580500 174350
rect 580448 174286 580500 174292
rect 580446 152688 580502 152697
rect 580446 152623 580502 152632
rect 580354 74760 580410 74769
rect 580354 74695 580410 74704
rect 580460 74458 580488 152623
rect 580552 142866 580580 630799
rect 580630 577688 580686 577697
rect 580630 577623 580686 577632
rect 580540 142860 580592 142866
rect 580540 142802 580592 142808
rect 580644 137290 580672 577623
rect 580814 524512 580870 524521
rect 580814 524447 580870 524456
rect 580722 484664 580778 484673
rect 580722 484599 580778 484608
rect 580632 137284 580684 137290
rect 580632 137226 580684 137232
rect 580538 112840 580594 112849
rect 580538 112775 580594 112784
rect 580552 74526 580580 112775
rect 580540 74520 580592 74526
rect 580540 74462 580592 74468
rect 580448 74452 580500 74458
rect 580448 74394 580500 74400
rect 580262 73128 580318 73137
rect 580736 73098 580764 484599
rect 580828 135998 580856 524447
rect 580906 431624 580962 431633
rect 580906 431559 580962 431568
rect 580816 135992 580868 135998
rect 580816 135934 580868 135940
rect 580920 74633 580948 431559
rect 580906 74624 580962 74633
rect 580906 74559 580962 74568
rect 580262 73063 580318 73072
rect 580724 73092 580776 73098
rect 580724 73034 580776 73040
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580184 72010 580212 72927
rect 581000 72480 581052 72486
rect 581000 72422 581052 72428
rect 581090 72448 581146 72457
rect 580172 72004 580224 72010
rect 580172 71946 580224 71952
rect 580264 71052 580316 71058
rect 580264 70994 580316 71000
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580276 33153 580304 70994
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 574100 32428 574152 32434
rect 574100 32370 574152 32376
rect 571340 28280 571392 28286
rect 571340 28222 571392 28228
rect 565820 25628 565872 25634
rect 565820 25570 565872 25576
rect 565832 16574 565860 25570
rect 567200 24200 567252 24206
rect 567200 24142 567252 24148
rect 567212 16574 567240 24142
rect 569960 24132 570012 24138
rect 569960 24074 570012 24080
rect 569972 16574 570000 24074
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 569972 16546 570368 16574
rect 564438 7576 564494 7585
rect 564438 7511 564494 7520
rect 562324 6860 562376 6866
rect 562324 6802 562376 6808
rect 563242 4992 563298 5001
rect 563242 4927 563298 4936
rect 563256 480 563284 4927
rect 564452 480 564480 7511
rect 565634 4856 565690 4865
rect 565634 4791 565690 4800
rect 565648 480 565676 4791
rect 566844 480 566872 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 569132 6248 569184 6254
rect 569132 6190 569184 6196
rect 569144 480 569172 6190
rect 570340 480 570368 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 28222
rect 572720 25560 572772 25566
rect 572720 25502 572772 25508
rect 572732 16574 572760 25502
rect 574112 16574 574140 32370
rect 580172 22772 580224 22778
rect 580172 22714 580224 22720
rect 580184 19825 580212 22714
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 572732 16546 573496 16574
rect 574112 16546 575152 16574
rect 572720 6180 572772 6186
rect 572720 6122 572772 6128
rect 572732 480 572760 6122
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 575124 480 575152 16546
rect 578606 8936 578662 8945
rect 578606 8871 578662 8880
rect 576306 6216 576362 6225
rect 576306 6151 576362 6160
rect 576320 480 576348 6151
rect 577412 4820 577464 4826
rect 577412 4762 577464 4768
rect 577424 480 577452 4762
rect 578620 480 578648 8871
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 581012 480 581040 72422
rect 581090 72383 581146 72392
rect 581104 16574 581132 72383
rect 581104 16546 581776 16574
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3330 566888 3386 566944
rect 2778 553852 2834 553888
rect 2778 553832 2780 553852
rect 2780 553832 2832 553852
rect 2832 553832 2834 553852
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 2778 501744 2834 501800
rect 2778 462596 2834 462632
rect 2778 462576 2780 462596
rect 2780 462576 2832 462596
rect 2832 462576 2834 462596
rect 2778 449520 2834 449576
rect 3146 410488 3202 410544
rect 2778 397468 2780 397488
rect 2780 397468 2832 397488
rect 2832 397468 2834 397488
rect 2778 397432 2834 397468
rect 3330 358400 3386 358456
rect 2778 345344 2834 345400
rect 3330 319232 3386 319288
rect 3238 306176 3294 306232
rect 3238 293120 3294 293176
rect 3238 267144 3294 267200
rect 3146 254088 3202 254144
rect 3054 241032 3110 241088
rect 3146 214920 3202 214976
rect 2962 201864 3018 201920
rect 3146 188808 3202 188864
rect 3146 162868 3148 162888
rect 3148 162868 3200 162888
rect 3200 162868 3202 162888
rect 3146 162832 3202 162868
rect 3146 149776 3202 149832
rect 3514 671200 3570 671256
rect 3606 632032 3662 632088
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3422 136720 3478 136776
rect 3330 84632 3386 84688
rect 2870 32408 2926 32464
rect 3698 579944 3754 580000
rect 3790 527856 3846 527912
rect 3974 475632 4030 475688
rect 3882 423544 3938 423600
rect 4066 371320 4122 371376
rect 3514 73752 3570 73808
rect 3514 71576 3570 71632
rect 3790 110608 3846 110664
rect 3698 97552 3754 97608
rect 4894 75112 4950 75168
rect 5170 75248 5226 75304
rect 4986 74024 5042 74080
rect 4802 73616 4858 73672
rect 395342 240080 395398 240136
rect 395526 239944 395582 240000
rect 392582 232328 392638 232384
rect 380162 231104 380218 231160
rect 22742 72528 22798 72584
rect 3606 58520 3662 58576
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3422 19352 3478 19408
rect 3514 6432 3570 6488
rect 1674 3440 1730 3496
rect 570 3304 626 3360
rect 18234 6160 18290 6216
rect 17038 3576 17094 3632
rect 34794 8880 34850 8936
rect 38382 9016 38438 9072
rect 37186 4800 37242 4856
rect 53746 9152 53802 9208
rect 52550 6296 52606 6352
rect 56046 6432 56102 6488
rect 54942 3712 54998 3768
rect 71502 10240 71558 10296
rect 70306 7520 70362 7576
rect 114006 138624 114062 138680
rect 113638 131164 113694 131200
rect 113638 131144 113640 131164
rect 113640 131144 113692 131164
rect 113692 131144 113694 131164
rect 113546 128968 113602 129024
rect 113546 127472 113602 127528
rect 113638 126792 113694 126848
rect 113638 125432 113694 125488
rect 113638 123800 113694 123856
rect 113638 122748 113640 122768
rect 113640 122748 113692 122768
rect 113692 122748 113694 122768
rect 113638 122712 113694 122748
rect 113638 121216 113694 121272
rect 113638 119720 113694 119776
rect 113638 118224 113694 118280
rect 113638 116728 113694 116784
rect 113546 115232 113602 115288
rect 113638 113092 113640 113112
rect 113640 113092 113692 113112
rect 113692 113092 113694 113112
rect 113638 113056 113694 113092
rect 113638 111732 113640 111752
rect 113640 111732 113692 111752
rect 113692 111732 113694 111752
rect 113638 111696 113694 111732
rect 113638 110372 113640 110392
rect 113640 110372 113692 110392
rect 113692 110372 113694 110392
rect 113638 110336 113694 110372
rect 113638 108840 113694 108896
rect 113638 107480 113694 107536
rect 113546 105848 113602 105904
rect 113638 104796 113640 104816
rect 113640 104796 113692 104816
rect 113692 104796 113694 104816
rect 113638 104760 113694 104796
rect 113730 103128 113786 103184
rect 113822 101768 113878 101824
rect 113914 91024 113970 91080
rect 114006 89664 114062 89720
rect 114098 88168 114154 88224
rect 114190 86808 114246 86864
rect 114282 85312 114338 85368
rect 115294 137264 115350 137320
rect 114466 82320 114522 82376
rect 114374 80824 114430 80880
rect 114466 78648 114522 78704
rect 114374 76608 114430 76664
rect 114466 75384 114522 75440
rect 115570 133184 115626 133240
rect 115294 100272 115350 100328
rect 115386 98776 115442 98832
rect 115478 93744 115534 93800
rect 115754 96668 115810 96724
rect 115662 95172 115718 95228
rect 115570 92384 115626 92440
rect 138110 195880 138166 195936
rect 140410 195880 140466 195936
rect 141422 195916 141424 195936
rect 141424 195916 141476 195936
rect 141476 195916 141478 195936
rect 141422 195880 141478 195916
rect 158902 195872 158958 195928
rect 160834 195880 160890 195936
rect 157154 195608 157210 195664
rect 139398 195472 139454 195528
rect 140870 191800 140926 191856
rect 140778 190848 140834 190904
rect 140962 191664 141018 191720
rect 144550 190984 144606 191040
rect 144458 190576 144514 190632
rect 145838 189760 145894 189816
rect 140962 184320 141018 184376
rect 140870 184184 140926 184240
rect 144734 183776 144790 183832
rect 144642 183640 144698 183696
rect 140778 182552 140834 182608
rect 145194 181192 145250 181248
rect 144642 180920 144698 180976
rect 149334 179424 149390 179480
rect 148046 179288 148102 179344
rect 142666 179016 142722 179072
rect 144090 178880 144146 178936
rect 141606 178744 141662 178800
rect 140502 175616 140558 175672
rect 139674 137944 139730 138000
rect 157798 179580 157854 179616
rect 157798 179560 157800 179580
rect 157800 179560 157852 179580
rect 157852 179560 157854 179580
rect 158534 179560 158590 179616
rect 157798 178084 157854 178120
rect 157798 178064 157800 178084
rect 157800 178064 157852 178084
rect 157852 178064 157854 178084
rect 158534 178064 158590 178120
rect 149334 175344 149390 175400
rect 154578 175344 154634 175400
rect 147494 174120 147550 174176
rect 161570 138760 161626 138816
rect 167826 137536 167882 137592
rect 169390 137400 169446 137456
rect 175462 132368 175518 132424
rect 175370 130056 175426 130112
rect 175554 128288 175610 128344
rect 115846 83204 115902 83260
rect 89166 10376 89222 10432
rect 87970 7656 88026 7712
rect 91558 7792 91614 7848
rect 90362 4936 90418 4992
rect 105726 9288 105782 9344
rect 109314 9424 109370 9480
rect 108118 6568 108174 6624
rect 121642 71984 121698 72040
rect 121550 71848 121606 71904
rect 121918 72528 121974 72584
rect 122838 71984 122894 72040
rect 122930 71848 122986 71904
rect 124218 72120 124274 72176
rect 124402 71984 124458 72040
rect 124494 71848 124550 71904
rect 125690 72256 125746 72312
rect 125598 72120 125654 72176
rect 125782 71984 125838 72040
rect 125874 71848 125930 71904
rect 127070 71984 127126 72040
rect 126978 71848 127034 71904
rect 128542 73072 128598 73128
rect 128450 72120 128506 72176
rect 128358 71984 128414 72040
rect 128634 71848 128690 71904
rect 129738 72120 129794 72176
rect 130014 71984 130070 72040
rect 129922 71848 129978 71904
rect 123482 3576 123538 3632
rect 124678 3440 124734 3496
rect 131210 71984 131266 72040
rect 131118 71848 131174 71904
rect 132222 71984 132278 72040
rect 132406 71848 132462 71904
rect 133694 72120 133750 72176
rect 133602 71984 133658 72040
rect 133786 71848 133842 71904
rect 135074 72120 135130 72176
rect 134982 71984 135038 72040
rect 135166 71848 135222 71904
rect 136454 72120 136510 72176
rect 136362 71984 136418 72040
rect 136178 71848 136234 71904
rect 136546 71848 136602 71904
rect 137834 71984 137890 72040
rect 137926 71848 137982 71904
rect 137650 3576 137706 3632
rect 139030 71984 139086 72040
rect 139306 72120 139362 72176
rect 138938 71848 138994 71904
rect 139122 71848 139178 71904
rect 140318 72120 140374 72176
rect 140594 71984 140650 72040
rect 140410 71848 140466 71904
rect 140686 71848 140742 71904
rect 141974 71984 142030 72040
rect 142066 71848 142122 71904
rect 143262 72120 143318 72176
rect 143354 71984 143410 72040
rect 143170 71848 143226 71904
rect 143446 71848 143502 71904
rect 144734 72120 144790 72176
rect 144642 71984 144698 72040
rect 144550 71848 144606 71904
rect 144826 71848 144882 71904
rect 146022 72120 146078 72176
rect 146206 71984 146262 72040
rect 146114 71848 146170 71904
rect 147494 72256 147550 72312
rect 147402 72120 147458 72176
rect 147586 71984 147642 72040
rect 147310 71848 147366 71904
rect 148690 72664 148746 72720
rect 148874 72800 148930 72856
rect 148966 72664 149022 72720
rect 148782 72392 148838 72448
rect 140042 3440 140098 3496
rect 149978 72664 150034 72720
rect 150346 72800 150402 72856
rect 150162 72528 150218 72584
rect 150070 72392 150126 72448
rect 151634 72800 151690 72856
rect 151542 72664 151598 72720
rect 151726 72392 151782 72448
rect 152922 72800 152978 72856
rect 153106 72936 153162 72992
rect 153014 72664 153070 72720
rect 152830 72528 152886 72584
rect 154118 72800 154174 72856
rect 154210 72664 154266 72720
rect 154302 72392 154358 72448
rect 154486 72528 154542 72584
rect 154762 74432 154818 74488
rect 155498 72936 155554 72992
rect 155866 72664 155922 72720
rect 155774 72392 155830 72448
rect 155682 72256 155738 72312
rect 156142 74568 156198 74624
rect 156970 72800 157026 72856
rect 156878 72664 156934 72720
rect 157062 72528 157118 72584
rect 157062 72256 157118 72312
rect 157246 72664 157302 72720
rect 157154 71984 157210 72040
rect 157798 71984 157854 72040
rect 158350 72800 158406 72856
rect 158534 72664 158590 72720
rect 158626 72528 158682 72584
rect 158442 72392 158498 72448
rect 158810 73072 158866 73128
rect 158902 72120 158958 72176
rect 155406 4936 155462 4992
rect 156602 4800 156658 4856
rect 157798 3304 157854 3360
rect 159638 72392 159694 72448
rect 159914 72800 159970 72856
rect 160006 72664 160062 72720
rect 160282 72256 160338 72312
rect 161018 72800 161074 72856
rect 161110 72664 161166 72720
rect 161294 73072 161350 73128
rect 161386 72664 161442 72720
rect 161202 72528 161258 72584
rect 161294 72392 161350 72448
rect 161662 74704 161718 74760
rect 161662 74468 161664 74488
rect 161664 74468 161716 74488
rect 161716 74468 161718 74488
rect 161662 74432 161718 74468
rect 161662 74160 161718 74216
rect 162398 73072 162454 73128
rect 162490 72664 162546 72720
rect 162490 72564 162492 72584
rect 162492 72564 162544 72584
rect 162544 72564 162546 72584
rect 162490 72528 162546 72564
rect 162674 72800 162730 72856
rect 162766 72664 162822 72720
rect 162582 72392 162638 72448
rect 163042 73072 163098 73128
rect 163318 72256 163374 72312
rect 163962 72800 164018 72856
rect 164238 74704 164294 74760
rect 164238 74432 164294 74488
rect 164146 72664 164202 72720
rect 164054 72528 164110 72584
rect 164422 74160 164478 74216
rect 164698 74704 164754 74760
rect 164882 74160 164938 74216
rect 164882 72800 164938 72856
rect 164698 71304 164754 71360
rect 165342 72800 165398 72856
rect 165250 72664 165306 72720
rect 165526 72664 165582 72720
rect 165434 72528 165490 72584
rect 165526 72256 165582 72312
rect 160834 3712 160890 3768
rect 165526 70080 165582 70136
rect 166354 72800 166410 72856
rect 166538 72664 166594 72720
rect 166814 73344 166870 73400
rect 167274 74432 167330 74488
rect 167366 74296 167422 74352
rect 167458 74160 167514 74216
rect 167458 74024 167514 74080
rect 167734 74840 167790 74896
rect 167274 72800 167330 72856
rect 168286 74840 168342 74896
rect 168194 74568 168250 74624
rect 168010 73072 168066 73128
rect 168562 72664 168618 72720
rect 168562 72120 168618 72176
rect 169114 73752 169170 73808
rect 169206 73616 169262 73672
rect 169390 74704 169446 74760
rect 169574 74704 169630 74760
rect 169482 73888 169538 73944
rect 169390 73752 169446 73808
rect 169298 73480 169354 73536
rect 172794 75112 172850 75168
rect 172610 74840 172666 74896
rect 170862 74024 170918 74080
rect 172334 74704 172390 74760
rect 172610 74568 172666 74624
rect 172794 74568 172850 74624
rect 172334 73752 172390 73808
rect 172886 72392 172942 72448
rect 176750 126928 176806 126984
rect 176658 119720 176714 119776
rect 178038 125432 178094 125488
rect 178130 122440 178186 122496
rect 176842 111696 176898 111752
rect 176658 110336 176714 110392
rect 175922 108976 175978 109032
rect 178498 124072 178554 124128
rect 178406 121216 178462 121272
rect 178590 118224 178646 118280
rect 178314 115232 178370 115288
rect 178866 131144 178922 131200
rect 178774 116728 178830 116784
rect 178682 113056 178738 113112
rect 178222 107480 178278 107536
rect 178038 105984 178094 106040
rect 178038 104488 178094 104544
rect 178038 102992 178094 103048
rect 178038 101632 178094 101688
rect 178038 100136 178094 100192
rect 178038 98776 178094 98832
rect 178038 97280 178094 97336
rect 178038 95140 178040 95160
rect 178040 95140 178092 95160
rect 178092 95140 178094 95160
rect 178038 95104 178094 95140
rect 178038 93780 178040 93800
rect 178040 93780 178092 93800
rect 178092 93780 178094 93800
rect 178038 93744 178094 93780
rect 178038 92248 178094 92304
rect 178038 90888 178094 90944
rect 178038 89392 178094 89448
rect 178038 88032 178094 88088
rect 178038 86536 178094 86592
rect 178038 85040 178094 85096
rect 178038 83680 178094 83736
rect 178038 82184 178094 82240
rect 178682 78648 178738 78704
rect 178038 76608 178094 76664
rect 179234 80824 179290 80880
rect 173898 32680 173954 32736
rect 172518 25608 172574 25664
rect 169666 8064 169722 8120
rect 187698 32544 187754 32600
rect 191838 32408 191894 32464
rect 190458 27104 190514 27160
rect 193310 4664 193366 4720
rect 209778 34040 209834 34096
rect 210974 12144 211030 12200
rect 223578 20168 223634 20224
rect 225142 12824 225198 12880
rect 228730 6840 228786 6896
rect 226430 6024 226486 6080
rect 241518 33904 241574 33960
rect 244278 20032 244334 20088
rect 242990 13640 243046 13696
rect 246394 6704 246450 6760
rect 262218 33768 262274 33824
rect 264150 15136 264206 15192
rect 278778 26968 278834 27024
rect 278318 7928 278374 7984
rect 280710 13504 280766 13560
rect 281906 7792 281962 7848
rect 298098 35264 298154 35320
rect 295614 16224 295670 16280
rect 297270 15000 297326 15056
rect 299662 9016 299718 9072
rect 314658 29552 314714 29608
rect 316038 17584 316094 17640
rect 316222 14864 316278 14920
rect 332598 35128 332654 35184
rect 331218 10376 331274 10432
rect 350538 21392 350594 21448
rect 332690 14728 332746 14784
rect 334622 10240 334678 10296
rect 349158 16088 349214 16144
rect 349250 12008 349306 12064
rect 352838 11872 352894 11928
rect 367098 26832 367154 26888
rect 365718 13368 365774 13424
rect 365810 11736 365866 11792
rect 370134 13232 370190 13288
rect 396998 74160 397054 74216
rect 386418 24384 386474 24440
rect 385958 6568 386014 6624
rect 387798 14592 387854 14648
rect 406014 15952 406070 16008
rect 402518 14456 402574 14512
rect 403622 11600 403678 11656
rect 404818 5480 404874 5536
rect 420918 17448 420974 17504
rect 420182 15816 420238 15872
rect 418526 13096 418582 13152
rect 423770 17312 423826 17368
rect 440238 22888 440294 22944
rect 440330 17176 440386 17232
rect 445022 31184 445078 31240
rect 445022 3984 445078 4040
rect 454038 22752 454094 22808
rect 455418 18808 455474 18864
rect 456890 25472 456946 25528
rect 458178 18672 458234 18728
rect 543462 699760 543518 699816
rect 580446 683848 580502 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580354 644000 580410 644056
rect 579986 617480 580042 617536
rect 580262 590960 580318 591016
rect 580170 564304 580226 564360
rect 580170 537784 580226 537840
rect 579802 511264 579858 511320
rect 580078 471416 580134 471472
rect 579986 458088 580042 458144
rect 579986 444760 580042 444816
rect 579986 404912 580042 404968
rect 579986 378392 580042 378448
rect 579986 365064 580042 365120
rect 579986 351908 579988 351928
rect 579988 351908 580040 351928
rect 580040 351908 580042 351928
rect 579986 351872 580042 351908
rect 579986 338544 580042 338600
rect 579802 325216 579858 325272
rect 579986 312024 580042 312080
rect 579986 298732 579988 298752
rect 579988 298732 580040 298752
rect 580040 298732 580042 298752
rect 579986 298696 580042 298732
rect 579986 285368 580042 285424
rect 579986 272176 580042 272232
rect 579986 258848 580042 258904
rect 579986 245520 580042 245576
rect 579802 232328 579858 232384
rect 579802 219000 579858 219056
rect 579986 205692 580042 205728
rect 579986 205672 579988 205692
rect 579988 205672 580040 205692
rect 580040 205672 580042 205692
rect 579986 179152 580042 179208
rect 579802 165824 579858 165880
rect 579986 139304 580042 139360
rect 580170 192480 580226 192536
rect 580078 125976 580134 126032
rect 580078 99456 580134 99512
rect 580078 86128 580134 86184
rect 527178 74976 527234 75032
rect 520922 74296 520978 74352
rect 478878 72800 478934 72856
rect 474738 65456 474794 65512
rect 473358 31048 473414 31104
rect 473450 19896 473506 19952
rect 476118 21256 476174 21312
rect 480258 72664 480314 72720
rect 498198 72528 498254 72584
rect 492678 30912 492734 30968
rect 494702 3848 494758 3904
rect 505374 3712 505430 3768
rect 509238 22616 509294 22672
rect 507214 12960 507270 13016
rect 508870 5344 508926 5400
rect 512458 5208 512514 5264
rect 527178 24248 527234 24304
rect 528558 18536 528614 18592
rect 526626 6432 526682 6488
rect 530122 6296 530178 6352
rect 533710 3576 533766 3632
rect 537206 3440 537262 3496
rect 545118 24112 545174 24168
rect 547878 5072 547934 5128
rect 562046 7656 562102 7712
rect 580170 74432 580226 74488
rect 580538 630808 580594 630864
rect 580446 152632 580502 152688
rect 580354 74704 580410 74760
rect 580630 577632 580686 577688
rect 580814 524456 580870 524512
rect 580722 484608 580778 484664
rect 580538 112784 580594 112840
rect 580262 73072 580318 73128
rect 580906 431568 580962 431624
rect 580906 74568 580962 74624
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580262 33088 580318 33144
rect 564438 7520 564494 7576
rect 563242 4936 563298 4992
rect 565634 4800 565690 4856
rect 580170 19760 580226 19816
rect 578606 8880 578662 8936
rect 576306 6160 576362 6216
rect 580170 6568 580226 6624
rect 581090 72392 581146 72448
rect 583390 3304 583446 3360
<< metal3 >>
rect 542670 699756 542676 699820
rect 542740 699818 542746 699820
rect 543457 699818 543523 699821
rect 542740 699816 543523 699818
rect 542740 699760 543462 699816
rect 543518 699760 543523 699816
rect 542740 699758 543523 699760
rect 542740 699756 542746 699758
rect 543457 699755 543523 699758
rect -960 697220 480 697460
rect 580206 697172 580212 697236
rect 580276 697234 580282 697236
rect 583520 697234 584960 697324
rect 580276 697174 584960 697234
rect 580276 697172 580282 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580441 683906 580507 683909
rect 583520 683906 584960 683996
rect 580441 683904 584960 683906
rect 580441 683848 580446 683904
rect 580502 683848 584960 683904
rect 580441 683846 584960 683848
rect 580441 683843 580507 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3366 658202 3372 658204
rect -960 658142 3372 658202
rect -960 658052 480 658142
rect 3366 658140 3372 658142
rect 3436 658140 3442 658204
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580349 644058 580415 644061
rect 583520 644058 584960 644148
rect 580349 644056 584960 644058
rect 580349 644000 580354 644056
rect 580410 644000 584960 644056
rect 580349 643998 584960 644000
rect 580349 643995 580415 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3601 632090 3667 632093
rect -960 632088 3667 632090
rect -960 632032 3606 632088
rect 3662 632032 3667 632088
rect -960 632030 3667 632032
rect -960 631940 480 632030
rect 3601 632027 3667 632030
rect 580533 630866 580599 630869
rect 583520 630866 584960 630956
rect 580533 630864 584960 630866
rect 580533 630808 580538 630864
rect 580594 630808 584960 630864
rect 580533 630806 584960 630808
rect 580533 630803 580599 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 579981 617538 580047 617541
rect 583520 617538 584960 617628
rect 579981 617536 584960 617538
rect 579981 617480 579986 617536
rect 580042 617480 584960 617536
rect 579981 617478 584960 617480
rect 579981 617475 580047 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580257 591018 580323 591021
rect 583520 591018 584960 591108
rect 580257 591016 584960 591018
rect 580257 590960 580262 591016
rect 580318 590960 584960 591016
rect 580257 590958 584960 590960
rect 580257 590955 580323 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3693 580002 3759 580005
rect -960 580000 3759 580002
rect -960 579944 3698 580000
rect 3754 579944 3759 580000
rect -960 579942 3759 579944
rect -960 579852 480 579942
rect 3693 579939 3759 579942
rect 580625 577690 580691 577693
rect 583520 577690 584960 577780
rect 580625 577688 584960 577690
rect 580625 577632 580630 577688
rect 580686 577632 584960 577688
rect 580625 577630 584960 577632
rect 580625 577627 580691 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3325 566946 3391 566949
rect -960 566944 3391 566946
rect -960 566888 3330 566944
rect 3386 566888 3391 566944
rect -960 566886 3391 566888
rect -960 566796 480 566886
rect 3325 566883 3391 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 2773 553890 2839 553893
rect -960 553888 2839 553890
rect -960 553832 2778 553888
rect 2834 553832 2839 553888
rect -960 553830 2839 553832
rect -960 553740 480 553830
rect 2773 553827 2839 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3785 527914 3851 527917
rect -960 527912 3851 527914
rect -960 527856 3790 527912
rect 3846 527856 3851 527912
rect -960 527854 3851 527856
rect -960 527764 480 527854
rect 3785 527851 3851 527854
rect 580809 524514 580875 524517
rect 583520 524514 584960 524604
rect 580809 524512 584960 524514
rect 580809 524456 580814 524512
rect 580870 524456 584960 524512
rect 580809 524454 584960 524456
rect 580809 524451 580875 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 579797 511322 579863 511325
rect 583520 511322 584960 511412
rect 579797 511320 584960 511322
rect 579797 511264 579802 511320
rect 579858 511264 584960 511320
rect 579797 511262 584960 511264
rect 579797 511259 579863 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 2773 501802 2839 501805
rect -960 501800 2839 501802
rect -960 501744 2778 501800
rect 2834 501744 2839 501800
rect -960 501742 2839 501744
rect -960 501652 480 501742
rect 2773 501739 2839 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580717 484666 580783 484669
rect 583520 484666 584960 484756
rect 580717 484664 584960 484666
rect 580717 484608 580722 484664
rect 580778 484608 584960 484664
rect 580717 484606 584960 484608
rect 580717 484603 580783 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3969 475690 4035 475693
rect -960 475688 4035 475690
rect -960 475632 3974 475688
rect 4030 475632 4035 475688
rect -960 475630 4035 475632
rect -960 475540 480 475630
rect 3969 475627 4035 475630
rect 580073 471474 580139 471477
rect 583520 471474 584960 471564
rect 580073 471472 584960 471474
rect 580073 471416 580078 471472
rect 580134 471416 584960 471472
rect 580073 471414 584960 471416
rect 580073 471411 580139 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 579981 458146 580047 458149
rect 583520 458146 584960 458236
rect 579981 458144 584960 458146
rect 579981 458088 579986 458144
rect 580042 458088 584960 458144
rect 579981 458086 584960 458088
rect 579981 458083 580047 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 2773 449578 2839 449581
rect -960 449576 2839 449578
rect -960 449520 2778 449576
rect 2834 449520 2839 449576
rect -960 449518 2839 449520
rect -960 449428 480 449518
rect 2773 449515 2839 449518
rect 579981 444818 580047 444821
rect 583520 444818 584960 444908
rect 579981 444816 584960 444818
rect 579981 444760 579986 444816
rect 580042 444760 584960 444816
rect 579981 444758 584960 444760
rect 579981 444755 580047 444758
rect 583520 444668 584960 444758
rect -960 436508 480 436748
rect 580901 431626 580967 431629
rect 583520 431626 584960 431716
rect 580901 431624 584960 431626
rect 580901 431568 580906 431624
rect 580962 431568 584960 431624
rect 580901 431566 584960 431568
rect 580901 431563 580967 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3877 423602 3943 423605
rect -960 423600 3943 423602
rect -960 423544 3882 423600
rect 3938 423544 3943 423600
rect -960 423542 3943 423544
rect -960 423452 480 423542
rect 3877 423539 3943 423542
rect 396574 418236 396580 418300
rect 396644 418298 396650 418300
rect 583520 418298 584960 418388
rect 396644 418238 584960 418298
rect 396644 418236 396650 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 579981 404970 580047 404973
rect 583520 404970 584960 405060
rect 579981 404968 584960 404970
rect 579981 404912 579986 404968
rect 580042 404912 584960 404968
rect 579981 404910 584960 404912
rect 579981 404907 580047 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 2773 397490 2839 397493
rect -960 397488 2839 397490
rect -960 397432 2778 397488
rect 2834 397432 2839 397488
rect -960 397430 2839 397432
rect -960 397340 480 397430
rect 2773 397427 2839 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 579981 378450 580047 378453
rect 583520 378450 584960 378540
rect 579981 378448 584960 378450
rect 579981 378392 579986 378448
rect 580042 378392 584960 378448
rect 579981 378390 584960 378392
rect 579981 378387 580047 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 4061 371378 4127 371381
rect -960 371376 4127 371378
rect -960 371320 4066 371376
rect 4122 371320 4127 371376
rect -960 371318 4127 371320
rect -960 371228 480 371318
rect 4061 371315 4127 371318
rect 579981 365122 580047 365125
rect 583520 365122 584960 365212
rect 579981 365120 584960 365122
rect 579981 365064 579986 365120
rect 580042 365064 584960 365120
rect 579981 365062 584960 365064
rect 579981 365059 580047 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 579981 351930 580047 351933
rect 583520 351930 584960 352020
rect 579981 351928 584960 351930
rect 579981 351872 579986 351928
rect 580042 351872 584960 351928
rect 579981 351870 584960 351872
rect 579981 351867 580047 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 2773 345402 2839 345405
rect -960 345400 2839 345402
rect -960 345344 2778 345400
rect 2834 345344 2839 345400
rect -960 345342 2839 345344
rect -960 345252 480 345342
rect 2773 345339 2839 345342
rect 579981 338602 580047 338605
rect 583520 338602 584960 338692
rect 579981 338600 584960 338602
rect 579981 338544 579986 338600
rect 580042 338544 584960 338600
rect 579981 338542 584960 338544
rect 579981 338539 580047 338542
rect 583520 338452 584960 338542
rect -960 332196 480 332436
rect 579797 325274 579863 325277
rect 583520 325274 584960 325364
rect 579797 325272 584960 325274
rect 579797 325216 579802 325272
rect 579858 325216 584960 325272
rect 579797 325214 584960 325216
rect 579797 325211 579863 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 579981 298754 580047 298757
rect 583520 298754 584960 298844
rect 579981 298752 584960 298754
rect 579981 298696 579986 298752
rect 580042 298696 584960 298752
rect 579981 298694 584960 298696
rect 579981 298691 580047 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3233 293178 3299 293181
rect -960 293176 3299 293178
rect -960 293120 3238 293176
rect 3294 293120 3299 293176
rect -960 293118 3299 293120
rect -960 293028 480 293118
rect 3233 293115 3299 293118
rect 579981 285426 580047 285429
rect 583520 285426 584960 285516
rect 579981 285424 584960 285426
rect 579981 285368 579986 285424
rect 580042 285368 584960 285424
rect 579981 285366 584960 285368
rect 579981 285363 580047 285366
rect 583520 285276 584960 285366
rect -960 279972 480 280212
rect 579981 272234 580047 272237
rect 583520 272234 584960 272324
rect 579981 272232 584960 272234
rect 579981 272176 579986 272232
rect 580042 272176 584960 272232
rect 579981 272174 584960 272176
rect 579981 272171 580047 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3233 267202 3299 267205
rect -960 267200 3299 267202
rect -960 267144 3238 267200
rect 3294 267144 3299 267200
rect -960 267142 3299 267144
rect -960 267052 480 267142
rect 3233 267139 3299 267142
rect 579981 258906 580047 258909
rect 583520 258906 584960 258996
rect 579981 258904 584960 258906
rect 579981 258848 579986 258904
rect 580042 258848 584960 258904
rect 579981 258846 584960 258848
rect 579981 258843 580047 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 579981 245578 580047 245581
rect 583520 245578 584960 245668
rect 579981 245576 584960 245578
rect 579981 245520 579986 245576
rect 580042 245520 584960 245576
rect 579981 245518 584960 245520
rect 579981 245515 580047 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3049 241090 3115 241093
rect -960 241088 3115 241090
rect -960 241032 3054 241088
rect 3110 241032 3115 241088
rect -960 241030 3115 241032
rect -960 240940 480 241030
rect 3049 241027 3115 241030
rect 395337 240138 395403 240141
rect 396758 240138 396764 240140
rect 395337 240136 396764 240138
rect 395337 240080 395342 240136
rect 395398 240080 396764 240136
rect 395337 240078 396764 240080
rect 395337 240075 395403 240078
rect 396758 240076 396764 240078
rect 396828 240076 396834 240140
rect 395521 240002 395587 240005
rect 396942 240002 396948 240004
rect 395521 240000 396948 240002
rect 395521 239944 395526 240000
rect 395582 239944 396948 240000
rect 395521 239942 396948 239944
rect 395521 239939 395587 239942
rect 396942 239940 396948 239942
rect 397012 239940 397018 240004
rect 392577 232386 392643 232389
rect 396758 232386 396764 232388
rect 392577 232384 396764 232386
rect 392577 232328 392582 232384
rect 392638 232328 396764 232384
rect 392577 232326 396764 232328
rect 392577 232323 392643 232326
rect 396758 232324 396764 232326
rect 396828 232324 396834 232388
rect 579797 232386 579863 232389
rect 583520 232386 584960 232476
rect 579797 232384 584960 232386
rect 579797 232328 579802 232384
rect 579858 232328 584960 232384
rect 579797 232326 584960 232328
rect 579797 232323 579863 232326
rect 583520 232236 584960 232326
rect 380157 231162 380223 231165
rect 396942 231162 396948 231164
rect 380157 231160 396948 231162
rect 380157 231104 380162 231160
rect 380218 231104 396948 231160
rect 380157 231102 396948 231104
rect 380157 231099 380223 231102
rect 396942 231100 396948 231102
rect 397012 231100 397018 231164
rect -960 227884 480 228124
rect 579797 219058 579863 219061
rect 583520 219058 584960 219148
rect 579797 219056 584960 219058
rect 579797 219000 579802 219056
rect 579858 219000 584960 219056
rect 579797 218998 584960 219000
rect 579797 218995 579863 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3141 214978 3207 214981
rect -960 214976 3207 214978
rect -960 214920 3146 214976
rect 3202 214920 3207 214976
rect -960 214918 3207 214920
rect -960 214828 480 214918
rect 3141 214915 3207 214918
rect 579981 205730 580047 205733
rect 583520 205730 584960 205820
rect 579981 205728 584960 205730
rect 579981 205672 579986 205728
rect 580042 205672 584960 205728
rect 579981 205670 584960 205672
rect 579981 205667 580047 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 2957 201922 3023 201925
rect -960 201920 3023 201922
rect -960 201864 2962 201920
rect 3018 201864 3023 201920
rect -960 201862 3023 201864
rect -960 201772 480 201862
rect 2957 201859 3023 201862
rect 138105 195938 138171 195941
rect 140405 195938 140471 195941
rect 138105 195936 140471 195938
rect 138105 195880 138110 195936
rect 138166 195880 140410 195936
rect 140466 195880 140471 195936
rect 138105 195878 140471 195880
rect 138105 195875 138171 195878
rect 140405 195875 140471 195878
rect 141417 195938 141483 195941
rect 160829 195938 160895 195941
rect 141417 195936 144194 195938
rect 141417 195880 141422 195936
rect 141478 195880 144194 195936
rect 141417 195878 144194 195880
rect 141417 195875 141483 195878
rect 144134 195644 144194 195878
rect 158854 195936 160895 195938
rect 158854 195928 160834 195936
rect 158854 195872 158902 195928
rect 158958 195880 160834 195928
rect 160890 195880 160895 195936
rect 158958 195878 160895 195880
rect 158958 195872 158963 195878
rect 160829 195875 160895 195878
rect 158854 195870 158963 195872
rect 158897 195867 158963 195870
rect 157149 195666 157215 195669
rect 155910 195664 157215 195666
rect 155910 195608 157154 195664
rect 157210 195608 157215 195664
rect 155910 195606 157215 195608
rect 139393 195530 139459 195533
rect 139393 195528 142170 195530
rect 139393 195472 139398 195528
rect 139454 195498 142170 195528
rect 139454 195472 142692 195498
rect 139393 195470 142692 195472
rect 139393 195467 139459 195470
rect 142110 195438 142692 195470
rect 155910 195340 155970 195606
rect 157149 195603 157215 195606
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 140865 191858 140931 191861
rect 143214 191858 143980 191900
rect 140865 191856 143980 191858
rect 140865 191800 140870 191856
rect 140926 191840 143980 191856
rect 140926 191800 143274 191840
rect 140865 191798 143274 191800
rect 140865 191795 140931 191798
rect 140957 191722 141023 191725
rect 143398 191722 143980 191760
rect 140957 191720 143980 191722
rect 140957 191664 140962 191720
rect 141018 191700 143980 191720
rect 141018 191664 143458 191700
rect 140957 191662 143458 191664
rect 140957 191659 141023 191662
rect 143574 191568 143580 191632
rect 143644 191630 143650 191632
rect 143644 191570 144164 191630
rect 143644 191568 143650 191570
rect 140773 190906 140839 190909
rect 144134 190906 144194 191460
rect 144545 191042 144611 191045
rect 144678 191042 144684 191044
rect 144545 191040 144684 191042
rect 144545 190984 144550 191040
rect 144606 190984 144684 191040
rect 144545 190982 144684 190984
rect 144545 190979 144611 190982
rect 144678 190980 144684 190982
rect 144748 190980 144754 191044
rect 140773 190904 144194 190906
rect 140773 190848 140778 190904
rect 140834 190848 144194 190904
rect 140773 190846 144194 190848
rect 140773 190843 140839 190846
rect 144453 190636 144519 190637
rect 144453 190632 144500 190636
rect 144564 190634 144570 190636
rect 144453 190576 144458 190632
rect 144453 190572 144500 190576
rect 144564 190574 144610 190634
rect 144564 190572 144570 190574
rect 144453 190571 144519 190572
rect 145833 189820 145899 189821
rect 145782 189818 145788 189820
rect 145742 189758 145788 189818
rect 145852 189816 145899 189820
rect 145894 189760 145899 189816
rect 145782 189756 145788 189758
rect 145852 189756 145899 189760
rect 145833 189755 145899 189756
rect -960 188866 480 188956
rect 3141 188866 3207 188869
rect -960 188864 3207 188866
rect -960 188808 3146 188864
rect 3202 188808 3207 188864
rect -960 188806 3207 188808
rect -960 188716 480 188806
rect 3141 188803 3207 188806
rect 140957 184378 141023 184381
rect 143022 184378 143028 184380
rect 140957 184376 143028 184378
rect 140957 184320 140962 184376
rect 141018 184320 143028 184376
rect 140957 184318 143028 184320
rect 140957 184315 141023 184318
rect 143022 184316 143028 184318
rect 143092 184316 143098 184380
rect 140865 184242 140931 184245
rect 141366 184242 141372 184244
rect 140865 184240 141372 184242
rect 140865 184184 140870 184240
rect 140926 184184 141372 184240
rect 140865 184182 141372 184184
rect 140865 184179 140931 184182
rect 141366 184180 141372 184182
rect 141436 184180 141442 184244
rect 144494 183772 144500 183836
rect 144564 183834 144570 183836
rect 144729 183834 144795 183837
rect 144564 183832 144795 183834
rect 144564 183776 144734 183832
rect 144790 183776 144795 183832
rect 144564 183774 144795 183776
rect 144564 183772 144570 183774
rect 144729 183771 144795 183774
rect 144637 183700 144703 183701
rect 144637 183698 144684 183700
rect 144592 183696 144684 183698
rect 144592 183640 144642 183696
rect 144592 183638 144684 183640
rect 144637 183636 144684 183638
rect 144748 183636 144754 183700
rect 144637 183635 144703 183636
rect 140630 182548 140636 182612
rect 140700 182610 140706 182612
rect 140773 182610 140839 182613
rect 140700 182608 140839 182610
rect 140700 182552 140778 182608
rect 140834 182552 140839 182608
rect 140700 182550 140839 182552
rect 140700 182548 140706 182550
rect 140773 182547 140839 182550
rect 145189 181250 145255 181253
rect 145966 181250 145972 181252
rect 145189 181248 145972 181250
rect 145189 181192 145194 181248
rect 145250 181192 145972 181248
rect 145189 181190 145972 181192
rect 145189 181187 145255 181190
rect 145966 181188 145972 181190
rect 146036 181188 146042 181252
rect 143390 180916 143396 180980
rect 143460 180978 143466 180980
rect 144637 180978 144703 180981
rect 143460 180976 144703 180978
rect 143460 180920 144642 180976
rect 144698 180920 144703 180976
rect 143460 180918 144703 180920
rect 143460 180916 143466 180918
rect 144637 180915 144703 180918
rect 157793 179618 157859 179621
rect 158529 179618 158595 179621
rect 157793 179616 158595 179618
rect 157793 179560 157798 179616
rect 157854 179560 158534 179616
rect 158590 179560 158595 179616
rect 157793 179558 158595 179560
rect 157793 179555 157859 179558
rect 158529 179555 158595 179558
rect 149329 179482 149395 179485
rect 149010 179480 149395 179482
rect 149010 179424 149334 179480
rect 149390 179424 149395 179480
rect 149010 179422 149395 179424
rect 148041 179346 148107 179349
rect 149010 179346 149070 179422
rect 149329 179419 149395 179422
rect 148041 179344 149070 179346
rect 148041 179288 148046 179344
rect 148102 179288 149070 179344
rect 148041 179286 149070 179288
rect 148041 179283 148107 179286
rect 579981 179210 580047 179213
rect 583520 179210 584960 179300
rect 579981 179208 584960 179210
rect 579981 179152 579986 179208
rect 580042 179152 584960 179208
rect 579981 179150 584960 179152
rect 579981 179147 580047 179150
rect 142286 179012 142292 179076
rect 142356 179074 142362 179076
rect 142661 179074 142727 179077
rect 142356 179072 142727 179074
rect 142356 179016 142666 179072
rect 142722 179016 142727 179072
rect 583520 179060 584960 179150
rect 142356 179014 142727 179016
rect 142356 179012 142362 179014
rect 142661 179011 142727 179014
rect 143022 178876 143028 178940
rect 143092 178938 143098 178940
rect 144085 178938 144151 178941
rect 143092 178936 144151 178938
rect 143092 178880 144090 178936
rect 144146 178880 144151 178936
rect 143092 178878 144151 178880
rect 143092 178876 143098 178878
rect 144085 178875 144151 178878
rect 141366 178740 141372 178804
rect 141436 178802 141442 178804
rect 141601 178802 141667 178805
rect 141436 178800 141667 178802
rect 141436 178744 141606 178800
rect 141662 178744 141667 178800
rect 141436 178742 141667 178744
rect 141436 178740 141442 178742
rect 141601 178739 141667 178742
rect 157793 178122 157859 178125
rect 158529 178122 158595 178125
rect 157793 178120 158595 178122
rect 157793 178064 157798 178120
rect 157854 178064 158534 178120
rect 158590 178064 158595 178120
rect 157793 178062 158595 178064
rect 157793 178059 157859 178062
rect 158529 178059 158595 178062
rect -960 175796 480 176036
rect 140497 175674 140563 175677
rect 140630 175674 140636 175676
rect 140497 175672 140636 175674
rect 140497 175616 140502 175672
rect 140558 175616 140636 175672
rect 140497 175614 140636 175616
rect 140497 175611 140563 175614
rect 140630 175612 140636 175614
rect 140700 175612 140706 175676
rect 149329 175402 149395 175405
rect 154573 175402 154639 175405
rect 149329 175400 154639 175402
rect 149329 175344 149334 175400
rect 149390 175344 154578 175400
rect 154634 175344 154639 175400
rect 149329 175342 154639 175344
rect 149329 175339 149395 175342
rect 154573 175339 154639 175342
rect 145966 174116 145972 174180
rect 146036 174178 146042 174180
rect 147489 174178 147555 174181
rect 146036 174176 147555 174178
rect 146036 174120 147494 174176
rect 147550 174120 147555 174176
rect 146036 174118 147555 174120
rect 146036 174116 146042 174118
rect 147489 174115 147555 174118
rect 579797 165882 579863 165885
rect 583520 165882 584960 165972
rect 579797 165880 584960 165882
rect 579797 165824 579802 165880
rect 579858 165824 584960 165880
rect 579797 165822 584960 165824
rect 579797 165819 579863 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3141 162890 3207 162893
rect -960 162888 3207 162890
rect -960 162832 3146 162888
rect 3202 162832 3207 162888
rect -960 162830 3207 162832
rect -960 162740 480 162830
rect 3141 162827 3207 162830
rect 580441 152690 580507 152693
rect 583520 152690 584960 152780
rect 580441 152688 584960 152690
rect 580441 152632 580446 152688
rect 580502 152632 584960 152688
rect 580441 152630 584960 152632
rect 580441 152627 580507 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3141 149834 3207 149837
rect -960 149832 3207 149834
rect -960 149776 3146 149832
rect 3202 149776 3207 149832
rect -960 149774 3207 149776
rect -960 149684 480 149774
rect 3141 149771 3207 149774
rect 579981 139362 580047 139365
rect 583520 139362 584960 139452
rect 579981 139360 584960 139362
rect 579981 139304 579986 139360
rect 580042 139304 584960 139360
rect 579981 139302 584960 139304
rect 579981 139299 580047 139302
rect 583520 139212 584960 139302
rect 143574 138756 143580 138820
rect 143644 138818 143650 138820
rect 161565 138818 161631 138821
rect 143644 138816 161631 138818
rect 143644 138760 161570 138816
rect 161626 138760 161631 138816
rect 143644 138758 161631 138760
rect 143644 138756 143650 138758
rect 161565 138755 161631 138758
rect 114001 138682 114067 138685
rect 396574 138682 396580 138684
rect 114001 138680 396580 138682
rect 114001 138624 114006 138680
rect 114062 138624 396580 138680
rect 114001 138622 396580 138624
rect 114001 138619 114067 138622
rect 396574 138620 396580 138622
rect 396644 138620 396650 138684
rect 139669 138002 139735 138005
rect 141918 138002 141924 138004
rect 139669 138000 141924 138002
rect 139669 137944 139674 138000
rect 139730 137944 141924 138000
rect 139669 137942 141924 137944
rect 139669 137939 139735 137942
rect 141918 137940 141924 137942
rect 141988 137940 141994 138004
rect 146150 137532 146156 137596
rect 146220 137594 146226 137596
rect 167821 137594 167887 137597
rect 146220 137592 167887 137594
rect 146220 137536 167826 137592
rect 167882 137536 167887 137592
rect 146220 137534 167887 137536
rect 146220 137532 146226 137534
rect 167821 137531 167887 137534
rect 143390 137396 143396 137460
rect 143460 137458 143466 137460
rect 169385 137458 169451 137461
rect 143460 137456 169451 137458
rect 143460 137400 169390 137456
rect 169446 137400 169451 137456
rect 143460 137398 169451 137400
rect 143460 137396 143466 137398
rect 169385 137395 169451 137398
rect 115289 137322 115355 137325
rect 542670 137322 542676 137324
rect 115289 137320 542676 137322
rect 115289 137264 115294 137320
rect 115350 137264 542676 137320
rect 115289 137262 542676 137264
rect 115289 137259 115355 137262
rect 542670 137260 542676 137262
rect 542740 137260 542746 137324
rect -960 136778 480 136868
rect 3417 136778 3483 136781
rect -960 136776 3483 136778
rect -960 136720 3422 136776
rect 3478 136720 3483 136776
rect -960 136718 3483 136720
rect -960 136628 480 136718
rect 3417 136715 3483 136718
rect 115565 133242 115631 133245
rect 115565 133240 116226 133242
rect 115565 133184 115570 133240
rect 115626 133184 116226 133240
rect 115565 133182 116226 133184
rect 115565 133179 115631 133182
rect 116166 132600 116226 133182
rect 175457 132426 175523 132429
rect 175598 132426 175658 132600
rect 175457 132424 175658 132426
rect 175457 132368 175462 132424
rect 175518 132368 175658 132424
rect 175457 132366 175658 132368
rect 175457 132363 175523 132366
rect 113633 131202 113699 131205
rect 178861 131202 178927 131205
rect 113633 131200 116226 131202
rect 113633 131144 113638 131200
rect 113694 131144 116226 131200
rect 113633 131142 116226 131144
rect 113633 131139 113699 131142
rect 116166 131104 116226 131142
rect 175782 131200 178927 131202
rect 175782 131144 178866 131200
rect 178922 131144 178927 131200
rect 175782 131142 178927 131144
rect 175782 131104 175842 131142
rect 178861 131139 178927 131142
rect 175365 130114 175431 130117
rect 175365 130112 175474 130114
rect 175365 130056 175370 130112
rect 175426 130056 175474 130112
rect 175365 130051 175474 130056
rect 175414 129608 175474 130051
rect 113541 129026 113607 129029
rect 116166 129026 116226 129608
rect 113541 129024 116226 129026
rect 113541 128968 113546 129024
rect 113602 128968 116226 129024
rect 113541 128966 116226 128968
rect 113541 128963 113607 128966
rect 175549 128346 175615 128349
rect 175549 128344 175658 128346
rect 175549 128288 175554 128344
rect 175610 128288 175658 128344
rect 175549 128283 175658 128288
rect 175598 128112 175658 128283
rect 113541 127530 113607 127533
rect 116166 127530 116226 128112
rect 113541 127528 116226 127530
rect 113541 127472 113546 127528
rect 113602 127472 116226 127528
rect 113541 127470 116226 127472
rect 113541 127467 113607 127470
rect 176745 126986 176811 126989
rect 175782 126984 176811 126986
rect 175782 126928 176750 126984
rect 176806 126928 176811 126984
rect 175782 126926 176811 126928
rect 113633 126850 113699 126853
rect 113633 126848 116226 126850
rect 113633 126792 113638 126848
rect 113694 126792 116226 126848
rect 113633 126790 116226 126792
rect 113633 126787 113699 126790
rect 116166 126616 116226 126790
rect 175782 126616 175842 126926
rect 176745 126923 176811 126926
rect 580073 126034 580139 126037
rect 583520 126034 584960 126124
rect 580073 126032 584960 126034
rect 580073 125976 580078 126032
rect 580134 125976 584960 126032
rect 580073 125974 584960 125976
rect 580073 125971 580139 125974
rect 583520 125884 584960 125974
rect 113633 125490 113699 125493
rect 178033 125490 178099 125493
rect 113633 125488 116226 125490
rect 113633 125432 113638 125488
rect 113694 125432 116226 125488
rect 113633 125430 116226 125432
rect 113633 125427 113699 125430
rect 116166 125120 116226 125430
rect 175782 125488 178099 125490
rect 175782 125432 178038 125488
rect 178094 125432 178099 125488
rect 175782 125430 178099 125432
rect 175782 125120 175842 125430
rect 178033 125427 178099 125430
rect 178493 124130 178559 124133
rect 175782 124128 178559 124130
rect 175782 124072 178498 124128
rect 178554 124072 178559 124128
rect 175782 124070 178559 124072
rect 113633 123858 113699 123861
rect 113633 123856 116226 123858
rect -960 123572 480 123812
rect 113633 123800 113638 123856
rect 113694 123800 116226 123856
rect 113633 123798 116226 123800
rect 113633 123795 113699 123798
rect 116166 123624 116226 123798
rect 175782 123624 175842 124070
rect 178493 124067 178559 124070
rect 113633 122770 113699 122773
rect 113633 122768 116226 122770
rect 113633 122712 113638 122768
rect 113694 122712 116226 122768
rect 113633 122710 116226 122712
rect 113633 122707 113699 122710
rect 116166 122128 116226 122710
rect 178125 122498 178191 122501
rect 175782 122496 178191 122498
rect 175782 122440 178130 122496
rect 178186 122440 178191 122496
rect 175782 122438 178191 122440
rect 175782 122128 175842 122438
rect 178125 122435 178191 122438
rect 113633 121274 113699 121277
rect 178401 121274 178467 121277
rect 113633 121272 116226 121274
rect 113633 121216 113638 121272
rect 113694 121216 116226 121272
rect 113633 121214 116226 121216
rect 113633 121211 113699 121214
rect 116166 120632 116226 121214
rect 175782 121272 178467 121274
rect 175782 121216 178406 121272
rect 178462 121216 178467 121272
rect 175782 121214 178467 121216
rect 175782 120632 175842 121214
rect 178401 121211 178467 121214
rect 113633 119778 113699 119781
rect 176653 119778 176719 119781
rect 113633 119776 116226 119778
rect 113633 119720 113638 119776
rect 113694 119720 116226 119776
rect 113633 119718 116226 119720
rect 113633 119715 113699 119718
rect 116166 119136 116226 119718
rect 175782 119776 176719 119778
rect 175782 119720 176658 119776
rect 176714 119720 176719 119776
rect 175782 119718 176719 119720
rect 175782 119136 175842 119718
rect 176653 119715 176719 119718
rect 113633 118282 113699 118285
rect 178585 118282 178651 118285
rect 113633 118280 116226 118282
rect 113633 118224 113638 118280
rect 113694 118224 116226 118280
rect 113633 118222 116226 118224
rect 113633 118219 113699 118222
rect 116166 117640 116226 118222
rect 175782 118280 178651 118282
rect 175782 118224 178590 118280
rect 178646 118224 178651 118280
rect 175782 118222 178651 118224
rect 175782 117640 175842 118222
rect 178585 118219 178651 118222
rect 113633 116786 113699 116789
rect 178769 116786 178835 116789
rect 113633 116784 116226 116786
rect 113633 116728 113638 116784
rect 113694 116728 116226 116784
rect 113633 116726 116226 116728
rect 113633 116723 113699 116726
rect 116166 116144 116226 116726
rect 175782 116784 178835 116786
rect 175782 116728 178774 116784
rect 178830 116728 178835 116784
rect 175782 116726 178835 116728
rect 175782 116144 175842 116726
rect 178769 116723 178835 116726
rect 113541 115290 113607 115293
rect 178309 115290 178375 115293
rect 113541 115288 116226 115290
rect 113541 115232 113546 115288
rect 113602 115232 116226 115288
rect 113541 115230 116226 115232
rect 113541 115227 113607 115230
rect 116166 114648 116226 115230
rect 175782 115288 178375 115290
rect 175782 115232 178314 115288
rect 178370 115232 178375 115288
rect 175782 115230 178375 115232
rect 175782 114648 175842 115230
rect 178309 115227 178375 115230
rect 113633 113114 113699 113117
rect 116166 113114 116226 113152
rect 113633 113112 116226 113114
rect 113633 113056 113638 113112
rect 113694 113056 116226 113112
rect 113633 113054 116226 113056
rect 175782 113114 175842 113152
rect 178677 113114 178743 113117
rect 175782 113112 178743 113114
rect 175782 113056 178682 113112
rect 178738 113056 178743 113112
rect 175782 113054 178743 113056
rect 113633 113051 113699 113054
rect 178677 113051 178743 113054
rect 580533 112842 580599 112845
rect 583520 112842 584960 112932
rect 580533 112840 584960 112842
rect 580533 112784 580538 112840
rect 580594 112784 584960 112840
rect 580533 112782 584960 112784
rect 580533 112779 580599 112782
rect 583520 112692 584960 112782
rect 113633 111754 113699 111757
rect 176837 111754 176903 111757
rect 113633 111752 116226 111754
rect 113633 111696 113638 111752
rect 113694 111696 116226 111752
rect 113633 111694 116226 111696
rect 113633 111691 113699 111694
rect 116166 111656 116226 111694
rect 175782 111752 176903 111754
rect 175782 111696 176842 111752
rect 176898 111696 176903 111752
rect 175782 111694 176903 111696
rect 175782 111656 175842 111694
rect 176837 111691 176903 111694
rect -960 110666 480 110756
rect 3785 110666 3851 110669
rect -960 110664 3851 110666
rect -960 110608 3790 110664
rect 3846 110608 3851 110664
rect -960 110606 3851 110608
rect -960 110516 480 110606
rect 3785 110603 3851 110606
rect 113633 110394 113699 110397
rect 176653 110394 176719 110397
rect 113633 110392 116226 110394
rect 113633 110336 113638 110392
rect 113694 110336 116226 110392
rect 113633 110334 116226 110336
rect 113633 110331 113699 110334
rect 116166 110160 116226 110334
rect 175782 110392 176719 110394
rect 175782 110336 176658 110392
rect 176714 110336 176719 110392
rect 175782 110334 176719 110336
rect 175782 110160 175842 110334
rect 176653 110331 176719 110334
rect 175917 109034 175983 109037
rect 175782 109032 175983 109034
rect 175782 108976 175922 109032
rect 175978 108976 175983 109032
rect 175782 108974 175983 108976
rect 113633 108898 113699 108901
rect 113633 108896 116226 108898
rect 113633 108840 113638 108896
rect 113694 108840 116226 108896
rect 113633 108838 116226 108840
rect 113633 108835 113699 108838
rect 116166 108664 116226 108838
rect 175782 108664 175842 108974
rect 175917 108971 175983 108974
rect 113633 107538 113699 107541
rect 178217 107538 178283 107541
rect 113633 107536 116226 107538
rect 113633 107480 113638 107536
rect 113694 107480 116226 107536
rect 113633 107478 116226 107480
rect 113633 107475 113699 107478
rect 116166 107168 116226 107478
rect 175782 107536 178283 107538
rect 175782 107480 178222 107536
rect 178278 107480 178283 107536
rect 175782 107478 178283 107480
rect 175782 107168 175842 107478
rect 178217 107475 178283 107478
rect 178033 106042 178099 106045
rect 175782 106040 178099 106042
rect 175782 105984 178038 106040
rect 178094 105984 178099 106040
rect 175782 105982 178099 105984
rect 113541 105906 113607 105909
rect 113541 105904 116226 105906
rect 113541 105848 113546 105904
rect 113602 105848 116226 105904
rect 113541 105846 116226 105848
rect 113541 105843 113607 105846
rect 116166 105672 116226 105846
rect 175782 105672 175842 105982
rect 178033 105979 178099 105982
rect 113633 104818 113699 104821
rect 113633 104816 116226 104818
rect 113633 104760 113638 104816
rect 113694 104760 116226 104816
rect 113633 104758 116226 104760
rect 113633 104755 113699 104758
rect 116166 104176 116226 104758
rect 178033 104546 178099 104549
rect 175782 104544 178099 104546
rect 175782 104488 178038 104544
rect 178094 104488 178099 104544
rect 175782 104486 178099 104488
rect 175782 104176 175842 104486
rect 178033 104483 178099 104486
rect 113725 103186 113791 103189
rect 113725 103184 116226 103186
rect 113725 103128 113730 103184
rect 113786 103128 116226 103184
rect 113725 103126 116226 103128
rect 113725 103123 113791 103126
rect 116166 102680 116226 103126
rect 178033 103050 178099 103053
rect 175782 103048 178099 103050
rect 175782 102992 178038 103048
rect 178094 102992 178099 103048
rect 175782 102990 178099 102992
rect 175782 102680 175842 102990
rect 178033 102987 178099 102990
rect 113817 101826 113883 101829
rect 113817 101824 116226 101826
rect 113817 101768 113822 101824
rect 113878 101768 116226 101824
rect 113817 101766 116226 101768
rect 113817 101763 113883 101766
rect 116166 101184 116226 101766
rect 178033 101690 178099 101693
rect 175782 101688 178099 101690
rect 175782 101632 178038 101688
rect 178094 101632 178099 101688
rect 175782 101630 178099 101632
rect 175782 101184 175842 101630
rect 178033 101627 178099 101630
rect 115289 100330 115355 100333
rect 115289 100328 116226 100330
rect 115289 100272 115294 100328
rect 115350 100272 116226 100328
rect 115289 100270 116226 100272
rect 115289 100267 115355 100270
rect 116166 99688 116226 100270
rect 178033 100194 178099 100197
rect 175782 100192 178099 100194
rect 175782 100136 178038 100192
rect 178094 100136 178099 100192
rect 175782 100134 178099 100136
rect 175782 99688 175842 100134
rect 178033 100131 178099 100134
rect 580073 99514 580139 99517
rect 583520 99514 584960 99604
rect 580073 99512 584960 99514
rect 580073 99456 580078 99512
rect 580134 99456 584960 99512
rect 580073 99454 584960 99456
rect 580073 99451 580139 99454
rect 583520 99364 584960 99454
rect 115381 98834 115447 98837
rect 178033 98834 178099 98837
rect 115381 98832 116226 98834
rect 115381 98776 115386 98832
rect 115442 98776 116226 98832
rect 115381 98774 116226 98776
rect 115381 98771 115447 98774
rect 116166 98192 116226 98774
rect 175782 98832 178099 98834
rect 175782 98776 178038 98832
rect 178094 98776 178099 98832
rect 175782 98774 178099 98776
rect 175782 98192 175842 98774
rect 178033 98771 178099 98774
rect -960 97610 480 97700
rect 3693 97610 3759 97613
rect -960 97608 3759 97610
rect -960 97552 3698 97608
rect 3754 97552 3759 97608
rect -960 97550 3759 97552
rect -960 97460 480 97550
rect 3693 97547 3759 97550
rect 178033 97338 178099 97341
rect 175782 97336 178099 97338
rect 175782 97280 178038 97336
rect 178094 97280 178099 97336
rect 175782 97278 178099 97280
rect 115749 96726 115815 96729
rect 115749 96724 116196 96726
rect 115749 96668 115754 96724
rect 115810 96668 116196 96724
rect 175782 96696 175842 97278
rect 178033 97275 178099 97278
rect 115749 96666 116196 96668
rect 115749 96663 115815 96666
rect 115657 95230 115723 95233
rect 115657 95228 116196 95230
rect 115657 95172 115662 95228
rect 115718 95172 116196 95228
rect 115657 95170 116196 95172
rect 115657 95167 115723 95170
rect 175782 95162 175842 95200
rect 178033 95162 178099 95165
rect 175782 95160 178099 95162
rect 175782 95104 178038 95160
rect 178094 95104 178099 95160
rect 175782 95102 178099 95104
rect 178033 95099 178099 95102
rect 115473 93802 115539 93805
rect 178033 93802 178099 93805
rect 115473 93800 116226 93802
rect 115473 93744 115478 93800
rect 115534 93744 116226 93800
rect 115473 93742 116226 93744
rect 115473 93739 115539 93742
rect 116166 93704 116226 93742
rect 175782 93800 178099 93802
rect 175782 93744 178038 93800
rect 178094 93744 178099 93800
rect 175782 93742 178099 93744
rect 175782 93704 175842 93742
rect 178033 93739 178099 93742
rect 115565 92442 115631 92445
rect 115565 92440 116226 92442
rect 115565 92384 115570 92440
rect 115626 92384 116226 92440
rect 115565 92382 116226 92384
rect 115565 92379 115631 92382
rect 116166 92208 116226 92382
rect 178033 92306 178099 92309
rect 175782 92304 178099 92306
rect 175782 92248 178038 92304
rect 178094 92248 178099 92304
rect 175782 92246 178099 92248
rect 175782 92208 175842 92246
rect 178033 92243 178099 92246
rect 113909 91082 113975 91085
rect 113909 91080 116226 91082
rect 113909 91024 113914 91080
rect 113970 91024 116226 91080
rect 113909 91022 116226 91024
rect 113909 91019 113975 91022
rect 116166 90712 116226 91022
rect 178033 90946 178099 90949
rect 175782 90944 178099 90946
rect 175782 90888 178038 90944
rect 178094 90888 178099 90944
rect 175782 90886 178099 90888
rect 175782 90712 175842 90886
rect 178033 90883 178099 90886
rect 114001 89722 114067 89725
rect 114001 89720 116226 89722
rect 114001 89664 114006 89720
rect 114062 89664 116226 89720
rect 114001 89662 116226 89664
rect 114001 89659 114067 89662
rect 116166 89216 116226 89662
rect 178033 89450 178099 89453
rect 175782 89448 178099 89450
rect 175782 89392 178038 89448
rect 178094 89392 178099 89448
rect 175782 89390 178099 89392
rect 175782 89216 175842 89390
rect 178033 89387 178099 89390
rect 114093 88226 114159 88229
rect 114093 88224 116226 88226
rect 114093 88168 114098 88224
rect 114154 88168 116226 88224
rect 114093 88166 116226 88168
rect 114093 88163 114159 88166
rect 116166 87720 116226 88166
rect 178033 88090 178099 88093
rect 175782 88088 178099 88090
rect 175782 88032 178038 88088
rect 178094 88032 178099 88088
rect 175782 88030 178099 88032
rect 175782 87720 175842 88030
rect 178033 88027 178099 88030
rect 114185 86866 114251 86869
rect 114185 86864 116226 86866
rect 114185 86808 114190 86864
rect 114246 86808 116226 86864
rect 114185 86806 116226 86808
rect 114185 86803 114251 86806
rect 116166 86224 116226 86806
rect 178033 86594 178099 86597
rect 175782 86592 178099 86594
rect 175782 86536 178038 86592
rect 178094 86536 178099 86592
rect 175782 86534 178099 86536
rect 175782 86224 175842 86534
rect 178033 86531 178099 86534
rect 580073 86186 580139 86189
rect 583520 86186 584960 86276
rect 580073 86184 584960 86186
rect 580073 86128 580078 86184
rect 580134 86128 584960 86184
rect 580073 86126 584960 86128
rect 580073 86123 580139 86126
rect 583520 86036 584960 86126
rect 114277 85370 114343 85373
rect 114277 85368 116226 85370
rect 114277 85312 114282 85368
rect 114338 85312 116226 85368
rect 114277 85310 116226 85312
rect 114277 85307 114343 85310
rect -960 84690 480 84780
rect 116166 84728 116226 85310
rect 178033 85098 178099 85101
rect 175782 85096 178099 85098
rect 175782 85040 178038 85096
rect 178094 85040 178099 85096
rect 175782 85038 178099 85040
rect 175782 84728 175842 85038
rect 178033 85035 178099 85038
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 178033 83738 178099 83741
rect 175782 83736 178099 83738
rect 175782 83680 178038 83736
rect 178094 83680 178099 83736
rect 175782 83678 178099 83680
rect 115841 83262 115907 83265
rect 115841 83260 116196 83262
rect 115841 83204 115846 83260
rect 115902 83204 116196 83260
rect 175782 83232 175842 83678
rect 178033 83675 178099 83678
rect 115841 83202 116196 83204
rect 115841 83199 115907 83202
rect 114461 82378 114527 82381
rect 114461 82376 116226 82378
rect 114461 82320 114466 82376
rect 114522 82320 116226 82376
rect 114461 82318 116226 82320
rect 114461 82315 114527 82318
rect 116166 81736 116226 82318
rect 178033 82242 178099 82245
rect 175782 82240 178099 82242
rect 175782 82184 178038 82240
rect 178094 82184 178099 82240
rect 175782 82182 178099 82184
rect 175782 81736 175842 82182
rect 178033 82179 178099 82182
rect 114369 80882 114435 80885
rect 179229 80882 179295 80885
rect 114369 80880 116226 80882
rect 114369 80824 114374 80880
rect 114430 80824 116226 80880
rect 114369 80822 116226 80824
rect 114369 80819 114435 80822
rect 116166 80240 116226 80822
rect 175782 80880 179295 80882
rect 175782 80824 179234 80880
rect 179290 80824 179295 80880
rect 175782 80822 179295 80824
rect 175782 80240 175842 80822
rect 179229 80819 179295 80822
rect 114461 78706 114527 78709
rect 116166 78706 116226 78744
rect 114461 78704 116226 78706
rect 114461 78648 114466 78704
rect 114522 78648 116226 78704
rect 114461 78646 116226 78648
rect 175782 78706 175842 78744
rect 178677 78706 178743 78709
rect 175782 78704 178743 78706
rect 175782 78648 178682 78704
rect 178738 78648 178743 78704
rect 175782 78646 178743 78648
rect 114461 78643 114527 78646
rect 178677 78643 178743 78646
rect 114369 76666 114435 76669
rect 116166 76666 116226 77248
rect 114369 76664 116226 76666
rect 114369 76608 114374 76664
rect 114430 76608 116226 76664
rect 114369 76606 116226 76608
rect 175782 76666 175842 77248
rect 178033 76666 178099 76669
rect 175782 76664 178099 76666
rect 175782 76608 178038 76664
rect 178094 76608 178099 76664
rect 175782 76606 178099 76608
rect 114369 76603 114435 76606
rect 178033 76603 178099 76606
rect 114461 75442 114527 75445
rect 116166 75442 116226 75752
rect 114461 75440 116226 75442
rect 114461 75384 114466 75440
rect 114522 75384 116226 75440
rect 114461 75382 116226 75384
rect 114461 75379 114527 75382
rect 5165 75306 5231 75309
rect 169518 75306 169524 75308
rect 5165 75304 169524 75306
rect 5165 75248 5170 75304
rect 5226 75248 169524 75304
rect 5165 75246 169524 75248
rect 5165 75243 5231 75246
rect 169518 75244 169524 75246
rect 169588 75244 169594 75308
rect 4889 75170 4955 75173
rect 4889 75168 167010 75170
rect 4889 75112 4894 75168
rect 4950 75112 167010 75168
rect 4889 75110 167010 75112
rect 4889 75107 4955 75110
rect 166950 75034 167010 75110
rect 167862 75108 167868 75172
rect 167932 75170 167938 75172
rect 172789 75170 172855 75173
rect 167932 75168 172855 75170
rect 167932 75112 172794 75168
rect 172850 75112 172855 75168
rect 167932 75110 172855 75112
rect 167932 75108 167938 75110
rect 172789 75107 172855 75110
rect 527173 75034 527239 75037
rect 166950 74974 168114 75034
rect 167494 74898 167500 74900
rect 157290 74838 167500 74898
rect 156137 74626 156203 74629
rect 157290 74626 157350 74838
rect 167494 74836 167500 74838
rect 167564 74836 167570 74900
rect 167729 74898 167795 74901
rect 167862 74898 167868 74900
rect 167729 74896 167868 74898
rect 167729 74840 167734 74896
rect 167790 74840 167868 74896
rect 167729 74838 167868 74840
rect 167729 74835 167795 74838
rect 167862 74836 167868 74838
rect 167932 74836 167938 74900
rect 161657 74764 161723 74765
rect 161606 74762 161612 74764
rect 161566 74702 161612 74762
rect 161676 74760 161723 74764
rect 164233 74762 164299 74765
rect 161718 74704 161723 74760
rect 161606 74700 161612 74702
rect 161676 74700 161723 74704
rect 161657 74699 161723 74700
rect 164190 74760 164299 74762
rect 164190 74704 164238 74760
rect 164294 74704 164299 74760
rect 164190 74699 164299 74704
rect 164693 74764 164759 74765
rect 164693 74760 164740 74764
rect 164804 74762 164810 74764
rect 168054 74762 168114 74974
rect 172470 75032 527239 75034
rect 172470 74976 527178 75032
rect 527234 74976 527239 75032
rect 172470 74974 527239 74976
rect 168281 74898 168347 74901
rect 172470 74898 172530 74974
rect 527173 74971 527239 74974
rect 168281 74896 172530 74898
rect 168281 74840 168286 74896
rect 168342 74840 172530 74896
rect 168281 74838 172530 74840
rect 172605 74898 172671 74901
rect 580206 74898 580212 74900
rect 172605 74896 580212 74898
rect 172605 74840 172610 74896
rect 172666 74840 580212 74896
rect 172605 74838 580212 74840
rect 168281 74835 168347 74838
rect 172605 74835 172671 74838
rect 580206 74836 580212 74838
rect 580276 74836 580282 74900
rect 169385 74762 169451 74765
rect 169569 74764 169635 74765
rect 164693 74704 164698 74760
rect 164693 74700 164740 74704
rect 164804 74702 164850 74762
rect 168054 74760 169451 74762
rect 168054 74704 169390 74760
rect 169446 74704 169451 74760
rect 168054 74702 169451 74704
rect 164804 74700 164810 74702
rect 164693 74699 164759 74700
rect 169385 74699 169451 74702
rect 169518 74700 169524 74764
rect 169588 74762 169635 74764
rect 172329 74762 172395 74765
rect 580349 74762 580415 74765
rect 169588 74760 169680 74762
rect 169630 74704 169680 74760
rect 169588 74702 169680 74704
rect 172329 74760 580415 74762
rect 172329 74704 172334 74760
rect 172390 74704 580354 74760
rect 580410 74704 580415 74760
rect 172329 74702 580415 74704
rect 169588 74700 169635 74702
rect 169569 74699 169635 74700
rect 172329 74699 172395 74702
rect 580349 74699 580415 74702
rect 156137 74624 157350 74626
rect 156137 74568 156142 74624
rect 156198 74568 157350 74624
rect 156137 74566 157350 74568
rect 156137 74563 156203 74566
rect 164190 74493 164250 74699
rect 168189 74626 168255 74629
rect 172605 74626 172671 74629
rect 168189 74624 172671 74626
rect 168189 74568 168194 74624
rect 168250 74568 172610 74624
rect 172666 74568 172671 74624
rect 168189 74566 172671 74568
rect 168189 74563 168255 74566
rect 172605 74563 172671 74566
rect 172789 74626 172855 74629
rect 580901 74626 580967 74629
rect 172789 74624 580967 74626
rect 172789 74568 172794 74624
rect 172850 74568 580906 74624
rect 580962 74568 580967 74624
rect 172789 74566 580967 74568
rect 172789 74563 172855 74566
rect 580901 74563 580967 74566
rect 154757 74490 154823 74493
rect 161657 74490 161723 74493
rect 154757 74488 161723 74490
rect 154757 74432 154762 74488
rect 154818 74432 161662 74488
rect 161718 74432 161723 74488
rect 154757 74430 161723 74432
rect 164190 74488 164299 74493
rect 164190 74432 164238 74488
rect 164294 74432 164299 74488
rect 164190 74430 164299 74432
rect 154757 74427 154823 74430
rect 161657 74427 161723 74430
rect 164233 74427 164299 74430
rect 167269 74490 167335 74493
rect 580165 74490 580231 74493
rect 167269 74488 580231 74490
rect 167269 74432 167274 74488
rect 167330 74432 580170 74488
rect 580226 74432 580231 74488
rect 167269 74430 580231 74432
rect 167269 74427 167335 74430
rect 580165 74427 580231 74430
rect 167361 74354 167427 74357
rect 520917 74354 520983 74357
rect 167361 74352 520983 74354
rect 167361 74296 167366 74352
rect 167422 74296 520922 74352
rect 520978 74296 520983 74352
rect 167361 74294 520983 74296
rect 167361 74291 167427 74294
rect 520917 74291 520983 74294
rect 161657 74218 161723 74221
rect 164417 74218 164483 74221
rect 161657 74216 164483 74218
rect 161657 74160 161662 74216
rect 161718 74160 164422 74216
rect 164478 74160 164483 74216
rect 161657 74158 164483 74160
rect 161657 74155 161723 74158
rect 164417 74155 164483 74158
rect 164877 74220 164943 74221
rect 164877 74216 164924 74220
rect 164988 74218 164994 74220
rect 167453 74218 167519 74221
rect 396993 74218 397059 74221
rect 164877 74160 164882 74216
rect 164877 74156 164924 74160
rect 164988 74158 165034 74218
rect 167453 74216 397059 74218
rect 167453 74160 167458 74216
rect 167514 74160 396998 74216
rect 397054 74160 397059 74216
rect 167453 74158 397059 74160
rect 164988 74156 164994 74158
rect 164877 74155 164943 74156
rect 167453 74155 167519 74158
rect 396993 74155 397059 74158
rect 4981 74082 5047 74085
rect 167453 74082 167519 74085
rect 170857 74082 170923 74085
rect 4981 74080 167010 74082
rect 4981 74024 4986 74080
rect 5042 74024 167010 74080
rect 4981 74022 167010 74024
rect 4981 74019 5047 74022
rect 3366 73884 3372 73948
rect 3436 73946 3442 73948
rect 166950 73946 167010 74022
rect 167453 74080 170923 74082
rect 167453 74024 167458 74080
rect 167514 74024 170862 74080
rect 170918 74024 170923 74080
rect 167453 74022 170923 74024
rect 167453 74019 167519 74022
rect 170857 74019 170923 74022
rect 169477 73946 169543 73949
rect 3436 73886 162226 73946
rect 166950 73944 169543 73946
rect 166950 73888 169482 73944
rect 169538 73888 169543 73944
rect 166950 73886 169543 73888
rect 3436 73884 3442 73886
rect 3509 73810 3575 73813
rect 162166 73810 162226 73886
rect 169477 73883 169543 73886
rect 169109 73810 169175 73813
rect 3509 73808 162042 73810
rect 3509 73752 3514 73808
rect 3570 73752 162042 73808
rect 3509 73750 162042 73752
rect 162166 73808 169175 73810
rect 162166 73752 169114 73808
rect 169170 73752 169175 73808
rect 162166 73750 169175 73752
rect 3509 73747 3575 73750
rect 4797 73674 4863 73677
rect 161982 73674 162042 73750
rect 169109 73747 169175 73750
rect 169385 73810 169451 73813
rect 172329 73810 172395 73813
rect 169385 73808 172395 73810
rect 169385 73752 169390 73808
rect 169446 73752 172334 73808
rect 172390 73752 172395 73808
rect 169385 73750 172395 73752
rect 169385 73747 169451 73750
rect 172329 73747 172395 73750
rect 169201 73674 169267 73677
rect 4797 73672 157350 73674
rect 4797 73616 4802 73672
rect 4858 73616 157350 73672
rect 4797 73614 157350 73616
rect 161982 73672 169267 73674
rect 161982 73616 169206 73672
rect 169262 73616 169267 73672
rect 161982 73614 169267 73616
rect 4797 73611 4863 73614
rect 157290 73538 157350 73614
rect 169201 73611 169267 73614
rect 169293 73538 169359 73541
rect 157290 73536 169359 73538
rect 157290 73480 169298 73536
rect 169354 73480 169359 73536
rect 157290 73478 169359 73480
rect 169293 73475 169359 73478
rect 166809 73404 166875 73405
rect 166758 73402 166764 73404
rect 166718 73342 166764 73402
rect 166828 73400 166875 73404
rect 166870 73344 166875 73400
rect 166758 73340 166764 73342
rect 166828 73340 166875 73344
rect 166809 73339 166875 73340
rect 161062 73206 167516 73266
rect 128537 73132 128603 73133
rect 128486 73130 128492 73132
rect 128446 73070 128492 73130
rect 128556 73128 128603 73132
rect 128598 73072 128603 73128
rect 128486 73068 128492 73070
rect 128556 73068 128603 73072
rect 128537 73067 128603 73068
rect 158805 73130 158871 73133
rect 161062 73130 161122 73206
rect 158805 73128 161122 73130
rect 158805 73072 158810 73128
rect 158866 73072 161122 73128
rect 158805 73070 161122 73072
rect 161289 73130 161355 73133
rect 162393 73130 162459 73133
rect 161289 73128 162459 73130
rect 161289 73072 161294 73128
rect 161350 73072 162398 73128
rect 162454 73072 162459 73128
rect 161289 73070 162459 73072
rect 158805 73067 158871 73070
rect 161289 73067 161355 73070
rect 162393 73067 162459 73070
rect 163037 73130 163103 73133
rect 165838 73130 165844 73132
rect 163037 73128 165844 73130
rect 163037 73072 163042 73128
rect 163098 73072 165844 73128
rect 163037 73070 165844 73072
rect 163037 73067 163103 73070
rect 165838 73068 165844 73070
rect 165908 73068 165914 73132
rect 152406 72932 152412 72996
rect 152476 72994 152482 72996
rect 153101 72994 153167 72997
rect 152476 72992 153167 72994
rect 152476 72936 153106 72992
rect 153162 72936 153167 72992
rect 152476 72934 153167 72936
rect 152476 72932 152482 72934
rect 153101 72931 153167 72934
rect 155493 72994 155559 72997
rect 155493 72992 166780 72994
rect 155493 72936 155498 72992
rect 155554 72936 166780 72992
rect 155493 72934 166780 72936
rect 155493 72931 155559 72934
rect 148358 72796 148364 72860
rect 148428 72858 148434 72860
rect 148869 72858 148935 72861
rect 148428 72856 148935 72858
rect 148428 72800 148874 72856
rect 148930 72800 148935 72856
rect 148428 72798 148935 72800
rect 148428 72796 148434 72798
rect 148869 72795 148935 72798
rect 149646 72796 149652 72860
rect 149716 72858 149722 72860
rect 150341 72858 150407 72861
rect 149716 72856 150407 72858
rect 149716 72800 150346 72856
rect 150402 72800 150407 72856
rect 149716 72798 150407 72800
rect 149716 72796 149722 72798
rect 150341 72795 150407 72798
rect 151302 72796 151308 72860
rect 151372 72858 151378 72860
rect 151629 72858 151695 72861
rect 151372 72856 151695 72858
rect 151372 72800 151634 72856
rect 151690 72800 151695 72856
rect 151372 72798 151695 72800
rect 151372 72796 151378 72798
rect 151629 72795 151695 72798
rect 152774 72796 152780 72860
rect 152844 72858 152850 72860
rect 152917 72858 152983 72861
rect 152844 72856 152983 72858
rect 152844 72800 152922 72856
rect 152978 72800 152983 72856
rect 152844 72798 152983 72800
rect 152844 72796 152850 72798
rect 152917 72795 152983 72798
rect 154113 72858 154179 72861
rect 156965 72860 157031 72861
rect 154430 72858 154436 72860
rect 154113 72856 154436 72858
rect 154113 72800 154118 72856
rect 154174 72800 154436 72856
rect 154113 72798 154436 72800
rect 154113 72795 154179 72798
rect 154430 72796 154436 72798
rect 154500 72796 154506 72860
rect 156965 72856 157012 72860
rect 157076 72858 157082 72860
rect 158345 72858 158411 72861
rect 158478 72858 158484 72860
rect 156965 72800 156970 72856
rect 156965 72796 157012 72800
rect 157076 72798 157122 72858
rect 158345 72856 158484 72858
rect 158345 72800 158350 72856
rect 158406 72800 158484 72856
rect 158345 72798 158484 72800
rect 157076 72796 157082 72798
rect 156965 72795 157031 72796
rect 158345 72795 158411 72798
rect 158478 72796 158484 72798
rect 158548 72796 158554 72860
rect 158846 72796 158852 72860
rect 158916 72858 158922 72860
rect 159909 72858 159975 72861
rect 158916 72856 159975 72858
rect 158916 72800 159914 72856
rect 159970 72800 159975 72856
rect 158916 72798 159975 72800
rect 158916 72796 158922 72798
rect 159909 72795 159975 72798
rect 160870 72796 160876 72860
rect 160940 72858 160946 72860
rect 161013 72858 161079 72861
rect 160940 72856 161079 72858
rect 160940 72800 161018 72856
rect 161074 72800 161079 72856
rect 160940 72798 161079 72800
rect 160940 72796 160946 72798
rect 161013 72795 161079 72798
rect 162342 72796 162348 72860
rect 162412 72858 162418 72860
rect 162669 72858 162735 72861
rect 162412 72856 162735 72858
rect 162412 72800 162674 72856
rect 162730 72800 162735 72856
rect 162412 72798 162735 72800
rect 162412 72796 162418 72798
rect 162669 72795 162735 72798
rect 163446 72796 163452 72860
rect 163516 72858 163522 72860
rect 163957 72858 164023 72861
rect 164877 72860 164943 72861
rect 165337 72860 165403 72861
rect 164877 72858 164924 72860
rect 163516 72856 164023 72858
rect 163516 72800 163962 72856
rect 164018 72800 164023 72856
rect 163516 72798 164023 72800
rect 164832 72856 164924 72858
rect 164832 72800 164882 72856
rect 164832 72798 164924 72800
rect 163516 72796 163522 72798
rect 163957 72795 164023 72798
rect 164877 72796 164924 72798
rect 164988 72796 164994 72860
rect 165286 72858 165292 72860
rect 165246 72798 165292 72858
rect 165356 72856 165403 72860
rect 165398 72800 165403 72856
rect 165286 72796 165292 72798
rect 165356 72796 165403 72800
rect 164877 72795 164943 72796
rect 165337 72795 165403 72796
rect 166349 72858 166415 72861
rect 166574 72858 166580 72860
rect 166349 72856 166580 72858
rect 166349 72800 166354 72856
rect 166410 72800 166580 72856
rect 166349 72798 166580 72800
rect 166349 72795 166415 72798
rect 166574 72796 166580 72798
rect 166644 72796 166650 72860
rect 166720 72858 166780 72934
rect 167269 72858 167335 72861
rect 166720 72856 167335 72858
rect 166720 72800 167274 72856
rect 167330 72800 167335 72856
rect 166720 72798 167335 72800
rect 167456 72858 167516 73206
rect 168005 73130 168071 73133
rect 580257 73130 580323 73133
rect 168005 73128 580323 73130
rect 168005 73072 168010 73128
rect 168066 73072 580262 73128
rect 580318 73072 580323 73128
rect 168005 73070 580323 73072
rect 168005 73067 168071 73070
rect 580257 73067 580323 73070
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 478873 72858 478939 72861
rect 167456 72856 478939 72858
rect 167456 72800 478878 72856
rect 478934 72800 478939 72856
rect 583520 72844 584960 72934
rect 167456 72798 478939 72800
rect 167269 72795 167335 72798
rect 478873 72795 478939 72798
rect 148685 72724 148751 72725
rect 148961 72724 149027 72725
rect 148685 72720 148732 72724
rect 148796 72722 148802 72724
rect 148685 72664 148690 72720
rect 148685 72660 148732 72664
rect 148796 72662 148842 72722
rect 148796 72660 148802 72662
rect 148910 72660 148916 72724
rect 148980 72722 149027 72724
rect 149973 72724 150039 72725
rect 148980 72720 149072 72722
rect 149022 72664 149072 72720
rect 148980 72662 149072 72664
rect 149973 72720 150020 72724
rect 150084 72722 150090 72724
rect 151537 72722 151603 72725
rect 153009 72724 153075 72725
rect 151670 72722 151676 72724
rect 149973 72664 149978 72720
rect 148980 72660 149027 72662
rect 148685 72659 148751 72660
rect 148961 72659 149027 72660
rect 149973 72660 150020 72664
rect 150084 72662 150130 72722
rect 151537 72720 151676 72722
rect 151537 72664 151542 72720
rect 151598 72664 151676 72720
rect 151537 72662 151676 72664
rect 150084 72660 150090 72662
rect 149973 72659 150039 72660
rect 151537 72659 151603 72662
rect 151670 72660 151676 72662
rect 151740 72660 151746 72724
rect 152958 72722 152964 72724
rect 152918 72662 152964 72722
rect 153028 72720 153075 72724
rect 153070 72664 153075 72720
rect 152958 72660 152964 72662
rect 153028 72660 153075 72664
rect 153009 72659 153075 72660
rect 154205 72724 154271 72725
rect 154205 72720 154252 72724
rect 154316 72722 154322 72724
rect 154205 72664 154210 72720
rect 154205 72660 154252 72664
rect 154316 72662 154362 72722
rect 154316 72660 154322 72662
rect 155718 72660 155724 72724
rect 155788 72722 155794 72724
rect 155861 72722 155927 72725
rect 156873 72724 156939 72725
rect 157241 72724 157307 72725
rect 156822 72722 156828 72724
rect 155788 72720 155927 72722
rect 155788 72664 155866 72720
rect 155922 72664 155927 72720
rect 155788 72662 155927 72664
rect 156782 72662 156828 72722
rect 156892 72720 156939 72724
rect 157190 72722 157196 72724
rect 156934 72664 156939 72720
rect 155788 72660 155794 72662
rect 154205 72659 154271 72660
rect 155861 72659 155927 72662
rect 156822 72660 156828 72662
rect 156892 72660 156939 72664
rect 157150 72662 157196 72722
rect 157260 72720 157307 72724
rect 157302 72664 157307 72720
rect 157190 72660 157196 72662
rect 157260 72660 157307 72664
rect 156873 72659 156939 72660
rect 157241 72659 157307 72660
rect 158529 72722 158595 72725
rect 158662 72722 158668 72724
rect 158529 72720 158668 72722
rect 158529 72664 158534 72720
rect 158590 72664 158668 72720
rect 158529 72662 158668 72664
rect 158529 72659 158595 72662
rect 158662 72660 158668 72662
rect 158732 72660 158738 72724
rect 159030 72660 159036 72724
rect 159100 72722 159106 72724
rect 160001 72722 160067 72725
rect 161105 72724 161171 72725
rect 161054 72722 161060 72724
rect 159100 72720 160067 72722
rect 159100 72664 160006 72720
rect 160062 72664 160067 72720
rect 159100 72662 160067 72664
rect 161014 72662 161060 72722
rect 161124 72720 161171 72724
rect 161166 72664 161171 72720
rect 159100 72660 159106 72662
rect 160001 72659 160067 72662
rect 161054 72660 161060 72662
rect 161124 72660 161171 72664
rect 161238 72660 161244 72724
rect 161308 72722 161314 72724
rect 161381 72722 161447 72725
rect 161308 72720 161447 72722
rect 161308 72664 161386 72720
rect 161442 72664 161447 72720
rect 161308 72662 161447 72664
rect 161308 72660 161314 72662
rect 161105 72659 161171 72660
rect 161381 72659 161447 72662
rect 162485 72724 162551 72725
rect 162761 72724 162827 72725
rect 162485 72720 162532 72724
rect 162596 72722 162602 72724
rect 162485 72664 162490 72720
rect 162485 72660 162532 72664
rect 162596 72662 162642 72722
rect 162596 72660 162602 72662
rect 162710 72660 162716 72724
rect 162780 72722 162827 72724
rect 162780 72720 162872 72722
rect 162822 72664 162872 72720
rect 162780 72662 162872 72664
rect 162780 72660 162827 72662
rect 163630 72660 163636 72724
rect 163700 72722 163706 72724
rect 164141 72722 164207 72725
rect 163700 72720 164207 72722
rect 163700 72664 164146 72720
rect 164202 72664 164207 72720
rect 163700 72662 164207 72664
rect 163700 72660 163706 72662
rect 162485 72659 162551 72660
rect 162761 72659 162827 72660
rect 164141 72659 164207 72662
rect 164918 72660 164924 72724
rect 164988 72722 164994 72724
rect 165245 72722 165311 72725
rect 165521 72724 165587 72725
rect 165470 72722 165476 72724
rect 164988 72720 165311 72722
rect 164988 72664 165250 72720
rect 165306 72664 165311 72720
rect 164988 72662 165311 72664
rect 165430 72662 165476 72722
rect 165540 72720 165587 72724
rect 165582 72664 165587 72720
rect 164988 72660 164994 72662
rect 165245 72659 165311 72662
rect 165470 72660 165476 72662
rect 165540 72660 165587 72664
rect 166390 72660 166396 72724
rect 166460 72722 166466 72724
rect 166533 72722 166599 72725
rect 166460 72720 166599 72722
rect 166460 72664 166538 72720
rect 166594 72664 166599 72720
rect 166460 72662 166599 72664
rect 166460 72660 166466 72662
rect 165521 72659 165587 72660
rect 166533 72659 166599 72662
rect 168557 72722 168623 72725
rect 480253 72722 480319 72725
rect 168557 72720 480319 72722
rect 168557 72664 168562 72720
rect 168618 72664 480258 72720
rect 480314 72664 480319 72720
rect 168557 72662 480319 72664
rect 168557 72659 168623 72662
rect 480253 72659 480319 72662
rect 22737 72586 22803 72589
rect 121913 72586 121979 72589
rect 22737 72584 121979 72586
rect 22737 72528 22742 72584
rect 22798 72528 121918 72584
rect 121974 72528 121979 72584
rect 22737 72526 121979 72528
rect 22737 72523 22803 72526
rect 121913 72523 121979 72526
rect 149462 72524 149468 72588
rect 149532 72586 149538 72588
rect 150157 72586 150223 72589
rect 149532 72584 150223 72586
rect 149532 72528 150162 72584
rect 150218 72528 150223 72584
rect 149532 72526 150223 72528
rect 149532 72524 149538 72526
rect 150157 72523 150223 72526
rect 152590 72524 152596 72588
rect 152660 72586 152666 72588
rect 152825 72586 152891 72589
rect 152660 72584 152891 72586
rect 152660 72528 152830 72584
rect 152886 72528 152891 72584
rect 152660 72526 152891 72528
rect 152660 72524 152666 72526
rect 152825 72523 152891 72526
rect 153878 72524 153884 72588
rect 153948 72586 153954 72588
rect 154481 72586 154547 72589
rect 153948 72584 154547 72586
rect 153948 72528 154486 72584
rect 154542 72528 154547 72584
rect 153948 72526 154547 72528
rect 153948 72524 153954 72526
rect 154481 72523 154547 72526
rect 156638 72524 156644 72588
rect 156708 72586 156714 72588
rect 157057 72586 157123 72589
rect 156708 72584 157123 72586
rect 156708 72528 157062 72584
rect 157118 72528 157123 72584
rect 156708 72526 157123 72528
rect 156708 72524 156714 72526
rect 157057 72523 157123 72526
rect 158294 72524 158300 72588
rect 158364 72586 158370 72588
rect 158621 72586 158687 72589
rect 158364 72584 158687 72586
rect 158364 72528 158626 72584
rect 158682 72528 158687 72584
rect 158364 72526 158687 72528
rect 158364 72524 158370 72526
rect 158621 72523 158687 72526
rect 160686 72524 160692 72588
rect 160756 72586 160762 72588
rect 161197 72586 161263 72589
rect 160756 72584 161263 72586
rect 160756 72528 161202 72584
rect 161258 72528 161263 72584
rect 160756 72526 161263 72528
rect 160756 72524 160762 72526
rect 161197 72523 161263 72526
rect 161606 72524 161612 72588
rect 161676 72586 161682 72588
rect 162485 72586 162551 72589
rect 161676 72584 162551 72586
rect 161676 72528 162490 72584
rect 162546 72528 162551 72584
rect 161676 72526 162551 72528
rect 161676 72524 161682 72526
rect 162485 72523 162551 72526
rect 163262 72524 163268 72588
rect 163332 72586 163338 72588
rect 164049 72586 164115 72589
rect 163332 72584 164115 72586
rect 163332 72528 164054 72584
rect 164110 72528 164115 72584
rect 163332 72526 164115 72528
rect 163332 72524 163338 72526
rect 164049 72523 164115 72526
rect 165102 72524 165108 72588
rect 165172 72586 165178 72588
rect 165429 72586 165495 72589
rect 498193 72586 498259 72589
rect 165172 72584 165495 72586
rect 165172 72528 165434 72584
rect 165490 72528 165495 72584
rect 165172 72526 165495 72528
rect 165172 72524 165178 72526
rect 165429 72523 165495 72526
rect 168974 72584 498259 72586
rect 168974 72528 498198 72584
rect 498254 72528 498259 72584
rect 168974 72526 498259 72528
rect 148542 72388 148548 72452
rect 148612 72450 148618 72452
rect 148777 72450 148843 72453
rect 148612 72448 148843 72450
rect 148612 72392 148782 72448
rect 148838 72392 148843 72448
rect 148612 72390 148843 72392
rect 148612 72388 148618 72390
rect 148777 72387 148843 72390
rect 149830 72388 149836 72452
rect 149900 72450 149906 72452
rect 150065 72450 150131 72453
rect 149900 72448 150131 72450
rect 149900 72392 150070 72448
rect 150126 72392 150131 72448
rect 149900 72390 150131 72392
rect 149900 72388 149906 72390
rect 150065 72387 150131 72390
rect 151486 72388 151492 72452
rect 151556 72450 151562 72452
rect 151721 72450 151787 72453
rect 151556 72448 151787 72450
rect 151556 72392 151726 72448
rect 151782 72392 151787 72448
rect 151556 72390 151787 72392
rect 151556 72388 151562 72390
rect 151721 72387 151787 72390
rect 154062 72388 154068 72452
rect 154132 72450 154138 72452
rect 154297 72450 154363 72453
rect 154132 72448 154363 72450
rect 154132 72392 154302 72448
rect 154358 72392 154363 72448
rect 154132 72390 154363 72392
rect 154132 72388 154138 72390
rect 154297 72387 154363 72390
rect 155534 72388 155540 72452
rect 155604 72450 155610 72452
rect 155769 72450 155835 72453
rect 155604 72448 155835 72450
rect 155604 72392 155774 72448
rect 155830 72392 155835 72448
rect 155604 72390 155835 72392
rect 155604 72388 155610 72390
rect 155769 72387 155835 72390
rect 158110 72388 158116 72452
rect 158180 72450 158186 72452
rect 158437 72450 158503 72453
rect 158180 72448 158503 72450
rect 158180 72392 158442 72448
rect 158498 72392 158503 72448
rect 158180 72390 158503 72392
rect 158180 72388 158186 72390
rect 158437 72387 158503 72390
rect 159633 72450 159699 72453
rect 161289 72450 161355 72453
rect 159633 72448 161355 72450
rect 159633 72392 159638 72448
rect 159694 72392 161294 72448
rect 161350 72392 161355 72448
rect 159633 72390 161355 72392
rect 159633 72387 159699 72390
rect 161289 72387 161355 72390
rect 162158 72388 162164 72452
rect 162228 72450 162234 72452
rect 162577 72450 162643 72453
rect 162228 72448 162643 72450
rect 162228 72392 162582 72448
rect 162638 72392 162643 72448
rect 162228 72390 162643 72392
rect 162228 72388 162234 72390
rect 162577 72387 162643 72390
rect 163086 72390 166596 72450
rect 125685 72314 125751 72317
rect 126094 72314 126100 72316
rect 125685 72312 126100 72314
rect 125685 72256 125690 72312
rect 125746 72256 126100 72312
rect 125685 72254 126100 72256
rect 125685 72251 125751 72254
rect 126094 72252 126100 72254
rect 126164 72252 126170 72316
rect 146886 72252 146892 72316
rect 146956 72314 146962 72316
rect 147489 72314 147555 72317
rect 146956 72312 147555 72314
rect 146956 72256 147494 72312
rect 147550 72256 147555 72312
rect 146956 72254 147555 72256
rect 146956 72252 146962 72254
rect 147489 72251 147555 72254
rect 155677 72314 155743 72317
rect 157057 72314 157123 72317
rect 155677 72312 157123 72314
rect 155677 72256 155682 72312
rect 155738 72256 157062 72312
rect 157118 72256 157123 72312
rect 155677 72254 157123 72256
rect 155677 72251 155743 72254
rect 157057 72251 157123 72254
rect 160277 72314 160343 72317
rect 163086 72314 163146 72390
rect 160277 72312 163146 72314
rect 160277 72256 160282 72312
rect 160338 72256 163146 72312
rect 160277 72254 163146 72256
rect 163313 72314 163379 72317
rect 165521 72314 165587 72317
rect 163313 72312 165587 72314
rect 163313 72256 163318 72312
rect 163374 72256 165526 72312
rect 165582 72256 165587 72312
rect 163313 72254 165587 72256
rect 166536 72314 166596 72390
rect 168974 72314 169034 72526
rect 498193 72523 498259 72526
rect 172881 72450 172947 72453
rect 581085 72450 581151 72453
rect 172881 72448 581151 72450
rect 172881 72392 172886 72448
rect 172942 72392 581090 72448
rect 581146 72392 581151 72448
rect 172881 72390 581151 72392
rect 172881 72387 172947 72390
rect 581085 72387 581151 72390
rect 166536 72254 169034 72314
rect 160277 72251 160343 72254
rect 163313 72251 163379 72254
rect 165521 72251 165587 72254
rect 124213 72178 124279 72181
rect 124622 72178 124628 72180
rect 124213 72176 124628 72178
rect 124213 72120 124218 72176
rect 124274 72120 124628 72176
rect 124213 72118 124628 72120
rect 124213 72115 124279 72118
rect 124622 72116 124628 72118
rect 124692 72116 124698 72180
rect 125593 72178 125659 72181
rect 125910 72178 125916 72180
rect 125593 72176 125916 72178
rect 125593 72120 125598 72176
rect 125654 72120 125916 72176
rect 125593 72118 125916 72120
rect 125593 72115 125659 72118
rect 125910 72116 125916 72118
rect 125980 72116 125986 72180
rect 128445 72178 128511 72181
rect 129038 72178 129044 72180
rect 128445 72176 129044 72178
rect 128445 72120 128450 72176
rect 128506 72120 129044 72176
rect 128445 72118 129044 72120
rect 128445 72115 128511 72118
rect 129038 72116 129044 72118
rect 129108 72116 129114 72180
rect 129733 72178 129799 72181
rect 129958 72178 129964 72180
rect 129733 72176 129964 72178
rect 129733 72120 129738 72176
rect 129794 72120 129964 72176
rect 129733 72118 129964 72120
rect 129733 72115 129799 72118
rect 129958 72116 129964 72118
rect 130028 72116 130034 72180
rect 133270 72116 133276 72180
rect 133340 72178 133346 72180
rect 133689 72178 133755 72181
rect 133340 72176 133755 72178
rect 133340 72120 133694 72176
rect 133750 72120 133755 72176
rect 133340 72118 133755 72120
rect 133340 72116 133346 72118
rect 133689 72115 133755 72118
rect 134742 72116 134748 72180
rect 134812 72178 134818 72180
rect 135069 72178 135135 72181
rect 134812 72176 135135 72178
rect 134812 72120 135074 72176
rect 135130 72120 135135 72176
rect 134812 72118 135135 72120
rect 134812 72116 134818 72118
rect 135069 72115 135135 72118
rect 135846 72116 135852 72180
rect 135916 72178 135922 72180
rect 136449 72178 136515 72181
rect 135916 72176 136515 72178
rect 135916 72120 136454 72176
rect 136510 72120 136515 72176
rect 135916 72118 136515 72120
rect 135916 72116 135922 72118
rect 136449 72115 136515 72118
rect 138974 72116 138980 72180
rect 139044 72178 139050 72180
rect 139301 72178 139367 72181
rect 139044 72176 139367 72178
rect 139044 72120 139306 72176
rect 139362 72120 139367 72176
rect 139044 72118 139367 72120
rect 139044 72116 139050 72118
rect 139301 72115 139367 72118
rect 140078 72116 140084 72180
rect 140148 72178 140154 72180
rect 140313 72178 140379 72181
rect 140148 72176 140379 72178
rect 140148 72120 140318 72176
rect 140374 72120 140379 72176
rect 140148 72118 140379 72120
rect 140148 72116 140154 72118
rect 140313 72115 140379 72118
rect 142838 72116 142844 72180
rect 142908 72178 142914 72180
rect 143257 72178 143323 72181
rect 142908 72176 143323 72178
rect 142908 72120 143262 72176
rect 143318 72120 143323 72176
rect 142908 72118 143323 72120
rect 142908 72116 142914 72118
rect 143257 72115 143323 72118
rect 144126 72116 144132 72180
rect 144196 72178 144202 72180
rect 144729 72178 144795 72181
rect 144196 72176 144795 72178
rect 144196 72120 144734 72176
rect 144790 72120 144795 72176
rect 144196 72118 144795 72120
rect 144196 72116 144202 72118
rect 144729 72115 144795 72118
rect 145230 72116 145236 72180
rect 145300 72178 145306 72180
rect 146017 72178 146083 72181
rect 145300 72176 146083 72178
rect 145300 72120 146022 72176
rect 146078 72120 146083 72176
rect 145300 72118 146083 72120
rect 145300 72116 145306 72118
rect 146017 72115 146083 72118
rect 147070 72116 147076 72180
rect 147140 72178 147146 72180
rect 147397 72178 147463 72181
rect 147140 72176 147463 72178
rect 147140 72120 147402 72176
rect 147458 72120 147463 72176
rect 147140 72118 147463 72120
rect 147140 72116 147146 72118
rect 147397 72115 147463 72118
rect 158897 72178 158963 72181
rect 168557 72178 168623 72181
rect 158897 72176 168623 72178
rect 158897 72120 158902 72176
rect 158958 72120 168562 72176
rect 168618 72120 168623 72176
rect 158897 72118 168623 72120
rect 158897 72115 158963 72118
rect 168557 72115 168623 72118
rect 121637 72044 121703 72045
rect 122833 72044 122899 72045
rect 121637 72042 121684 72044
rect 121592 72040 121684 72042
rect 121592 71984 121642 72040
rect 121592 71982 121684 71984
rect 121637 71980 121684 71982
rect 121748 71980 121754 72044
rect 122782 71980 122788 72044
rect 122852 72042 122899 72044
rect 122852 72040 122944 72042
rect 122894 71984 122944 72040
rect 122852 71982 122944 71984
rect 122852 71980 122899 71982
rect 124254 71980 124260 72044
rect 124324 72042 124330 72044
rect 124397 72042 124463 72045
rect 124324 72040 124463 72042
rect 124324 71984 124402 72040
rect 124458 71984 124463 72040
rect 124324 71982 124463 71984
rect 124324 71980 124330 71982
rect 121637 71979 121703 71980
rect 122833 71979 122899 71980
rect 124397 71979 124463 71982
rect 125542 71980 125548 72044
rect 125612 72042 125618 72044
rect 125777 72042 125843 72045
rect 125612 72040 125843 72042
rect 125612 71984 125782 72040
rect 125838 71984 125843 72040
rect 125612 71982 125843 71984
rect 125612 71980 125618 71982
rect 125777 71979 125843 71982
rect 127065 72042 127131 72045
rect 127198 72042 127204 72044
rect 127065 72040 127204 72042
rect 127065 71984 127070 72040
rect 127126 71984 127204 72040
rect 127065 71982 127204 71984
rect 127065 71979 127131 71982
rect 127198 71980 127204 71982
rect 127268 71980 127274 72044
rect 128353 72042 128419 72045
rect 128854 72042 128860 72044
rect 128353 72040 128860 72042
rect 128353 71984 128358 72040
rect 128414 71984 128860 72040
rect 128353 71982 128860 71984
rect 128353 71979 128419 71982
rect 128854 71980 128860 71982
rect 128924 71980 128930 72044
rect 130009 72042 130075 72045
rect 130142 72042 130148 72044
rect 130009 72040 130148 72042
rect 130009 71984 130014 72040
rect 130070 71984 130148 72040
rect 130009 71982 130148 71984
rect 130009 71979 130075 71982
rect 130142 71980 130148 71982
rect 130212 71980 130218 72044
rect 131062 71980 131068 72044
rect 131132 72042 131138 72044
rect 131205 72042 131271 72045
rect 131132 72040 131271 72042
rect 131132 71984 131210 72040
rect 131266 71984 131271 72040
rect 131132 71982 131271 71984
rect 131132 71980 131138 71982
rect 131205 71979 131271 71982
rect 131798 71980 131804 72044
rect 131868 72042 131874 72044
rect 132217 72042 132283 72045
rect 131868 72040 132283 72042
rect 131868 71984 132222 72040
rect 132278 71984 132283 72040
rect 131868 71982 132283 71984
rect 131868 71980 131874 71982
rect 132217 71979 132283 71982
rect 133454 71980 133460 72044
rect 133524 72042 133530 72044
rect 133597 72042 133663 72045
rect 134977 72044 135043 72045
rect 134926 72042 134932 72044
rect 133524 72040 133663 72042
rect 133524 71984 133602 72040
rect 133658 71984 133663 72040
rect 133524 71982 133663 71984
rect 134886 71982 134932 72042
rect 134996 72040 135043 72044
rect 135038 71984 135043 72040
rect 133524 71980 133530 71982
rect 133597 71979 133663 71982
rect 134926 71980 134932 71982
rect 134996 71980 135043 71984
rect 136214 71980 136220 72044
rect 136284 72042 136290 72044
rect 136357 72042 136423 72045
rect 136284 72040 136423 72042
rect 136284 71984 136362 72040
rect 136418 71984 136423 72040
rect 136284 71982 136423 71984
rect 136284 71980 136290 71982
rect 134977 71979 135043 71980
rect 136357 71979 136423 71982
rect 137686 71980 137692 72044
rect 137756 72042 137762 72044
rect 137829 72042 137895 72045
rect 137756 72040 137895 72042
rect 137756 71984 137834 72040
rect 137890 71984 137895 72040
rect 137756 71982 137895 71984
rect 137756 71980 137762 71982
rect 137829 71979 137895 71982
rect 138790 71980 138796 72044
rect 138860 72042 138866 72044
rect 139025 72042 139091 72045
rect 138860 72040 139091 72042
rect 138860 71984 139030 72040
rect 139086 71984 139091 72040
rect 138860 71982 139091 71984
rect 138860 71980 138866 71982
rect 139025 71979 139091 71982
rect 140262 71980 140268 72044
rect 140332 72042 140338 72044
rect 140589 72042 140655 72045
rect 140332 72040 140655 72042
rect 140332 71984 140594 72040
rect 140650 71984 140655 72040
rect 140332 71982 140655 71984
rect 140332 71980 140338 71982
rect 140589 71979 140655 71982
rect 140814 71980 140820 72044
rect 140884 72042 140890 72044
rect 141969 72042 142035 72045
rect 140884 72040 142035 72042
rect 140884 71984 141974 72040
rect 142030 71984 142035 72040
rect 140884 71982 142035 71984
rect 140884 71980 140890 71982
rect 141969 71979 142035 71982
rect 143022 71980 143028 72044
rect 143092 72042 143098 72044
rect 143349 72042 143415 72045
rect 143092 72040 143415 72042
rect 143092 71984 143354 72040
rect 143410 71984 143415 72040
rect 143092 71982 143415 71984
rect 143092 71980 143098 71982
rect 143349 71979 143415 71982
rect 144494 71980 144500 72044
rect 144564 72042 144570 72044
rect 144637 72042 144703 72045
rect 144564 72040 144703 72042
rect 144564 71984 144642 72040
rect 144698 71984 144703 72040
rect 144564 71982 144703 71984
rect 144564 71980 144570 71982
rect 144637 71979 144703 71982
rect 145414 71980 145420 72044
rect 145484 72042 145490 72044
rect 146201 72042 146267 72045
rect 145484 72040 146267 72042
rect 145484 71984 146206 72040
rect 146262 71984 146267 72040
rect 145484 71982 146267 71984
rect 145484 71980 145490 71982
rect 146201 71979 146267 71982
rect 147254 71980 147260 72044
rect 147324 72042 147330 72044
rect 147581 72042 147647 72045
rect 147324 72040 147647 72042
rect 147324 71984 147586 72040
rect 147642 71984 147647 72040
rect 147324 71982 147647 71984
rect 147324 71980 147330 71982
rect 147581 71979 147647 71982
rect 157149 72042 157215 72045
rect 157793 72042 157859 72045
rect 157149 72040 157859 72042
rect 157149 71984 157154 72040
rect 157210 71984 157798 72040
rect 157854 71984 157859 72040
rect 157149 71982 157859 71984
rect 157149 71979 157215 71982
rect 157793 71979 157859 71982
rect 121545 71908 121611 71909
rect 121494 71906 121500 71908
rect 121454 71846 121500 71906
rect 121564 71904 121611 71908
rect 122925 71908 122991 71909
rect 124489 71908 124555 71909
rect 122925 71906 122972 71908
rect 121606 71848 121611 71904
rect 121494 71844 121500 71846
rect 121564 71844 121611 71848
rect 122880 71904 122972 71906
rect 122880 71848 122930 71904
rect 122880 71846 122972 71848
rect 121545 71843 121611 71844
rect 122925 71844 122972 71846
rect 123036 71844 123042 71908
rect 124438 71906 124444 71908
rect 124398 71846 124444 71906
rect 124508 71904 124555 71908
rect 124550 71848 124555 71904
rect 124438 71844 124444 71846
rect 124508 71844 124555 71848
rect 125726 71844 125732 71908
rect 125796 71906 125802 71908
rect 125869 71906 125935 71909
rect 126973 71908 127039 71909
rect 128629 71908 128695 71909
rect 126973 71906 127020 71908
rect 125796 71904 125935 71906
rect 125796 71848 125874 71904
rect 125930 71848 125935 71904
rect 125796 71846 125935 71848
rect 126928 71904 127020 71906
rect 126928 71848 126978 71904
rect 126928 71846 127020 71848
rect 125796 71844 125802 71846
rect 122925 71843 122991 71844
rect 124489 71843 124555 71844
rect 125869 71843 125935 71846
rect 126973 71844 127020 71846
rect 127084 71844 127090 71908
rect 128629 71906 128676 71908
rect 128584 71904 128676 71906
rect 128584 71848 128634 71904
rect 128584 71846 128676 71848
rect 128629 71844 128676 71846
rect 128740 71844 128746 71908
rect 129774 71844 129780 71908
rect 129844 71906 129850 71908
rect 129917 71906 129983 71909
rect 129844 71904 129983 71906
rect 129844 71848 129922 71904
rect 129978 71848 129983 71904
rect 129844 71846 129983 71848
rect 129844 71844 129850 71846
rect 126973 71843 127039 71844
rect 128629 71843 128695 71844
rect 129917 71843 129983 71846
rect 131113 71906 131179 71909
rect 131246 71906 131252 71908
rect 131113 71904 131252 71906
rect 131113 71848 131118 71904
rect 131174 71848 131252 71904
rect 131113 71846 131252 71848
rect 131113 71843 131179 71846
rect 131246 71844 131252 71846
rect 131316 71844 131322 71908
rect 131982 71844 131988 71908
rect 132052 71906 132058 71908
rect 132401 71906 132467 71909
rect 132052 71904 132467 71906
rect 132052 71848 132406 71904
rect 132462 71848 132467 71904
rect 132052 71846 132467 71848
rect 132052 71844 132058 71846
rect 132401 71843 132467 71846
rect 133638 71844 133644 71908
rect 133708 71906 133714 71908
rect 133781 71906 133847 71909
rect 135161 71908 135227 71909
rect 135110 71906 135116 71908
rect 133708 71904 133847 71906
rect 133708 71848 133786 71904
rect 133842 71848 133847 71904
rect 133708 71846 133847 71848
rect 135070 71846 135116 71906
rect 135180 71904 135227 71908
rect 135222 71848 135227 71904
rect 133708 71844 133714 71846
rect 133781 71843 133847 71846
rect 135110 71844 135116 71846
rect 135180 71844 135227 71848
rect 136030 71844 136036 71908
rect 136100 71906 136106 71908
rect 136173 71906 136239 71909
rect 136100 71904 136239 71906
rect 136100 71848 136178 71904
rect 136234 71848 136239 71904
rect 136100 71846 136239 71848
rect 136100 71844 136106 71846
rect 135161 71843 135227 71844
rect 136173 71843 136239 71846
rect 136398 71844 136404 71908
rect 136468 71906 136474 71908
rect 136541 71906 136607 71909
rect 137921 71908 137987 71909
rect 137870 71906 137876 71908
rect 136468 71904 136607 71906
rect 136468 71848 136546 71904
rect 136602 71848 136607 71904
rect 136468 71846 136607 71848
rect 137830 71846 137876 71906
rect 137940 71904 137987 71908
rect 137982 71848 137987 71904
rect 136468 71844 136474 71846
rect 136541 71843 136607 71846
rect 137870 71844 137876 71846
rect 137940 71844 137987 71848
rect 138606 71844 138612 71908
rect 138676 71906 138682 71908
rect 138933 71906 138999 71909
rect 139117 71908 139183 71909
rect 140405 71908 140471 71909
rect 140681 71908 140747 71909
rect 139117 71906 139164 71908
rect 138676 71904 138999 71906
rect 138676 71848 138938 71904
rect 138994 71848 138999 71904
rect 138676 71846 138999 71848
rect 139072 71904 139164 71906
rect 139072 71848 139122 71904
rect 139072 71846 139164 71848
rect 138676 71844 138682 71846
rect 137921 71843 137987 71844
rect 138933 71843 138999 71846
rect 139117 71844 139164 71846
rect 139228 71844 139234 71908
rect 140405 71906 140452 71908
rect 140360 71904 140452 71906
rect 140360 71848 140410 71904
rect 140360 71846 140452 71848
rect 140405 71844 140452 71846
rect 140516 71844 140522 71908
rect 140630 71844 140636 71908
rect 140700 71906 140747 71908
rect 140700 71904 140792 71906
rect 140742 71848 140792 71904
rect 140700 71846 140792 71848
rect 140700 71844 140747 71846
rect 140998 71844 141004 71908
rect 141068 71906 141074 71908
rect 142061 71906 142127 71909
rect 143165 71908 143231 71909
rect 143441 71908 143507 71909
rect 143165 71906 143212 71908
rect 141068 71904 142127 71906
rect 141068 71848 142066 71904
rect 142122 71848 142127 71904
rect 141068 71846 142127 71848
rect 143120 71904 143212 71906
rect 143120 71848 143170 71904
rect 143120 71846 143212 71848
rect 141068 71844 141074 71846
rect 139117 71843 139183 71844
rect 140405 71843 140471 71844
rect 140681 71843 140747 71844
rect 142061 71843 142127 71846
rect 143165 71844 143212 71846
rect 143276 71844 143282 71908
rect 143390 71906 143396 71908
rect 143350 71846 143396 71906
rect 143460 71904 143507 71908
rect 143502 71848 143507 71904
rect 143390 71844 143396 71846
rect 143460 71844 143507 71848
rect 144310 71844 144316 71908
rect 144380 71906 144386 71908
rect 144545 71906 144611 71909
rect 144380 71904 144611 71906
rect 144380 71848 144550 71904
rect 144606 71848 144611 71904
rect 144380 71846 144611 71848
rect 144380 71844 144386 71846
rect 143165 71843 143231 71844
rect 143441 71843 143507 71844
rect 144545 71843 144611 71846
rect 144678 71844 144684 71908
rect 144748 71906 144754 71908
rect 144821 71906 144887 71909
rect 144748 71904 144887 71906
rect 144748 71848 144826 71904
rect 144882 71848 144887 71904
rect 144748 71846 144887 71848
rect 144748 71844 144754 71846
rect 144821 71843 144887 71846
rect 145598 71844 145604 71908
rect 145668 71906 145674 71908
rect 146109 71906 146175 71909
rect 145668 71904 146175 71906
rect 145668 71848 146114 71904
rect 146170 71848 146175 71904
rect 145668 71846 146175 71848
rect 145668 71844 145674 71846
rect 146109 71843 146175 71846
rect 147305 71906 147371 71909
rect 147438 71906 147444 71908
rect 147305 71904 147444 71906
rect 147305 71848 147310 71904
rect 147366 71848 147444 71904
rect 147305 71846 147444 71848
rect 147305 71843 147371 71846
rect 147438 71844 147444 71846
rect 147508 71844 147514 71908
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 164693 71364 164759 71365
rect 164693 71362 164740 71364
rect 164648 71360 164740 71362
rect 164648 71304 164698 71360
rect 164648 71302 164740 71304
rect 164693 71300 164740 71302
rect 164804 71300 164810 71364
rect 164693 71299 164759 71300
rect 165838 71164 165844 71228
rect 165908 71226 165914 71228
rect 167862 71226 167868 71228
rect 165908 71166 167868 71226
rect 165908 71164 165914 71166
rect 167862 71164 167868 71166
rect 167932 71164 167938 71228
rect 165521 70138 165587 70141
rect 167678 70138 167684 70140
rect 165521 70136 167684 70138
rect 165521 70080 165526 70136
rect 165582 70080 167684 70136
rect 165521 70078 167684 70080
rect 165521 70075 165587 70078
rect 167678 70076 167684 70078
rect 167748 70076 167754 70140
rect 158662 65452 158668 65516
rect 158732 65514 158738 65516
rect 474733 65514 474799 65517
rect 158732 65512 474799 65514
rect 158732 65456 474738 65512
rect 474794 65456 474799 65512
rect 158732 65454 474799 65456
rect 158732 65452 158738 65454
rect 474733 65451 474799 65454
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3601 58578 3667 58581
rect -960 58576 3667 58578
rect -960 58520 3606 58576
rect 3662 58520 3667 58576
rect -960 58518 3667 58520
rect -960 58428 480 58518
rect 3601 58515 3667 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 144126 35260 144132 35324
rect 144196 35322 144202 35324
rect 298093 35322 298159 35325
rect 144196 35320 298159 35322
rect 144196 35264 298098 35320
rect 298154 35264 298159 35320
rect 144196 35262 298159 35264
rect 144196 35260 144202 35262
rect 298093 35259 298159 35262
rect 146886 35124 146892 35188
rect 146956 35186 146962 35188
rect 332593 35186 332659 35189
rect 146956 35184 332659 35186
rect 146956 35128 332598 35184
rect 332654 35128 332659 35184
rect 146956 35126 332659 35128
rect 146956 35124 146962 35126
rect 332593 35123 332659 35126
rect 137686 34036 137692 34100
rect 137756 34098 137762 34100
rect 209773 34098 209839 34101
rect 137756 34096 209839 34098
rect 137756 34040 209778 34096
rect 209834 34040 209839 34096
rect 137756 34038 209839 34040
rect 137756 34036 137762 34038
rect 209773 34035 209839 34038
rect 140078 33900 140084 33964
rect 140148 33962 140154 33964
rect 241513 33962 241579 33965
rect 140148 33960 241579 33962
rect 140148 33904 241518 33960
rect 241574 33904 241579 33960
rect 140148 33902 241579 33904
rect 140148 33900 140154 33902
rect 241513 33899 241579 33902
rect 140814 33764 140820 33828
rect 140884 33826 140890 33828
rect 262213 33826 262279 33829
rect 140884 33824 262279 33826
rect 140884 33768 262218 33824
rect 262274 33768 262279 33824
rect 140884 33766 262279 33768
rect 140884 33764 140890 33766
rect 262213 33763 262279 33766
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect 134742 32676 134748 32740
rect 134812 32738 134818 32740
rect 173893 32738 173959 32741
rect 134812 32736 173959 32738
rect 134812 32680 173898 32736
rect 173954 32680 173959 32736
rect 134812 32678 173959 32680
rect 134812 32676 134818 32678
rect 173893 32675 173959 32678
rect -960 32466 480 32556
rect 136030 32540 136036 32604
rect 136100 32602 136106 32604
rect 187693 32602 187759 32605
rect 136100 32600 187759 32602
rect 136100 32544 187698 32600
rect 187754 32544 187759 32600
rect 136100 32542 187759 32544
rect 136100 32540 136106 32542
rect 187693 32539 187759 32542
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 135846 32404 135852 32468
rect 135916 32466 135922 32468
rect 191833 32466 191899 32469
rect 135916 32464 191899 32466
rect 135916 32408 191838 32464
rect 191894 32408 191899 32464
rect 135916 32406 191899 32408
rect 135916 32404 135922 32406
rect 191833 32403 191899 32406
rect 163262 31180 163268 31244
rect 163332 31242 163338 31244
rect 445017 31242 445083 31245
rect 163332 31240 445083 31242
rect 163332 31184 445022 31240
rect 445078 31184 445083 31240
rect 163332 31182 445083 31184
rect 163332 31180 163338 31182
rect 445017 31179 445083 31182
rect 158110 31044 158116 31108
rect 158180 31106 158186 31108
rect 473353 31106 473419 31109
rect 158180 31104 473419 31106
rect 158180 31048 473358 31104
rect 473414 31048 473419 31104
rect 158180 31046 473419 31048
rect 158180 31044 158186 31046
rect 473353 31043 473419 31046
rect 158846 30908 158852 30972
rect 158916 30970 158922 30972
rect 492673 30970 492739 30973
rect 158916 30968 492739 30970
rect 158916 30912 492678 30968
rect 492734 30912 492739 30968
rect 158916 30910 492739 30912
rect 158916 30908 158922 30910
rect 492673 30907 492739 30910
rect 145230 29548 145236 29612
rect 145300 29610 145306 29612
rect 314653 29610 314719 29613
rect 145300 29608 314719 29610
rect 145300 29552 314658 29608
rect 314714 29552 314719 29608
rect 145300 29550 314719 29552
rect 145300 29548 145306 29550
rect 314653 29547 314719 29550
rect 136214 27100 136220 27164
rect 136284 27162 136290 27164
rect 190453 27162 190519 27165
rect 136284 27160 190519 27162
rect 136284 27104 190458 27160
rect 190514 27104 190519 27160
rect 136284 27102 190519 27104
rect 136284 27100 136290 27102
rect 190453 27099 190519 27102
rect 142838 26964 142844 27028
rect 142908 27026 142914 27028
rect 278773 27026 278839 27029
rect 142908 27024 278839 27026
rect 142908 26968 278778 27024
rect 278834 26968 278839 27024
rect 142908 26966 278839 26968
rect 142908 26964 142914 26966
rect 278773 26963 278839 26966
rect 149462 26828 149468 26892
rect 149532 26890 149538 26892
rect 367093 26890 367159 26893
rect 149532 26888 367159 26890
rect 149532 26832 367098 26888
rect 367154 26832 367159 26888
rect 149532 26830 367159 26832
rect 149532 26828 149538 26830
rect 367093 26827 367159 26830
rect 134926 25604 134932 25668
rect 134996 25666 135002 25668
rect 172513 25666 172579 25669
rect 134996 25664 172579 25666
rect 134996 25608 172518 25664
rect 172574 25608 172579 25664
rect 134996 25606 172579 25608
rect 134996 25604 135002 25606
rect 172513 25603 172579 25606
rect 156638 25468 156644 25532
rect 156708 25530 156714 25532
rect 456885 25530 456951 25533
rect 156708 25528 456951 25530
rect 156708 25472 456890 25528
rect 456946 25472 456951 25528
rect 156708 25470 456951 25472
rect 156708 25468 156714 25470
rect 456885 25467 456951 25470
rect 151302 24380 151308 24444
rect 151372 24442 151378 24444
rect 386413 24442 386479 24445
rect 151372 24440 386479 24442
rect 151372 24384 386418 24440
rect 386474 24384 386479 24440
rect 151372 24382 386479 24384
rect 151372 24380 151378 24382
rect 386413 24379 386479 24382
rect 162158 24244 162164 24308
rect 162228 24306 162234 24308
rect 527173 24306 527239 24309
rect 162228 24304 527239 24306
rect 162228 24248 527178 24304
rect 527234 24248 527239 24304
rect 162228 24246 527239 24248
rect 162228 24244 162234 24246
rect 527173 24243 527239 24246
rect 163446 24108 163452 24172
rect 163516 24170 163522 24172
rect 545113 24170 545179 24173
rect 163516 24168 545179 24170
rect 163516 24112 545118 24168
rect 545174 24112 545179 24168
rect 163516 24110 545179 24112
rect 163516 24108 163522 24110
rect 545113 24107 545179 24110
rect 155534 22884 155540 22948
rect 155604 22946 155610 22948
rect 440233 22946 440299 22949
rect 155604 22944 440299 22946
rect 155604 22888 440238 22944
rect 440294 22888 440299 22944
rect 155604 22886 440299 22888
rect 155604 22884 155610 22886
rect 440233 22883 440299 22886
rect 156822 22748 156828 22812
rect 156892 22810 156898 22812
rect 454033 22810 454099 22813
rect 156892 22808 454099 22810
rect 156892 22752 454038 22808
rect 454094 22752 454099 22808
rect 156892 22750 454099 22752
rect 156892 22748 156898 22750
rect 454033 22747 454099 22750
rect 160686 22612 160692 22676
rect 160756 22674 160762 22676
rect 509233 22674 509299 22677
rect 160756 22672 509299 22674
rect 160756 22616 509238 22672
rect 509294 22616 509299 22672
rect 160756 22614 509299 22616
rect 160756 22612 160762 22614
rect 509233 22611 509299 22614
rect 148358 21388 148364 21452
rect 148428 21450 148434 21452
rect 350533 21450 350599 21453
rect 148428 21448 350599 21450
rect 148428 21392 350538 21448
rect 350594 21392 350599 21448
rect 148428 21390 350599 21392
rect 148428 21388 148434 21390
rect 350533 21387 350599 21390
rect 158294 21252 158300 21316
rect 158364 21314 158370 21316
rect 476113 21314 476179 21317
rect 158364 21312 476179 21314
rect 158364 21256 476118 21312
rect 476174 21256 476179 21312
rect 158364 21254 476179 21256
rect 158364 21252 158370 21254
rect 476113 21251 476179 21254
rect 138606 20164 138612 20228
rect 138676 20226 138682 20228
rect 223573 20226 223639 20229
rect 138676 20224 223639 20226
rect 138676 20168 223578 20224
rect 223634 20168 223639 20224
rect 138676 20166 223639 20168
rect 138676 20164 138682 20166
rect 223573 20163 223639 20166
rect 140262 20028 140268 20092
rect 140332 20090 140338 20092
rect 244273 20090 244339 20093
rect 140332 20088 244339 20090
rect 140332 20032 244278 20088
rect 244334 20032 244339 20088
rect 140332 20030 244339 20032
rect 140332 20028 140338 20030
rect 244273 20027 244339 20030
rect 158478 19892 158484 19956
rect 158548 19954 158554 19956
rect 473445 19954 473511 19957
rect 158548 19952 473511 19954
rect 158548 19896 473450 19952
rect 473506 19896 473511 19952
rect 158548 19894 473511 19896
rect 158548 19892 158554 19894
rect 473445 19891 473511 19894
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 157006 18804 157012 18868
rect 157076 18866 157082 18868
rect 455413 18866 455479 18869
rect 157076 18864 455479 18866
rect 157076 18808 455418 18864
rect 455474 18808 455479 18864
rect 157076 18806 455479 18808
rect 157076 18804 157082 18806
rect 455413 18803 455479 18806
rect 157190 18668 157196 18732
rect 157260 18730 157266 18732
rect 458173 18730 458239 18733
rect 157260 18728 458239 18730
rect 157260 18672 458178 18728
rect 458234 18672 458239 18728
rect 157260 18670 458239 18672
rect 157260 18668 157266 18670
rect 458173 18667 458239 18670
rect 162342 18532 162348 18596
rect 162412 18594 162418 18596
rect 528553 18594 528619 18597
rect 162412 18592 528619 18594
rect 162412 18536 528558 18592
rect 528614 18536 528619 18592
rect 162412 18534 528619 18536
rect 162412 18532 162418 18534
rect 528553 18531 528619 18534
rect 145414 17580 145420 17644
rect 145484 17642 145490 17644
rect 316033 17642 316099 17645
rect 145484 17640 316099 17642
rect 145484 17584 316038 17640
rect 316094 17584 316099 17640
rect 145484 17582 316099 17584
rect 145484 17580 145490 17582
rect 316033 17579 316099 17582
rect 154062 17444 154068 17508
rect 154132 17506 154138 17508
rect 420913 17506 420979 17509
rect 154132 17504 420979 17506
rect 154132 17448 420918 17504
rect 420974 17448 420979 17504
rect 154132 17446 420979 17448
rect 154132 17444 154138 17446
rect 420913 17443 420979 17446
rect 153878 17308 153884 17372
rect 153948 17370 153954 17372
rect 423765 17370 423831 17373
rect 153948 17368 423831 17370
rect 153948 17312 423770 17368
rect 423826 17312 423831 17368
rect 153948 17310 423831 17312
rect 153948 17308 153954 17310
rect 423765 17307 423831 17310
rect 155718 17172 155724 17236
rect 155788 17234 155794 17236
rect 440325 17234 440391 17237
rect 155788 17232 440391 17234
rect 155788 17176 440330 17232
rect 440386 17176 440391 17232
rect 155788 17174 440391 17176
rect 155788 17172 155794 17174
rect 440325 17171 440391 17174
rect 144310 16220 144316 16284
rect 144380 16282 144386 16284
rect 295609 16282 295675 16285
rect 144380 16280 295675 16282
rect 144380 16224 295614 16280
rect 295670 16224 295675 16280
rect 144380 16222 295675 16224
rect 144380 16220 144386 16222
rect 295609 16219 295675 16222
rect 148542 16084 148548 16148
rect 148612 16146 148618 16148
rect 349153 16146 349219 16149
rect 148612 16144 349219 16146
rect 148612 16088 349158 16144
rect 349214 16088 349219 16144
rect 148612 16086 349219 16088
rect 148612 16084 148618 16086
rect 349153 16083 349219 16086
rect 152406 15948 152412 16012
rect 152476 16010 152482 16012
rect 406009 16010 406075 16013
rect 152476 16008 406075 16010
rect 152476 15952 406014 16008
rect 406070 15952 406075 16008
rect 152476 15950 406075 15952
rect 152476 15948 152482 15950
rect 406009 15947 406075 15950
rect 154246 15812 154252 15876
rect 154316 15874 154322 15876
rect 420177 15874 420243 15877
rect 154316 15872 420243 15874
rect 154316 15816 420182 15872
rect 420238 15816 420243 15872
rect 154316 15814 420243 15816
rect 154316 15812 154322 15814
rect 420177 15811 420243 15814
rect 140998 15132 141004 15196
rect 141068 15194 141074 15196
rect 264145 15194 264211 15197
rect 141068 15192 264211 15194
rect 141068 15136 264150 15192
rect 264206 15136 264211 15192
rect 141068 15134 264211 15136
rect 141068 15132 141074 15134
rect 264145 15131 264211 15134
rect 144494 14996 144500 15060
rect 144564 15058 144570 15060
rect 297265 15058 297331 15061
rect 144564 15056 297331 15058
rect 144564 15000 297270 15056
rect 297326 15000 297331 15056
rect 144564 14998 297331 15000
rect 144564 14996 144570 14998
rect 297265 14995 297331 14998
rect 145598 14860 145604 14924
rect 145668 14922 145674 14924
rect 316217 14922 316283 14925
rect 145668 14920 316283 14922
rect 145668 14864 316222 14920
rect 316278 14864 316283 14920
rect 145668 14862 316283 14864
rect 145668 14860 145674 14862
rect 316217 14859 316283 14862
rect 147070 14724 147076 14788
rect 147140 14786 147146 14788
rect 332685 14786 332751 14789
rect 147140 14784 332751 14786
rect 147140 14728 332690 14784
rect 332746 14728 332751 14784
rect 147140 14726 332751 14728
rect 147140 14724 147146 14726
rect 332685 14723 332751 14726
rect 151486 14588 151492 14652
rect 151556 14650 151562 14652
rect 387793 14650 387859 14653
rect 151556 14648 387859 14650
rect 151556 14592 387798 14648
rect 387854 14592 387859 14648
rect 151556 14590 387859 14592
rect 151556 14588 151562 14590
rect 387793 14587 387859 14590
rect 152590 14452 152596 14516
rect 152660 14514 152666 14516
rect 402513 14514 402579 14517
rect 152660 14512 402579 14514
rect 152660 14456 402518 14512
rect 402574 14456 402579 14512
rect 152660 14454 402579 14456
rect 152660 14452 152666 14454
rect 402513 14451 402579 14454
rect 140446 13636 140452 13700
rect 140516 13698 140522 13700
rect 242985 13698 243051 13701
rect 140516 13696 243051 13698
rect 140516 13640 242990 13696
rect 243046 13640 243051 13696
rect 140516 13638 243051 13640
rect 140516 13636 140522 13638
rect 242985 13635 243051 13638
rect 143022 13500 143028 13564
rect 143092 13562 143098 13564
rect 280705 13562 280771 13565
rect 143092 13560 280771 13562
rect 143092 13504 280710 13560
rect 280766 13504 280771 13560
rect 143092 13502 280771 13504
rect 143092 13500 143098 13502
rect 280705 13499 280771 13502
rect 149830 13364 149836 13428
rect 149900 13426 149906 13428
rect 365713 13426 365779 13429
rect 149900 13424 365779 13426
rect 149900 13368 365718 13424
rect 365774 13368 365779 13424
rect 149900 13366 365779 13368
rect 149900 13364 149906 13366
rect 365713 13363 365779 13366
rect 149646 13228 149652 13292
rect 149716 13290 149722 13292
rect 370129 13290 370195 13293
rect 149716 13288 370195 13290
rect 149716 13232 370134 13288
rect 370190 13232 370195 13288
rect 149716 13230 370195 13232
rect 149716 13228 149722 13230
rect 370129 13227 370195 13230
rect 154430 13092 154436 13156
rect 154500 13154 154506 13156
rect 418521 13154 418587 13157
rect 154500 13152 418587 13154
rect 154500 13096 418526 13152
rect 418582 13096 418587 13152
rect 154500 13094 418587 13096
rect 154500 13092 154506 13094
rect 418521 13091 418587 13094
rect 160870 12956 160876 13020
rect 160940 13018 160946 13020
rect 507209 13018 507275 13021
rect 160940 13016 507275 13018
rect 160940 12960 507214 13016
rect 507270 12960 507275 13016
rect 160940 12958 507275 12960
rect 160940 12956 160946 12958
rect 507209 12955 507275 12958
rect 138790 12820 138796 12884
rect 138860 12882 138866 12884
rect 225137 12882 225203 12885
rect 138860 12880 225203 12882
rect 138860 12824 225142 12880
rect 225198 12824 225203 12880
rect 138860 12822 225203 12824
rect 138860 12820 138866 12822
rect 225137 12819 225203 12822
rect 137870 12140 137876 12204
rect 137940 12202 137946 12204
rect 210969 12202 211035 12205
rect 137940 12200 211035 12202
rect 137940 12144 210974 12200
rect 211030 12144 211035 12200
rect 137940 12142 211035 12144
rect 137940 12140 137946 12142
rect 210969 12139 211035 12142
rect 148726 12004 148732 12068
rect 148796 12066 148802 12068
rect 349245 12066 349311 12069
rect 148796 12064 349311 12066
rect 148796 12008 349250 12064
rect 349306 12008 349311 12064
rect 148796 12006 349311 12008
rect 148796 12004 148802 12006
rect 349245 12003 349311 12006
rect 148910 11868 148916 11932
rect 148980 11930 148986 11932
rect 352833 11930 352899 11933
rect 148980 11928 352899 11930
rect 148980 11872 352838 11928
rect 352894 11872 352899 11928
rect 148980 11870 352899 11872
rect 148980 11868 148986 11870
rect 352833 11867 352899 11870
rect 150014 11732 150020 11796
rect 150084 11794 150090 11796
rect 365805 11794 365871 11797
rect 150084 11792 365871 11794
rect 150084 11736 365810 11792
rect 365866 11736 365871 11792
rect 150084 11734 365871 11736
rect 150084 11732 150090 11734
rect 365805 11731 365871 11734
rect 152774 11596 152780 11660
rect 152844 11658 152850 11660
rect 403617 11658 403683 11661
rect 152844 11656 403683 11658
rect 152844 11600 403622 11656
rect 403678 11600 403683 11656
rect 152844 11598 403683 11600
rect 152844 11596 152850 11598
rect 403617 11595 403683 11598
rect 89161 10434 89227 10437
rect 129038 10434 129044 10436
rect 89161 10432 129044 10434
rect 89161 10376 89166 10432
rect 89222 10376 129044 10432
rect 89161 10374 129044 10376
rect 89161 10371 89227 10374
rect 129038 10372 129044 10374
rect 129108 10372 129114 10436
rect 147438 10372 147444 10436
rect 147508 10434 147514 10436
rect 331213 10434 331279 10437
rect 147508 10432 331279 10434
rect 147508 10376 331218 10432
rect 331274 10376 331279 10432
rect 147508 10374 331279 10376
rect 147508 10372 147514 10374
rect 331213 10371 331279 10374
rect 71497 10298 71563 10301
rect 127198 10298 127204 10300
rect 71497 10296 127204 10298
rect 71497 10240 71502 10296
rect 71558 10240 127204 10296
rect 71497 10238 127204 10240
rect 71497 10235 71563 10238
rect 127198 10236 127204 10238
rect 127268 10236 127274 10300
rect 147254 10236 147260 10300
rect 147324 10298 147330 10300
rect 334617 10298 334683 10301
rect 147324 10296 334683 10298
rect 147324 10240 334622 10296
rect 334678 10240 334683 10296
rect 147324 10238 334683 10240
rect 147324 10236 147330 10238
rect 334617 10235 334683 10238
rect 109309 9482 109375 9485
rect 130142 9482 130148 9484
rect 109309 9480 130148 9482
rect 109309 9424 109314 9480
rect 109370 9424 130148 9480
rect 109309 9422 130148 9424
rect 109309 9419 109375 9422
rect 130142 9420 130148 9422
rect 130212 9420 130218 9484
rect 105721 9346 105787 9349
rect 129958 9346 129964 9348
rect 105721 9344 129964 9346
rect 105721 9288 105726 9344
rect 105782 9288 129964 9344
rect 105721 9286 129964 9288
rect 105721 9283 105787 9286
rect 129958 9284 129964 9286
rect 130028 9284 130034 9348
rect 53741 9210 53807 9213
rect 126094 9210 126100 9212
rect 53741 9208 126100 9210
rect 53741 9152 53746 9208
rect 53802 9152 126100 9208
rect 53741 9150 126100 9152
rect 53741 9147 53807 9150
rect 126094 9148 126100 9150
rect 126164 9148 126170 9212
rect 38377 9074 38443 9077
rect 124438 9074 124444 9076
rect 38377 9072 124444 9074
rect 38377 9016 38382 9072
rect 38438 9016 124444 9072
rect 38377 9014 124444 9016
rect 38377 9011 38443 9014
rect 124438 9012 124444 9014
rect 124508 9012 124514 9076
rect 144678 9012 144684 9076
rect 144748 9074 144754 9076
rect 299657 9074 299723 9077
rect 144748 9072 299723 9074
rect 144748 9016 299662 9072
rect 299718 9016 299723 9072
rect 144748 9014 299723 9016
rect 144748 9012 144754 9014
rect 299657 9011 299723 9014
rect 34789 8938 34855 8941
rect 124622 8938 124628 8940
rect 34789 8936 124628 8938
rect 34789 8880 34794 8936
rect 34850 8880 124628 8936
rect 34789 8878 124628 8880
rect 34789 8875 34855 8878
rect 124622 8876 124628 8878
rect 124692 8876 124698 8940
rect 166390 8876 166396 8940
rect 166460 8938 166466 8940
rect 578601 8938 578667 8941
rect 166460 8936 578667 8938
rect 166460 8880 578606 8936
rect 578662 8880 578667 8936
rect 166460 8878 578667 8880
rect 166460 8876 166466 8878
rect 578601 8875 578667 8878
rect 135110 8060 135116 8124
rect 135180 8122 135186 8124
rect 169661 8122 169727 8125
rect 135180 8120 169727 8122
rect 135180 8064 169666 8120
rect 169722 8064 169727 8120
rect 135180 8062 169727 8064
rect 135180 8060 135186 8062
rect 169661 8059 169727 8062
rect 143206 7924 143212 7988
rect 143276 7986 143282 7988
rect 278313 7986 278379 7989
rect 143276 7984 278379 7986
rect 143276 7928 278318 7984
rect 278374 7928 278379 7984
rect 143276 7926 278379 7928
rect 143276 7924 143282 7926
rect 278313 7923 278379 7926
rect 91553 7850 91619 7853
rect 128670 7850 128676 7852
rect 91553 7848 128676 7850
rect 91553 7792 91558 7848
rect 91614 7792 128676 7848
rect 91553 7790 128676 7792
rect 91553 7787 91619 7790
rect 128670 7788 128676 7790
rect 128740 7788 128746 7852
rect 143390 7788 143396 7852
rect 143460 7850 143466 7852
rect 281901 7850 281967 7853
rect 143460 7848 281967 7850
rect 143460 7792 281906 7848
rect 281962 7792 281967 7848
rect 143460 7790 281967 7792
rect 143460 7788 143466 7790
rect 281901 7787 281967 7790
rect 87965 7714 88031 7717
rect 128854 7714 128860 7716
rect 87965 7712 128860 7714
rect 87965 7656 87970 7712
rect 88026 7656 128860 7712
rect 87965 7654 128860 7656
rect 87965 7651 88031 7654
rect 128854 7652 128860 7654
rect 128924 7652 128930 7716
rect 164918 7652 164924 7716
rect 164988 7714 164994 7716
rect 562041 7714 562107 7717
rect 164988 7712 562107 7714
rect 164988 7656 562046 7712
rect 562102 7656 562107 7712
rect 164988 7654 562107 7656
rect 164988 7652 164994 7654
rect 562041 7651 562107 7654
rect 70301 7578 70367 7581
rect 127014 7578 127020 7580
rect 70301 7576 127020 7578
rect 70301 7520 70306 7576
rect 70362 7520 127020 7576
rect 70301 7518 127020 7520
rect 70301 7515 70367 7518
rect 127014 7516 127020 7518
rect 127084 7516 127090 7580
rect 165102 7516 165108 7580
rect 165172 7578 165178 7580
rect 564433 7578 564499 7581
rect 165172 7576 564499 7578
rect 165172 7520 564438 7576
rect 564494 7520 564499 7576
rect 165172 7518 564499 7520
rect 165172 7516 165178 7518
rect 564433 7515 564499 7518
rect 138974 6836 138980 6900
rect 139044 6898 139050 6900
rect 228725 6898 228791 6901
rect 139044 6896 228791 6898
rect 139044 6840 228730 6896
rect 228786 6840 228791 6896
rect 139044 6838 228791 6840
rect 139044 6836 139050 6838
rect 228725 6835 228791 6838
rect 140630 6700 140636 6764
rect 140700 6762 140706 6764
rect 246389 6762 246455 6765
rect 140700 6760 246455 6762
rect 140700 6704 246394 6760
rect 246450 6704 246455 6760
rect 140700 6702 246455 6704
rect 140700 6700 140706 6702
rect 246389 6699 246455 6702
rect 108113 6626 108179 6629
rect 129774 6626 129780 6628
rect 108113 6624 129780 6626
rect -960 6490 480 6580
rect 108113 6568 108118 6624
rect 108174 6568 129780 6624
rect 108113 6566 129780 6568
rect 108113 6563 108179 6566
rect 129774 6564 129780 6566
rect 129844 6564 129850 6628
rect 151670 6564 151676 6628
rect 151740 6626 151746 6628
rect 385953 6626 386019 6629
rect 151740 6624 386019 6626
rect 151740 6568 385958 6624
rect 386014 6568 386019 6624
rect 151740 6566 386019 6568
rect 151740 6564 151746 6566
rect 385953 6563 386019 6566
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3509 6490 3575 6493
rect -960 6488 3575 6490
rect -960 6432 3514 6488
rect 3570 6432 3575 6488
rect -960 6430 3575 6432
rect -960 6340 480 6430
rect 3509 6427 3575 6430
rect 56041 6490 56107 6493
rect 125726 6490 125732 6492
rect 56041 6488 125732 6490
rect 56041 6432 56046 6488
rect 56102 6432 125732 6488
rect 56041 6430 125732 6432
rect 56041 6427 56107 6430
rect 125726 6428 125732 6430
rect 125796 6428 125802 6492
rect 162526 6428 162532 6492
rect 162596 6490 162602 6492
rect 526621 6490 526687 6493
rect 162596 6488 526687 6490
rect 162596 6432 526626 6488
rect 526682 6432 526687 6488
rect 583520 6476 584960 6566
rect 162596 6430 526687 6432
rect 162596 6428 162602 6430
rect 526621 6427 526687 6430
rect 52545 6354 52611 6357
rect 125910 6354 125916 6356
rect 52545 6352 125916 6354
rect 52545 6296 52550 6352
rect 52606 6296 125916 6352
rect 52545 6294 125916 6296
rect 52545 6291 52611 6294
rect 125910 6292 125916 6294
rect 125980 6292 125986 6356
rect 162710 6292 162716 6356
rect 162780 6354 162786 6356
rect 530117 6354 530183 6357
rect 162780 6352 530183 6354
rect 162780 6296 530122 6352
rect 530178 6296 530183 6352
rect 162780 6294 530183 6296
rect 162780 6292 162786 6294
rect 530117 6291 530183 6294
rect 18229 6218 18295 6221
rect 122966 6218 122972 6220
rect 18229 6216 122972 6218
rect 18229 6160 18234 6216
rect 18290 6160 122972 6216
rect 18229 6158 122972 6160
rect 18229 6155 18295 6158
rect 122966 6156 122972 6158
rect 123036 6156 123042 6220
rect 166574 6156 166580 6220
rect 166644 6218 166650 6220
rect 576301 6218 576367 6221
rect 166644 6216 576367 6218
rect 166644 6160 576306 6216
rect 576362 6160 576367 6216
rect 166644 6158 576367 6160
rect 166644 6156 166650 6158
rect 576301 6155 576367 6158
rect 139158 6020 139164 6084
rect 139228 6082 139234 6084
rect 226425 6082 226491 6085
rect 139228 6080 226491 6082
rect 139228 6024 226430 6080
rect 226486 6024 226491 6080
rect 139228 6022 226491 6024
rect 139228 6020 139234 6022
rect 226425 6019 226491 6022
rect 152958 5476 152964 5540
rect 153028 5538 153034 5540
rect 404813 5538 404879 5541
rect 153028 5536 404879 5538
rect 153028 5480 404818 5536
rect 404874 5480 404879 5536
rect 153028 5478 404879 5480
rect 153028 5476 153034 5478
rect 404813 5475 404879 5478
rect 161054 5340 161060 5404
rect 161124 5402 161130 5404
rect 508865 5402 508931 5405
rect 161124 5400 508931 5402
rect 161124 5344 508870 5400
rect 508926 5344 508931 5400
rect 161124 5342 508931 5344
rect 161124 5340 161130 5342
rect 508865 5339 508931 5342
rect 161238 5204 161244 5268
rect 161308 5266 161314 5268
rect 512453 5266 512519 5269
rect 161308 5264 512519 5266
rect 161308 5208 512458 5264
rect 512514 5208 512519 5264
rect 161308 5206 512519 5208
rect 161308 5204 161314 5206
rect 512453 5203 512519 5206
rect 163630 5068 163636 5132
rect 163700 5130 163706 5132
rect 547873 5130 547939 5133
rect 163700 5128 547939 5130
rect 163700 5072 547878 5128
rect 547934 5072 547939 5128
rect 163700 5070 547939 5072
rect 163700 5068 163706 5070
rect 547873 5067 547939 5070
rect 90357 4994 90423 4997
rect 128670 4994 128676 4996
rect 90357 4992 128676 4994
rect 90357 4936 90362 4992
rect 90418 4936 128676 4992
rect 90357 4934 128676 4936
rect 90357 4931 90423 4934
rect 128670 4932 128676 4934
rect 128740 4932 128746 4996
rect 133454 4932 133460 4996
rect 133524 4994 133530 4996
rect 155401 4994 155467 4997
rect 133524 4992 155467 4994
rect 133524 4936 155406 4992
rect 155462 4936 155467 4992
rect 133524 4934 155467 4936
rect 133524 4932 133530 4934
rect 155401 4931 155467 4934
rect 165286 4932 165292 4996
rect 165356 4994 165362 4996
rect 563237 4994 563303 4997
rect 165356 4992 563303 4994
rect 165356 4936 563242 4992
rect 563298 4936 563303 4992
rect 165356 4934 563303 4936
rect 165356 4932 165362 4934
rect 563237 4931 563303 4934
rect 37181 4858 37247 4861
rect 124254 4858 124260 4860
rect 37181 4856 124260 4858
rect 37181 4800 37186 4856
rect 37242 4800 124260 4856
rect 37181 4798 124260 4800
rect 37181 4795 37247 4798
rect 124254 4796 124260 4798
rect 124324 4796 124330 4860
rect 133270 4796 133276 4860
rect 133340 4858 133346 4860
rect 156597 4858 156663 4861
rect 133340 4856 156663 4858
rect 133340 4800 156602 4856
rect 156658 4800 156663 4856
rect 133340 4798 156663 4800
rect 133340 4796 133346 4798
rect 156597 4795 156663 4798
rect 165470 4796 165476 4860
rect 165540 4858 165546 4860
rect 565629 4858 565695 4861
rect 165540 4856 565695 4858
rect 165540 4800 565634 4856
rect 565690 4800 565695 4856
rect 165540 4798 565695 4800
rect 165540 4796 165546 4798
rect 565629 4795 565695 4798
rect 136398 4660 136404 4724
rect 136468 4722 136474 4724
rect 193305 4722 193371 4725
rect 136468 4720 193371 4722
rect 136468 4664 193310 4720
rect 193366 4664 193371 4720
rect 136468 4662 193371 4664
rect 136468 4660 136474 4662
rect 193305 4659 193371 4662
rect 167494 3980 167500 4044
rect 167564 4042 167570 4044
rect 445017 4042 445083 4045
rect 167564 4040 445083 4042
rect 167564 3984 445022 4040
rect 445078 3984 445083 4040
rect 167564 3982 445083 3984
rect 167564 3980 167570 3982
rect 445017 3979 445083 3982
rect 159030 3844 159036 3908
rect 159100 3906 159106 3908
rect 494697 3906 494763 3909
rect 159100 3904 494763 3906
rect 159100 3848 494702 3904
rect 494758 3848 494763 3904
rect 159100 3846 494763 3848
rect 159100 3844 159106 3846
rect 494697 3843 494763 3846
rect 54937 3770 55003 3773
rect 125542 3770 125548 3772
rect 54937 3768 125548 3770
rect 54937 3712 54942 3768
rect 54998 3712 125548 3768
rect 54937 3710 125548 3712
rect 54937 3707 55003 3710
rect 125542 3708 125548 3710
rect 125612 3708 125618 3772
rect 160829 3770 160895 3773
rect 505369 3770 505435 3773
rect 160829 3768 505435 3770
rect 160829 3712 160834 3768
rect 160890 3712 505374 3768
rect 505430 3712 505435 3768
rect 160829 3710 505435 3712
rect 160829 3707 160895 3710
rect 505369 3707 505435 3710
rect 17033 3634 17099 3637
rect 122598 3634 122604 3636
rect 17033 3632 122604 3634
rect 17033 3576 17038 3632
rect 17094 3576 122604 3632
rect 17033 3574 122604 3576
rect 17033 3571 17099 3574
rect 122598 3572 122604 3574
rect 122668 3572 122674 3636
rect 123477 3634 123543 3637
rect 131246 3634 131252 3636
rect 123477 3632 131252 3634
rect 123477 3576 123482 3632
rect 123538 3576 131252 3632
rect 123477 3574 131252 3576
rect 123477 3571 123543 3574
rect 131246 3572 131252 3574
rect 131316 3572 131322 3636
rect 131798 3572 131804 3636
rect 131868 3634 131874 3636
rect 137645 3634 137711 3637
rect 131868 3632 137711 3634
rect 131868 3576 137650 3632
rect 137706 3576 137711 3632
rect 131868 3574 137711 3576
rect 131868 3572 131874 3574
rect 137645 3571 137711 3574
rect 167862 3572 167868 3636
rect 167932 3634 167938 3636
rect 533705 3634 533771 3637
rect 167932 3632 533771 3634
rect 167932 3576 533710 3632
rect 533766 3576 533771 3632
rect 167932 3574 533771 3576
rect 167932 3572 167938 3574
rect 533705 3571 533771 3574
rect 1669 3498 1735 3501
rect 121678 3498 121684 3500
rect 1669 3496 121684 3498
rect 1669 3440 1674 3496
rect 1730 3440 121684 3496
rect 1669 3438 121684 3440
rect 1669 3435 1735 3438
rect 121678 3436 121684 3438
rect 121748 3436 121754 3500
rect 124673 3498 124739 3501
rect 131062 3498 131068 3500
rect 124673 3496 131068 3498
rect 124673 3440 124678 3496
rect 124734 3440 131068 3496
rect 124673 3438 131068 3440
rect 124673 3435 124739 3438
rect 131062 3436 131068 3438
rect 131132 3436 131138 3500
rect 131982 3436 131988 3500
rect 132052 3498 132058 3500
rect 140037 3498 140103 3501
rect 132052 3496 140103 3498
rect 132052 3440 140042 3496
rect 140098 3440 140103 3496
rect 132052 3438 140103 3440
rect 132052 3436 132058 3438
rect 140037 3435 140103 3438
rect 167678 3436 167684 3500
rect 167748 3498 167754 3500
rect 537201 3498 537267 3501
rect 167748 3496 537267 3498
rect 167748 3440 537206 3496
rect 537262 3440 537267 3496
rect 167748 3438 537267 3440
rect 167748 3436 167754 3438
rect 537201 3435 537267 3438
rect 565 3362 631 3365
rect 121494 3362 121500 3364
rect 565 3360 121500 3362
rect 565 3304 570 3360
rect 626 3304 121500 3360
rect 565 3302 121500 3304
rect 565 3299 631 3302
rect 121494 3300 121500 3302
rect 121564 3300 121570 3364
rect 133638 3300 133644 3364
rect 133708 3362 133714 3364
rect 157793 3362 157859 3365
rect 133708 3360 157859 3362
rect 133708 3304 157798 3360
rect 157854 3304 157859 3360
rect 133708 3302 157859 3304
rect 133708 3300 133714 3302
rect 157793 3299 157859 3302
rect 166758 3300 166764 3364
rect 166828 3362 166834 3364
rect 583385 3362 583451 3365
rect 166828 3360 583451 3362
rect 166828 3304 583390 3360
rect 583446 3304 583451 3360
rect 166828 3302 583451 3304
rect 166828 3300 166834 3302
rect 583385 3299 583451 3302
<< via3 >>
rect 542676 699756 542740 699820
rect 580212 697172 580276 697236
rect 3372 658140 3436 658204
rect 396580 418236 396644 418300
rect 396764 240076 396828 240140
rect 396948 239940 397012 240004
rect 396764 232324 396828 232388
rect 396948 231100 397012 231164
rect 143580 191568 143644 191632
rect 144684 190980 144748 191044
rect 144500 190632 144564 190636
rect 144500 190576 144514 190632
rect 144514 190576 144564 190632
rect 144500 190572 144564 190576
rect 145788 189816 145852 189820
rect 145788 189760 145838 189816
rect 145838 189760 145852 189816
rect 145788 189756 145852 189760
rect 143028 184316 143092 184380
rect 141372 184180 141436 184244
rect 144500 183772 144564 183836
rect 144684 183696 144748 183700
rect 144684 183640 144698 183696
rect 144698 183640 144748 183696
rect 144684 183636 144748 183640
rect 140636 182548 140700 182612
rect 145972 181188 146036 181252
rect 143396 180916 143460 180980
rect 142292 179012 142356 179076
rect 143028 178876 143092 178940
rect 141372 178740 141436 178804
rect 140636 175612 140700 175676
rect 145972 174116 146036 174180
rect 143580 138756 143644 138820
rect 396580 138620 396644 138684
rect 141924 137940 141988 138004
rect 146156 137532 146220 137596
rect 143396 137396 143460 137460
rect 542676 137260 542740 137324
rect 169524 75244 169588 75308
rect 167868 75108 167932 75172
rect 167500 74836 167564 74900
rect 167868 74836 167932 74900
rect 161612 74760 161676 74764
rect 161612 74704 161662 74760
rect 161662 74704 161676 74760
rect 161612 74700 161676 74704
rect 164740 74760 164804 74764
rect 580212 74836 580276 74900
rect 164740 74704 164754 74760
rect 164754 74704 164804 74760
rect 164740 74700 164804 74704
rect 169524 74760 169588 74764
rect 169524 74704 169574 74760
rect 169574 74704 169588 74760
rect 169524 74700 169588 74704
rect 164924 74216 164988 74220
rect 164924 74160 164938 74216
rect 164938 74160 164988 74216
rect 164924 74156 164988 74160
rect 3372 73884 3436 73948
rect 166764 73400 166828 73404
rect 166764 73344 166814 73400
rect 166814 73344 166828 73400
rect 166764 73340 166828 73344
rect 128492 73128 128556 73132
rect 128492 73072 128542 73128
rect 128542 73072 128556 73128
rect 128492 73068 128556 73072
rect 165844 73068 165908 73132
rect 152412 72932 152476 72996
rect 148364 72796 148428 72860
rect 149652 72796 149716 72860
rect 151308 72796 151372 72860
rect 152780 72796 152844 72860
rect 154436 72796 154500 72860
rect 157012 72856 157076 72860
rect 157012 72800 157026 72856
rect 157026 72800 157076 72856
rect 157012 72796 157076 72800
rect 158484 72796 158548 72860
rect 158852 72796 158916 72860
rect 160876 72796 160940 72860
rect 162348 72796 162412 72860
rect 163452 72796 163516 72860
rect 164924 72856 164988 72860
rect 164924 72800 164938 72856
rect 164938 72800 164988 72856
rect 164924 72796 164988 72800
rect 165292 72856 165356 72860
rect 165292 72800 165342 72856
rect 165342 72800 165356 72856
rect 165292 72796 165356 72800
rect 166580 72796 166644 72860
rect 148732 72720 148796 72724
rect 148732 72664 148746 72720
rect 148746 72664 148796 72720
rect 148732 72660 148796 72664
rect 148916 72720 148980 72724
rect 148916 72664 148966 72720
rect 148966 72664 148980 72720
rect 148916 72660 148980 72664
rect 150020 72720 150084 72724
rect 150020 72664 150034 72720
rect 150034 72664 150084 72720
rect 150020 72660 150084 72664
rect 151676 72660 151740 72724
rect 152964 72720 153028 72724
rect 152964 72664 153014 72720
rect 153014 72664 153028 72720
rect 152964 72660 153028 72664
rect 154252 72720 154316 72724
rect 154252 72664 154266 72720
rect 154266 72664 154316 72720
rect 154252 72660 154316 72664
rect 155724 72660 155788 72724
rect 156828 72720 156892 72724
rect 156828 72664 156878 72720
rect 156878 72664 156892 72720
rect 156828 72660 156892 72664
rect 157196 72720 157260 72724
rect 157196 72664 157246 72720
rect 157246 72664 157260 72720
rect 157196 72660 157260 72664
rect 158668 72660 158732 72724
rect 159036 72660 159100 72724
rect 161060 72720 161124 72724
rect 161060 72664 161110 72720
rect 161110 72664 161124 72720
rect 161060 72660 161124 72664
rect 161244 72660 161308 72724
rect 162532 72720 162596 72724
rect 162532 72664 162546 72720
rect 162546 72664 162596 72720
rect 162532 72660 162596 72664
rect 162716 72720 162780 72724
rect 162716 72664 162766 72720
rect 162766 72664 162780 72720
rect 162716 72660 162780 72664
rect 163636 72660 163700 72724
rect 164924 72660 164988 72724
rect 165476 72720 165540 72724
rect 165476 72664 165526 72720
rect 165526 72664 165540 72720
rect 165476 72660 165540 72664
rect 166396 72660 166460 72724
rect 149468 72524 149532 72588
rect 152596 72524 152660 72588
rect 153884 72524 153948 72588
rect 156644 72524 156708 72588
rect 158300 72524 158364 72588
rect 160692 72524 160756 72588
rect 161612 72524 161676 72588
rect 163268 72524 163332 72588
rect 165108 72524 165172 72588
rect 148548 72388 148612 72452
rect 149836 72388 149900 72452
rect 151492 72388 151556 72452
rect 154068 72388 154132 72452
rect 155540 72388 155604 72452
rect 158116 72388 158180 72452
rect 162164 72388 162228 72452
rect 126100 72252 126164 72316
rect 146892 72252 146956 72316
rect 124628 72116 124692 72180
rect 125916 72116 125980 72180
rect 129044 72116 129108 72180
rect 129964 72116 130028 72180
rect 133276 72116 133340 72180
rect 134748 72116 134812 72180
rect 135852 72116 135916 72180
rect 138980 72116 139044 72180
rect 140084 72116 140148 72180
rect 142844 72116 142908 72180
rect 144132 72116 144196 72180
rect 145236 72116 145300 72180
rect 147076 72116 147140 72180
rect 121684 72040 121748 72044
rect 121684 71984 121698 72040
rect 121698 71984 121748 72040
rect 121684 71980 121748 71984
rect 122788 72040 122852 72044
rect 122788 71984 122838 72040
rect 122838 71984 122852 72040
rect 122788 71980 122852 71984
rect 124260 71980 124324 72044
rect 125548 71980 125612 72044
rect 127204 71980 127268 72044
rect 128860 71980 128924 72044
rect 130148 71980 130212 72044
rect 131068 71980 131132 72044
rect 131804 71980 131868 72044
rect 133460 71980 133524 72044
rect 134932 72040 134996 72044
rect 134932 71984 134982 72040
rect 134982 71984 134996 72040
rect 134932 71980 134996 71984
rect 136220 71980 136284 72044
rect 137692 71980 137756 72044
rect 138796 71980 138860 72044
rect 140268 71980 140332 72044
rect 140820 71980 140884 72044
rect 143028 71980 143092 72044
rect 144500 71980 144564 72044
rect 145420 71980 145484 72044
rect 147260 71980 147324 72044
rect 121500 71904 121564 71908
rect 121500 71848 121550 71904
rect 121550 71848 121564 71904
rect 121500 71844 121564 71848
rect 122972 71904 123036 71908
rect 122972 71848 122986 71904
rect 122986 71848 123036 71904
rect 122972 71844 123036 71848
rect 124444 71904 124508 71908
rect 124444 71848 124494 71904
rect 124494 71848 124508 71904
rect 124444 71844 124508 71848
rect 125732 71844 125796 71908
rect 127020 71904 127084 71908
rect 127020 71848 127034 71904
rect 127034 71848 127084 71904
rect 127020 71844 127084 71848
rect 128676 71904 128740 71908
rect 128676 71848 128690 71904
rect 128690 71848 128740 71904
rect 128676 71844 128740 71848
rect 129780 71844 129844 71908
rect 131252 71844 131316 71908
rect 131988 71844 132052 71908
rect 133644 71844 133708 71908
rect 135116 71904 135180 71908
rect 135116 71848 135166 71904
rect 135166 71848 135180 71904
rect 135116 71844 135180 71848
rect 136036 71844 136100 71908
rect 136404 71844 136468 71908
rect 137876 71904 137940 71908
rect 137876 71848 137926 71904
rect 137926 71848 137940 71904
rect 137876 71844 137940 71848
rect 138612 71844 138676 71908
rect 139164 71904 139228 71908
rect 139164 71848 139178 71904
rect 139178 71848 139228 71904
rect 139164 71844 139228 71848
rect 140452 71904 140516 71908
rect 140452 71848 140466 71904
rect 140466 71848 140516 71904
rect 140452 71844 140516 71848
rect 140636 71904 140700 71908
rect 140636 71848 140686 71904
rect 140686 71848 140700 71904
rect 140636 71844 140700 71848
rect 141004 71844 141068 71908
rect 143212 71904 143276 71908
rect 143212 71848 143226 71904
rect 143226 71848 143276 71904
rect 143212 71844 143276 71848
rect 143396 71904 143460 71908
rect 143396 71848 143446 71904
rect 143446 71848 143460 71904
rect 143396 71844 143460 71848
rect 144316 71844 144380 71908
rect 144684 71844 144748 71908
rect 145604 71844 145668 71908
rect 147444 71844 147508 71908
rect 164740 71360 164804 71364
rect 164740 71304 164754 71360
rect 164754 71304 164804 71360
rect 164740 71300 164804 71304
rect 165844 71164 165908 71228
rect 167868 71164 167932 71228
rect 167684 70076 167748 70140
rect 158668 65452 158732 65516
rect 144132 35260 144196 35324
rect 146892 35124 146956 35188
rect 137692 34036 137756 34100
rect 140084 33900 140148 33964
rect 140820 33764 140884 33828
rect 134748 32676 134812 32740
rect 136036 32540 136100 32604
rect 135852 32404 135916 32468
rect 163268 31180 163332 31244
rect 158116 31044 158180 31108
rect 158852 30908 158916 30972
rect 145236 29548 145300 29612
rect 136220 27100 136284 27164
rect 142844 26964 142908 27028
rect 149468 26828 149532 26892
rect 134932 25604 134996 25668
rect 156644 25468 156708 25532
rect 151308 24380 151372 24444
rect 162164 24244 162228 24308
rect 163452 24108 163516 24172
rect 155540 22884 155604 22948
rect 156828 22748 156892 22812
rect 160692 22612 160756 22676
rect 148364 21388 148428 21452
rect 158300 21252 158364 21316
rect 138612 20164 138676 20228
rect 140268 20028 140332 20092
rect 158484 19892 158548 19956
rect 157012 18804 157076 18868
rect 157196 18668 157260 18732
rect 162348 18532 162412 18596
rect 145420 17580 145484 17644
rect 154068 17444 154132 17508
rect 153884 17308 153948 17372
rect 155724 17172 155788 17236
rect 144316 16220 144380 16284
rect 148548 16084 148612 16148
rect 152412 15948 152476 16012
rect 154252 15812 154316 15876
rect 141004 15132 141068 15196
rect 144500 14996 144564 15060
rect 145604 14860 145668 14924
rect 147076 14724 147140 14788
rect 151492 14588 151556 14652
rect 152596 14452 152660 14516
rect 140452 13636 140516 13700
rect 143028 13500 143092 13564
rect 149836 13364 149900 13428
rect 149652 13228 149716 13292
rect 154436 13092 154500 13156
rect 160876 12956 160940 13020
rect 138796 12820 138860 12884
rect 137876 12140 137940 12204
rect 148732 12004 148796 12068
rect 148916 11868 148980 11932
rect 150020 11732 150084 11796
rect 152780 11596 152844 11660
rect 129044 10372 129108 10436
rect 147444 10372 147508 10436
rect 127204 10236 127268 10300
rect 147260 10236 147324 10300
rect 130148 9420 130212 9484
rect 129964 9284 130028 9348
rect 126100 9148 126164 9212
rect 124444 9012 124508 9076
rect 144684 9012 144748 9076
rect 124628 8876 124692 8940
rect 166396 8876 166460 8940
rect 135116 8060 135180 8124
rect 143212 7924 143276 7988
rect 128676 7788 128740 7852
rect 143396 7788 143460 7852
rect 128860 7652 128924 7716
rect 164924 7652 164988 7716
rect 127020 7516 127084 7580
rect 165108 7516 165172 7580
rect 138980 6836 139044 6900
rect 140636 6700 140700 6764
rect 129780 6564 129844 6628
rect 151676 6564 151740 6628
rect 125732 6428 125796 6492
rect 162532 6428 162596 6492
rect 125916 6292 125980 6356
rect 162716 6292 162780 6356
rect 122972 6156 123036 6220
rect 166580 6156 166644 6220
rect 139164 6020 139228 6084
rect 152964 5476 153028 5540
rect 161060 5340 161124 5404
rect 161244 5204 161308 5268
rect 163636 5068 163700 5132
rect 128676 4932 128740 4996
rect 133460 4932 133524 4996
rect 165292 4932 165356 4996
rect 124260 4796 124324 4860
rect 133276 4796 133340 4860
rect 165476 4796 165540 4860
rect 136404 4660 136468 4724
rect 167500 3980 167564 4044
rect 159036 3844 159100 3908
rect 125548 3708 125612 3772
rect 122604 3572 122668 3636
rect 131252 3572 131316 3636
rect 131804 3572 131868 3636
rect 167868 3572 167932 3636
rect 121684 3436 121748 3500
rect 131068 3436 131132 3500
rect 131988 3436 132052 3500
rect 167684 3436 167748 3500
rect 121500 3300 121564 3364
rect 133644 3300 133708 3364
rect 166764 3300 166828 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 3371 658204 3437 658205
rect 3371 658140 3372 658204
rect 3436 658140 3437 658204
rect 3371 658139 3437 658140
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 3374 73949 3434 658139
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 3371 73948 3437 73949
rect 3371 73884 3372 73948
rect 3436 73884 3437 73948
rect 3371 73883 3437 73884
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 248684 47414 263898
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 248684 51914 268398
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 248684 56414 272898
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 248684 60914 277398
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 248684 65414 281898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 248684 69914 250398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 248684 74414 254898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 248684 78914 259398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 248684 83414 263898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 248684 87914 268398
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 248684 92414 272898
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 248684 96914 277398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 248684 101414 281898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 248684 105914 250398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 248684 110414 254898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 248684 114914 259398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 248684 119414 263898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 248684 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 248684 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 248684 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 248684 137414 281898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 248684 141914 250398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 248684 146414 254898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 248684 150914 259398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 248684 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 248684 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 248684 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 248684 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 248684 173414 281898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 248684 177914 250398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 248684 182414 254898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 248684 186914 259398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 248684 191414 263898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 248684 195914 268398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 248684 200414 272898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 248684 204914 277398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 248684 209414 281898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 248684 213914 250398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 248684 218414 254898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 248684 222914 259398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 248684 227414 263898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 248684 231914 268398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 248684 236414 272898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 248684 240914 277398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 248684 245414 281898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 248684 249914 250398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 248684 254414 254898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 248684 258914 259398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 248684 263414 263898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 248684 267914 268398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 248684 272414 272898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 248684 276914 277398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 248684 281414 281898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 248684 285914 250398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 248684 290414 254898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 248684 294914 259398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 248684 299414 263898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 248684 303914 268398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 248684 308414 272898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 248684 312914 277398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 248684 317414 281898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 248684 321914 250398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 248684 326414 254898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 248684 330914 259398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 248684 335414 263898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 248684 339914 268398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 248684 344414 272898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 248684 348914 277398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 248684 353414 281898
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 248684 357914 250398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 248684 362414 254898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 248684 366914 259398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 248684 371414 263898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 248684 375914 268398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 248684 380414 272898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 248684 384914 277398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 248684 389414 281898
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 396579 418300 396645 418301
rect 396579 418236 396580 418300
rect 396644 418236 396645 418300
rect 396579 418235 396645 418236
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 248684 393914 250398
rect 65300 246303 70100 246486
rect 65300 246067 65342 246303
rect 65578 246067 65662 246303
rect 65898 246067 65982 246303
rect 66218 246067 66302 246303
rect 66538 246067 66622 246303
rect 66858 246067 66942 246303
rect 67178 246067 67262 246303
rect 67498 246067 67582 246303
rect 67818 246067 67902 246303
rect 68138 246067 68222 246303
rect 68458 246067 68542 246303
rect 68778 246067 68862 246303
rect 69098 246067 69182 246303
rect 69418 246067 69502 246303
rect 69738 246067 69822 246303
rect 70058 246067 70100 246303
rect 65300 245884 70100 246067
rect 65300 241953 71300 241984
rect 65300 241717 65462 241953
rect 65698 241717 65782 241953
rect 66018 241717 66102 241953
rect 66338 241717 66422 241953
rect 66658 241717 66742 241953
rect 66978 241717 67062 241953
rect 67298 241717 67382 241953
rect 67618 241717 67702 241953
rect 67938 241717 68022 241953
rect 68258 241717 68342 241953
rect 68578 241717 68662 241953
rect 68898 241717 68982 241953
rect 69218 241717 69302 241953
rect 69538 241717 69622 241953
rect 69858 241717 69942 241953
rect 70178 241717 70262 241953
rect 70498 241717 70582 241953
rect 70818 241717 70902 241953
rect 71138 241717 71300 241953
rect 65300 241633 71300 241717
rect 65300 241397 65462 241633
rect 65698 241397 65782 241633
rect 66018 241397 66102 241633
rect 66338 241397 66422 241633
rect 66658 241397 66742 241633
rect 66978 241397 67062 241633
rect 67298 241397 67382 241633
rect 67618 241397 67702 241633
rect 67938 241397 68022 241633
rect 68258 241397 68342 241633
rect 68578 241397 68662 241633
rect 68898 241397 68982 241633
rect 69218 241397 69302 241633
rect 69538 241397 69622 241633
rect 69858 241397 69942 241633
rect 70178 241397 70262 241633
rect 70498 241397 70582 241633
rect 70818 241397 70902 241633
rect 71138 241397 71300 241633
rect 65300 241366 71300 241397
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 228453 47414 228484
rect 46794 228217 46826 228453
rect 47062 228217 47146 228453
rect 47382 228217 47414 228453
rect 46794 228133 47414 228217
rect 46794 227897 46826 228133
rect 47062 227897 47146 228133
rect 47382 227897 47414 228133
rect 46794 192454 47414 227897
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 196954 51914 228484
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 201454 56414 228484
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 205954 60914 228484
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 210454 65414 228484
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 214954 69914 228484
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 219454 74414 228484
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 223954 78914 228484
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 228453 83414 228484
rect 82794 228217 82826 228453
rect 83062 228217 83146 228453
rect 83382 228217 83414 228453
rect 82794 228133 83414 228217
rect 82794 227897 82826 228133
rect 83062 227897 83146 228133
rect 83382 227897 83414 228133
rect 82794 192454 83414 227897
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 196954 87914 228484
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 201454 92414 228484
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 205954 96914 228484
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 210454 101414 228484
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 214954 105914 228484
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 219454 110414 228484
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 114294 223954 114914 228484
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 137000 114914 151398
rect 118794 228453 119414 228484
rect 118794 228217 118826 228453
rect 119062 228217 119146 228453
rect 119382 228217 119414 228453
rect 118794 228133 119414 228217
rect 118794 227897 118826 228133
rect 119062 227897 119146 228133
rect 119382 227897 119414 228133
rect 118794 192454 119414 227897
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 137000 119414 155898
rect 123294 196954 123914 228484
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 137000 123914 160398
rect 127794 201454 128414 228484
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 137000 128414 164898
rect 132294 205954 132914 228484
rect 172794 210454 173414 228484
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 135914 205861 165514 205986
rect 135914 205625 136036 205861
rect 136272 205625 136356 205861
rect 136592 205625 136676 205861
rect 136912 205625 136996 205861
rect 137232 205625 137316 205861
rect 137552 205625 137636 205861
rect 137872 205625 137956 205861
rect 138192 205625 138276 205861
rect 138512 205625 138596 205861
rect 138832 205625 138916 205861
rect 139152 205625 139236 205861
rect 139472 205625 139556 205861
rect 139792 205625 139876 205861
rect 140112 205625 140196 205861
rect 140432 205625 140516 205861
rect 140752 205625 140836 205861
rect 141072 205625 141156 205861
rect 141392 205625 141476 205861
rect 141712 205625 141796 205861
rect 142032 205625 142116 205861
rect 142352 205625 142436 205861
rect 142672 205625 142756 205861
rect 142992 205625 143076 205861
rect 143312 205625 143396 205861
rect 143632 205625 143716 205861
rect 143952 205625 144036 205861
rect 144272 205625 144356 205861
rect 144592 205625 144676 205861
rect 144912 205625 144996 205861
rect 145232 205625 145316 205861
rect 145552 205625 145636 205861
rect 145872 205625 145956 205861
rect 146192 205625 146276 205861
rect 146512 205625 146596 205861
rect 146832 205625 146916 205861
rect 147152 205625 147236 205861
rect 147472 205625 147556 205861
rect 147792 205625 147876 205861
rect 148112 205625 148196 205861
rect 148432 205625 148516 205861
rect 148752 205625 148836 205861
rect 149072 205625 149156 205861
rect 149392 205625 149476 205861
rect 149712 205625 149796 205861
rect 150032 205625 150116 205861
rect 150352 205625 150436 205861
rect 150672 205625 150756 205861
rect 150992 205625 151076 205861
rect 151312 205625 151396 205861
rect 151632 205625 151716 205861
rect 151952 205625 152036 205861
rect 152272 205625 152356 205861
rect 152592 205625 152676 205861
rect 152912 205625 152996 205861
rect 153232 205625 153316 205861
rect 153552 205625 153636 205861
rect 153872 205625 153956 205861
rect 154192 205625 154276 205861
rect 154512 205625 154596 205861
rect 154832 205625 154916 205861
rect 155152 205625 155236 205861
rect 155472 205625 155556 205861
rect 155792 205625 155876 205861
rect 156112 205625 156196 205861
rect 156432 205625 156516 205861
rect 156752 205625 156836 205861
rect 157072 205625 157156 205861
rect 157392 205625 157476 205861
rect 157712 205625 157796 205861
rect 158032 205625 158116 205861
rect 158352 205625 158436 205861
rect 158672 205625 158756 205861
rect 158992 205625 159076 205861
rect 159312 205625 159396 205861
rect 159632 205625 159716 205861
rect 159952 205625 160036 205861
rect 160272 205625 160356 205861
rect 160592 205625 160676 205861
rect 160912 205625 160996 205861
rect 161232 205625 161316 205861
rect 161552 205625 161636 205861
rect 161872 205625 161956 205861
rect 162192 205625 162276 205861
rect 162512 205625 162596 205861
rect 162832 205625 162916 205861
rect 163152 205625 163236 205861
rect 163472 205625 163556 205861
rect 163792 205625 163876 205861
rect 164112 205625 164196 205861
rect 164432 205625 164516 205861
rect 164752 205625 164836 205861
rect 165072 205625 165156 205861
rect 165392 205625 165514 205861
rect 135914 205500 165514 205625
rect 132294 169954 132914 205398
rect 137314 201411 165514 201486
rect 137314 201175 137376 201411
rect 137612 201175 137696 201411
rect 137932 201175 138016 201411
rect 138252 201175 138336 201411
rect 138572 201175 138656 201411
rect 138892 201175 138976 201411
rect 139212 201175 139296 201411
rect 139532 201175 139616 201411
rect 139852 201175 139936 201411
rect 140172 201175 140256 201411
rect 140492 201175 140576 201411
rect 140812 201175 140896 201411
rect 141132 201175 141216 201411
rect 141452 201175 141536 201411
rect 141772 201175 141856 201411
rect 142092 201175 142176 201411
rect 142412 201175 142496 201411
rect 142732 201175 142816 201411
rect 143052 201175 143136 201411
rect 143372 201175 143456 201411
rect 143692 201175 143776 201411
rect 144012 201175 144096 201411
rect 144332 201175 144416 201411
rect 144652 201175 144736 201411
rect 144972 201175 145056 201411
rect 145292 201175 145376 201411
rect 145612 201175 145696 201411
rect 145932 201175 146016 201411
rect 146252 201175 146336 201411
rect 146572 201175 146656 201411
rect 146892 201175 146976 201411
rect 147212 201175 147296 201411
rect 147532 201175 147616 201411
rect 147852 201175 147936 201411
rect 148172 201175 148256 201411
rect 148492 201175 148576 201411
rect 148812 201175 148896 201411
rect 149132 201175 149216 201411
rect 149452 201175 149536 201411
rect 149772 201175 149856 201411
rect 150092 201175 150176 201411
rect 150412 201175 150496 201411
rect 150732 201175 150816 201411
rect 151052 201175 151136 201411
rect 151372 201175 151456 201411
rect 151692 201175 151776 201411
rect 152012 201175 152096 201411
rect 152332 201175 152416 201411
rect 152652 201175 152736 201411
rect 152972 201175 153056 201411
rect 153292 201175 153376 201411
rect 153612 201175 153696 201411
rect 153932 201175 154016 201411
rect 154252 201175 154336 201411
rect 154572 201175 154656 201411
rect 154892 201175 154976 201411
rect 155212 201175 155296 201411
rect 155532 201175 155616 201411
rect 155852 201175 155936 201411
rect 156172 201175 156256 201411
rect 156492 201175 156576 201411
rect 156812 201175 156896 201411
rect 157132 201175 157216 201411
rect 157452 201175 157536 201411
rect 157772 201175 157856 201411
rect 158092 201175 158176 201411
rect 158412 201175 158496 201411
rect 158732 201175 158816 201411
rect 159052 201175 159136 201411
rect 159372 201175 159456 201411
rect 159692 201175 159776 201411
rect 160012 201175 160096 201411
rect 160332 201175 160416 201411
rect 160652 201175 160736 201411
rect 160972 201175 161056 201411
rect 161292 201175 161376 201411
rect 161612 201175 161696 201411
rect 161932 201175 162016 201411
rect 162252 201175 162336 201411
rect 162572 201175 162656 201411
rect 162892 201175 162976 201411
rect 163212 201175 163296 201411
rect 163532 201175 163616 201411
rect 163852 201175 163936 201411
rect 164172 201175 164256 201411
rect 164492 201175 164576 201411
rect 164812 201175 164896 201411
rect 165132 201175 165216 201411
rect 165452 201175 165514 201411
rect 137314 201100 165514 201175
rect 143579 191632 143645 191633
rect 143579 191568 143580 191632
rect 143644 191568 143645 191632
rect 143579 191567 143645 191568
rect 143027 184380 143093 184381
rect 143027 184316 143028 184380
rect 143092 184316 143093 184380
rect 143027 184315 143093 184316
rect 141371 184244 141437 184245
rect 141371 184180 141372 184244
rect 141436 184180 141437 184244
rect 141371 184179 141437 184180
rect 140635 182612 140701 182613
rect 140635 182548 140636 182612
rect 140700 182548 140701 182612
rect 140635 182547 140701 182548
rect 140638 175677 140698 182547
rect 141374 178805 141434 184179
rect 142291 179076 142357 179077
rect 142291 179012 142292 179076
rect 142356 179012 142357 179076
rect 142291 179011 142357 179012
rect 141371 178804 141437 178805
rect 141371 178740 141372 178804
rect 141436 178740 141437 178804
rect 141371 178739 141437 178740
rect 142294 176670 142354 179011
rect 143030 178941 143090 184315
rect 143395 180980 143461 180981
rect 143395 180916 143396 180980
rect 143460 180916 143461 180980
rect 143395 180915 143461 180916
rect 143027 178940 143093 178941
rect 143027 178876 143028 178940
rect 143092 178876 143093 178940
rect 143027 178875 143093 178876
rect 142110 176610 142354 176670
rect 140635 175676 140701 175677
rect 140635 175612 140636 175676
rect 140700 175612 140701 175676
rect 140635 175611 140701 175612
rect 137014 174454 141514 174486
rect 137014 174218 137066 174454
rect 137302 174218 137386 174454
rect 137622 174218 137706 174454
rect 137942 174218 138026 174454
rect 138262 174218 138346 174454
rect 138582 174218 138666 174454
rect 138902 174218 138986 174454
rect 139222 174218 139306 174454
rect 139542 174218 139626 174454
rect 139862 174218 139946 174454
rect 140182 174218 140266 174454
rect 140502 174218 140586 174454
rect 140822 174218 140906 174454
rect 141142 174218 141226 174454
rect 141462 174218 141514 174454
rect 137014 174134 141514 174218
rect 137014 173898 137066 174134
rect 137302 173898 137386 174134
rect 137622 173898 137706 174134
rect 137942 173898 138026 174134
rect 138262 173898 138346 174134
rect 138582 173898 138666 174134
rect 138902 173898 138986 174134
rect 139222 173898 139306 174134
rect 139542 173898 139626 174134
rect 139862 173898 139946 174134
rect 140182 173898 140266 174134
rect 140502 173898 140586 174134
rect 140822 173898 140906 174134
rect 141142 173898 141226 174134
rect 141462 173898 141514 174134
rect 137014 173866 141514 173898
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 137000 132914 169398
rect 142110 167010 142170 176610
rect 141926 166950 142170 167010
rect 141926 138005 141986 166950
rect 141923 138004 141989 138005
rect 141923 137940 141924 138004
rect 141988 137940 141989 138004
rect 141923 137939 141989 137940
rect 143398 137461 143458 180915
rect 143582 138821 143642 191567
rect 144683 191044 144749 191045
rect 144683 190980 144684 191044
rect 144748 190980 144749 191044
rect 144683 190979 144749 190980
rect 144499 190636 144565 190637
rect 144499 190572 144500 190636
rect 144564 190572 144565 190636
rect 144499 190571 144565 190572
rect 144502 183837 144562 190571
rect 144499 183836 144565 183837
rect 144499 183772 144500 183836
rect 144564 183772 144565 183836
rect 144499 183771 144565 183772
rect 144686 183701 144746 190979
rect 145787 189820 145853 189821
rect 145787 189756 145788 189820
rect 145852 189756 145853 189820
rect 145787 189755 145853 189756
rect 145790 184950 145850 189755
rect 145790 184890 146218 184950
rect 144683 183700 144749 183701
rect 144683 183636 144684 183700
rect 144748 183636 144749 183700
rect 144683 183635 144749 183636
rect 145971 181252 146037 181253
rect 145971 181188 145972 181252
rect 146036 181188 146037 181252
rect 145971 181187 146037 181188
rect 145974 174181 146034 181187
rect 145971 174180 146037 174181
rect 145971 174116 145972 174180
rect 146036 174116 146037 174180
rect 145971 174115 146037 174116
rect 143579 138820 143645 138821
rect 143579 138756 143580 138820
rect 143644 138756 143645 138820
rect 143579 138755 143645 138756
rect 146158 137597 146218 184890
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 146155 137596 146221 137597
rect 146155 137532 146156 137596
rect 146220 137532 146221 137596
rect 146155 137531 146221 137532
rect 143395 137460 143461 137461
rect 143395 137396 143396 137460
rect 143460 137396 143461 137460
rect 143395 137395 143461 137396
rect 172794 137000 173414 137898
rect 177294 214954 177914 228484
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 137000 177914 142398
rect 181794 219454 182414 228484
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 135568 115954 135888 115986
rect 135568 115718 135610 115954
rect 135846 115718 135888 115954
rect 135568 115634 135888 115718
rect 135568 115398 135610 115634
rect 135846 115398 135888 115634
rect 135568 115366 135888 115398
rect 166288 115954 166608 115986
rect 166288 115718 166330 115954
rect 166566 115718 166608 115954
rect 166288 115634 166608 115718
rect 166288 115398 166330 115634
rect 166566 115398 166608 115634
rect 166288 115366 166608 115398
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 120208 111454 120528 111486
rect 120208 111218 120250 111454
rect 120486 111218 120528 111454
rect 120208 111134 120528 111218
rect 120208 110898 120250 111134
rect 120486 110898 120528 111134
rect 120208 110866 120528 110898
rect 150928 111454 151248 111486
rect 150928 111218 150970 111454
rect 151206 111218 151248 111454
rect 150928 111134 151248 111218
rect 150928 110898 150970 111134
rect 151206 110898 151248 111134
rect 150928 110866 151248 110898
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 135568 79954 135888 79986
rect 135568 79718 135610 79954
rect 135846 79718 135888 79954
rect 135568 79634 135888 79718
rect 135568 79398 135610 79634
rect 135846 79398 135888 79634
rect 135568 79366 135888 79398
rect 166288 79954 166608 79986
rect 166288 79718 166330 79954
rect 166566 79718 166608 79954
rect 166288 79634 166608 79718
rect 166288 79398 166330 79634
rect 166566 79398 166608 79634
rect 166288 79366 166608 79398
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 181794 75454 182414 110898
rect 169523 75308 169589 75309
rect 169523 75244 169524 75308
rect 169588 75244 169589 75308
rect 169523 75243 169589 75244
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 167867 75172 167933 75173
rect 167867 75108 167868 75172
rect 167932 75108 167933 75172
rect 167867 75107 167933 75108
rect 167870 74901 167930 75107
rect 109794 39454 110414 74898
rect 167499 74900 167565 74901
rect 167499 74836 167500 74900
rect 167564 74836 167565 74900
rect 167499 74835 167565 74836
rect 167867 74900 167933 74901
rect 167867 74836 167868 74900
rect 167932 74836 167933 74900
rect 167867 74835 167933 74836
rect 161611 74764 161677 74765
rect 161611 74700 161612 74764
rect 161676 74700 161677 74764
rect 161611 74699 161677 74700
rect 164739 74764 164805 74765
rect 164739 74700 164740 74764
rect 164804 74700 164805 74764
rect 164739 74699 164805 74700
rect 128491 73132 128557 73133
rect 128491 73068 128492 73132
rect 128556 73068 128557 73132
rect 128491 73067 128557 73068
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 43954 114914 73000
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 73000
rect 121683 72044 121749 72045
rect 121683 71980 121684 72044
rect 121748 71980 121749 72044
rect 121683 71979 121749 71980
rect 122787 72044 122853 72045
rect 122787 71980 122788 72044
rect 122852 71980 122853 72044
rect 122787 71979 122853 71980
rect 121499 71908 121565 71909
rect 121499 71844 121500 71908
rect 121564 71844 121565 71908
rect 121499 71843 121565 71844
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 121502 3365 121562 71843
rect 121686 3501 121746 71979
rect 122790 71770 122850 71979
rect 122971 71908 123037 71909
rect 122971 71844 122972 71908
rect 123036 71844 123037 71908
rect 122971 71843 123037 71844
rect 122606 71710 122850 71770
rect 122606 3637 122666 71710
rect 122974 6221 123034 71843
rect 123294 52954 123914 73000
rect 126099 72316 126165 72317
rect 126099 72252 126100 72316
rect 126164 72252 126165 72316
rect 126099 72251 126165 72252
rect 124627 72180 124693 72181
rect 124627 72116 124628 72180
rect 124692 72116 124693 72180
rect 124627 72115 124693 72116
rect 125915 72180 125981 72181
rect 125915 72116 125916 72180
rect 125980 72116 125981 72180
rect 125915 72115 125981 72116
rect 124259 72044 124325 72045
rect 124259 71980 124260 72044
rect 124324 71980 124325 72044
rect 124259 71979 124325 71980
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 122971 6220 123037 6221
rect 122971 6156 122972 6220
rect 123036 6156 123037 6220
rect 122971 6155 123037 6156
rect 122603 3636 122669 3637
rect 122603 3572 122604 3636
rect 122668 3572 122669 3636
rect 122603 3571 122669 3572
rect 121683 3500 121749 3501
rect 121683 3436 121684 3500
rect 121748 3436 121749 3500
rect 121683 3435 121749 3436
rect 121499 3364 121565 3365
rect 121499 3300 121500 3364
rect 121564 3300 121565 3364
rect 121499 3299 121565 3300
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 -3226 123914 16398
rect 124262 4861 124322 71979
rect 124443 71908 124509 71909
rect 124443 71844 124444 71908
rect 124508 71844 124509 71908
rect 124443 71843 124509 71844
rect 124446 9077 124506 71843
rect 124443 9076 124509 9077
rect 124443 9012 124444 9076
rect 124508 9012 124509 9076
rect 124443 9011 124509 9012
rect 124630 8941 124690 72115
rect 125547 72044 125613 72045
rect 125547 71980 125548 72044
rect 125612 71980 125613 72044
rect 125547 71979 125613 71980
rect 124627 8940 124693 8941
rect 124627 8876 124628 8940
rect 124692 8876 124693 8940
rect 124627 8875 124693 8876
rect 124259 4860 124325 4861
rect 124259 4796 124260 4860
rect 124324 4796 124325 4860
rect 124259 4795 124325 4796
rect 125550 3773 125610 71979
rect 125731 71908 125797 71909
rect 125731 71844 125732 71908
rect 125796 71844 125797 71908
rect 125731 71843 125797 71844
rect 125734 6493 125794 71843
rect 125731 6492 125797 6493
rect 125731 6428 125732 6492
rect 125796 6428 125797 6492
rect 125731 6427 125797 6428
rect 125918 6357 125978 72115
rect 126102 9213 126162 72251
rect 127203 72044 127269 72045
rect 127203 71980 127204 72044
rect 127268 71980 127269 72044
rect 127203 71979 127269 71980
rect 127019 71908 127085 71909
rect 127019 71844 127020 71908
rect 127084 71844 127085 71908
rect 127019 71843 127085 71844
rect 126099 9212 126165 9213
rect 126099 9148 126100 9212
rect 126164 9148 126165 9212
rect 126099 9147 126165 9148
rect 127022 7581 127082 71843
rect 127206 10301 127266 71979
rect 127794 57454 128414 73000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127203 10300 127269 10301
rect 127203 10236 127204 10300
rect 127268 10236 127269 10300
rect 127203 10235 127269 10236
rect 127019 7580 127085 7581
rect 127019 7516 127020 7580
rect 127084 7516 127085 7580
rect 127019 7515 127085 7516
rect 125915 6356 125981 6357
rect 125915 6292 125916 6356
rect 125980 6292 125981 6356
rect 125915 6291 125981 6292
rect 125547 3772 125613 3773
rect 125547 3708 125548 3772
rect 125612 3708 125613 3772
rect 125547 3707 125613 3708
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 -4186 128414 20898
rect 128494 6930 128554 73067
rect 129043 72180 129109 72181
rect 129043 72116 129044 72180
rect 129108 72116 129109 72180
rect 129043 72115 129109 72116
rect 129963 72180 130029 72181
rect 129963 72116 129964 72180
rect 130028 72116 130029 72180
rect 129963 72115 130029 72116
rect 128859 72044 128925 72045
rect 128859 71980 128860 72044
rect 128924 71980 128925 72044
rect 128859 71979 128925 71980
rect 128675 71908 128741 71909
rect 128675 71844 128676 71908
rect 128740 71844 128741 71908
rect 128675 71843 128741 71844
rect 128678 7853 128738 71843
rect 128675 7852 128741 7853
rect 128675 7788 128676 7852
rect 128740 7788 128741 7852
rect 128675 7787 128741 7788
rect 128862 7717 128922 71979
rect 129046 10437 129106 72115
rect 129779 71908 129845 71909
rect 129779 71844 129780 71908
rect 129844 71844 129845 71908
rect 129779 71843 129845 71844
rect 129043 10436 129109 10437
rect 129043 10372 129044 10436
rect 129108 10372 129109 10436
rect 129043 10371 129109 10372
rect 128859 7716 128925 7717
rect 128859 7652 128860 7716
rect 128924 7652 128925 7716
rect 128859 7651 128925 7652
rect 128494 6870 128738 6930
rect 128678 4997 128738 6870
rect 129782 6629 129842 71843
rect 129966 9349 130026 72115
rect 130147 72044 130213 72045
rect 130147 71980 130148 72044
rect 130212 71980 130213 72044
rect 130147 71979 130213 71980
rect 131067 72044 131133 72045
rect 131067 71980 131068 72044
rect 131132 71980 131133 72044
rect 131067 71979 131133 71980
rect 131803 72044 131869 72045
rect 131803 71980 131804 72044
rect 131868 71980 131869 72044
rect 131803 71979 131869 71980
rect 130150 9485 130210 71979
rect 130147 9484 130213 9485
rect 130147 9420 130148 9484
rect 130212 9420 130213 9484
rect 130147 9419 130213 9420
rect 129963 9348 130029 9349
rect 129963 9284 129964 9348
rect 130028 9284 130029 9348
rect 129963 9283 130029 9284
rect 129779 6628 129845 6629
rect 129779 6564 129780 6628
rect 129844 6564 129845 6628
rect 129779 6563 129845 6564
rect 128675 4996 128741 4997
rect 128675 4932 128676 4996
rect 128740 4932 128741 4996
rect 128675 4931 128741 4932
rect 131070 3501 131130 71979
rect 131251 71908 131317 71909
rect 131251 71844 131252 71908
rect 131316 71844 131317 71908
rect 131251 71843 131317 71844
rect 131254 3637 131314 71843
rect 131806 3637 131866 71979
rect 131987 71908 132053 71909
rect 131987 71844 131988 71908
rect 132052 71844 132053 71908
rect 131987 71843 132053 71844
rect 131251 3636 131317 3637
rect 131251 3572 131252 3636
rect 131316 3572 131317 3636
rect 131251 3571 131317 3572
rect 131803 3636 131869 3637
rect 131803 3572 131804 3636
rect 131868 3572 131869 3636
rect 131803 3571 131869 3572
rect 131990 3501 132050 71843
rect 132294 61954 132914 73000
rect 133275 72180 133341 72181
rect 133275 72116 133276 72180
rect 133340 72116 133341 72180
rect 133275 72115 133341 72116
rect 134747 72180 134813 72181
rect 134747 72116 134748 72180
rect 134812 72116 134813 72180
rect 134747 72115 134813 72116
rect 135851 72180 135917 72181
rect 135851 72116 135852 72180
rect 135916 72116 135917 72180
rect 135851 72115 135917 72116
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 131067 3500 131133 3501
rect 131067 3436 131068 3500
rect 131132 3436 131133 3500
rect 131067 3435 131133 3436
rect 131987 3500 132053 3501
rect 131987 3436 131988 3500
rect 132052 3436 132053 3500
rect 131987 3435 132053 3436
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 -5146 132914 25398
rect 133278 4861 133338 72115
rect 133459 72044 133525 72045
rect 133459 71980 133460 72044
rect 133524 71980 133525 72044
rect 133459 71979 133525 71980
rect 133462 4997 133522 71979
rect 133643 71908 133709 71909
rect 133643 71844 133644 71908
rect 133708 71844 133709 71908
rect 133643 71843 133709 71844
rect 133459 4996 133525 4997
rect 133459 4932 133460 4996
rect 133524 4932 133525 4996
rect 133459 4931 133525 4932
rect 133275 4860 133341 4861
rect 133275 4796 133276 4860
rect 133340 4796 133341 4860
rect 133275 4795 133341 4796
rect 133646 3365 133706 71843
rect 134750 32741 134810 72115
rect 134931 72044 134997 72045
rect 134931 71980 134932 72044
rect 134996 71980 134997 72044
rect 134931 71979 134997 71980
rect 134747 32740 134813 32741
rect 134747 32676 134748 32740
rect 134812 32676 134813 32740
rect 134747 32675 134813 32676
rect 134934 25669 134994 71979
rect 135115 71908 135181 71909
rect 135115 71844 135116 71908
rect 135180 71844 135181 71908
rect 135115 71843 135181 71844
rect 134931 25668 134997 25669
rect 134931 25604 134932 25668
rect 134996 25604 134997 25668
rect 134931 25603 134997 25604
rect 135118 8125 135178 71843
rect 135854 32469 135914 72115
rect 136219 72044 136285 72045
rect 136219 71980 136220 72044
rect 136284 71980 136285 72044
rect 136219 71979 136285 71980
rect 136035 71908 136101 71909
rect 136035 71844 136036 71908
rect 136100 71844 136101 71908
rect 136035 71843 136101 71844
rect 136038 32605 136098 71843
rect 136035 32604 136101 32605
rect 136035 32540 136036 32604
rect 136100 32540 136101 32604
rect 136035 32539 136101 32540
rect 135851 32468 135917 32469
rect 135851 32404 135852 32468
rect 135916 32404 135917 32468
rect 135851 32403 135917 32404
rect 136222 27165 136282 71979
rect 136403 71908 136469 71909
rect 136403 71844 136404 71908
rect 136468 71844 136469 71908
rect 136403 71843 136469 71844
rect 136219 27164 136285 27165
rect 136219 27100 136220 27164
rect 136284 27100 136285 27164
rect 136219 27099 136285 27100
rect 135115 8124 135181 8125
rect 135115 8060 135116 8124
rect 135180 8060 135181 8124
rect 135115 8059 135181 8060
rect 136406 4725 136466 71843
rect 136794 66454 137414 73000
rect 138979 72180 139045 72181
rect 138979 72116 138980 72180
rect 139044 72116 139045 72180
rect 138979 72115 139045 72116
rect 140083 72180 140149 72181
rect 140083 72116 140084 72180
rect 140148 72116 140149 72180
rect 140083 72115 140149 72116
rect 137691 72044 137757 72045
rect 137691 71980 137692 72044
rect 137756 71980 137757 72044
rect 137691 71979 137757 71980
rect 138795 72044 138861 72045
rect 138795 71980 138796 72044
rect 138860 71980 138861 72044
rect 138795 71979 138861 71980
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 137694 34101 137754 71979
rect 137875 71908 137941 71909
rect 137875 71844 137876 71908
rect 137940 71844 137941 71908
rect 137875 71843 137941 71844
rect 138611 71908 138677 71909
rect 138611 71844 138612 71908
rect 138676 71844 138677 71908
rect 138611 71843 138677 71844
rect 137691 34100 137757 34101
rect 137691 34036 137692 34100
rect 137756 34036 137757 34100
rect 137691 34035 137757 34036
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136403 4724 136469 4725
rect 136403 4660 136404 4724
rect 136468 4660 136469 4724
rect 136403 4659 136469 4660
rect 133643 3364 133709 3365
rect 133643 3300 133644 3364
rect 133708 3300 133709 3364
rect 133643 3299 133709 3300
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 -6106 137414 29898
rect 137878 12205 137938 71843
rect 138614 20229 138674 71843
rect 138611 20228 138677 20229
rect 138611 20164 138612 20228
rect 138676 20164 138677 20228
rect 138611 20163 138677 20164
rect 138798 12885 138858 71979
rect 138795 12884 138861 12885
rect 138795 12820 138796 12884
rect 138860 12820 138861 12884
rect 138795 12819 138861 12820
rect 137875 12204 137941 12205
rect 137875 12140 137876 12204
rect 137940 12140 137941 12204
rect 137875 12139 137941 12140
rect 138982 6901 139042 72115
rect 139163 71908 139229 71909
rect 139163 71844 139164 71908
rect 139228 71844 139229 71908
rect 139163 71843 139229 71844
rect 138979 6900 139045 6901
rect 138979 6836 138980 6900
rect 139044 6836 139045 6900
rect 138979 6835 139045 6836
rect 139166 6085 139226 71843
rect 140086 33965 140146 72115
rect 140267 72044 140333 72045
rect 140267 71980 140268 72044
rect 140332 71980 140333 72044
rect 140267 71979 140333 71980
rect 140819 72044 140885 72045
rect 140819 71980 140820 72044
rect 140884 71980 140885 72044
rect 140819 71979 140885 71980
rect 140083 33964 140149 33965
rect 140083 33900 140084 33964
rect 140148 33900 140149 33964
rect 140083 33899 140149 33900
rect 140270 20093 140330 71979
rect 140451 71908 140517 71909
rect 140451 71844 140452 71908
rect 140516 71844 140517 71908
rect 140451 71843 140517 71844
rect 140635 71908 140701 71909
rect 140635 71844 140636 71908
rect 140700 71844 140701 71908
rect 140635 71843 140701 71844
rect 140267 20092 140333 20093
rect 140267 20028 140268 20092
rect 140332 20028 140333 20092
rect 140267 20027 140333 20028
rect 140454 13701 140514 71843
rect 140451 13700 140517 13701
rect 140451 13636 140452 13700
rect 140516 13636 140517 13700
rect 140451 13635 140517 13636
rect 140638 6765 140698 71843
rect 140822 33829 140882 71979
rect 141003 71908 141069 71909
rect 141003 71844 141004 71908
rect 141068 71844 141069 71908
rect 141003 71843 141069 71844
rect 140819 33828 140885 33829
rect 140819 33764 140820 33828
rect 140884 33764 140885 33828
rect 140819 33763 140885 33764
rect 141006 15197 141066 71843
rect 141294 70954 141914 73000
rect 142843 72180 142909 72181
rect 142843 72116 142844 72180
rect 142908 72116 142909 72180
rect 142843 72115 142909 72116
rect 144131 72180 144197 72181
rect 144131 72116 144132 72180
rect 144196 72116 144197 72180
rect 144131 72115 144197 72116
rect 145235 72180 145301 72181
rect 145235 72116 145236 72180
rect 145300 72116 145301 72180
rect 145235 72115 145301 72116
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141003 15196 141069 15197
rect 141003 15132 141004 15196
rect 141068 15132 141069 15196
rect 141003 15131 141069 15132
rect 140635 6764 140701 6765
rect 140635 6700 140636 6764
rect 140700 6700 140701 6764
rect 140635 6699 140701 6700
rect 139163 6084 139229 6085
rect 139163 6020 139164 6084
rect 139228 6020 139229 6084
rect 139163 6019 139229 6020
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 -7066 141914 34398
rect 142846 27029 142906 72115
rect 143027 72044 143093 72045
rect 143027 71980 143028 72044
rect 143092 71980 143093 72044
rect 143027 71979 143093 71980
rect 142843 27028 142909 27029
rect 142843 26964 142844 27028
rect 142908 26964 142909 27028
rect 142843 26963 142909 26964
rect 143030 13565 143090 71979
rect 143211 71908 143277 71909
rect 143211 71844 143212 71908
rect 143276 71844 143277 71908
rect 143211 71843 143277 71844
rect 143395 71908 143461 71909
rect 143395 71844 143396 71908
rect 143460 71844 143461 71908
rect 143395 71843 143461 71844
rect 143027 13564 143093 13565
rect 143027 13500 143028 13564
rect 143092 13500 143093 13564
rect 143027 13499 143093 13500
rect 143214 7989 143274 71843
rect 143211 7988 143277 7989
rect 143211 7924 143212 7988
rect 143276 7924 143277 7988
rect 143211 7923 143277 7924
rect 143398 7853 143458 71843
rect 144134 35325 144194 72115
rect 144499 72044 144565 72045
rect 144499 71980 144500 72044
rect 144564 71980 144565 72044
rect 144499 71979 144565 71980
rect 144315 71908 144381 71909
rect 144315 71844 144316 71908
rect 144380 71844 144381 71908
rect 144315 71843 144381 71844
rect 144131 35324 144197 35325
rect 144131 35260 144132 35324
rect 144196 35260 144197 35324
rect 144131 35259 144197 35260
rect 144318 16285 144378 71843
rect 144315 16284 144381 16285
rect 144315 16220 144316 16284
rect 144380 16220 144381 16284
rect 144315 16219 144381 16220
rect 144502 15061 144562 71979
rect 144683 71908 144749 71909
rect 144683 71844 144684 71908
rect 144748 71844 144749 71908
rect 144683 71843 144749 71844
rect 144499 15060 144565 15061
rect 144499 14996 144500 15060
rect 144564 14996 144565 15060
rect 144499 14995 144565 14996
rect 144686 9077 144746 71843
rect 145238 29613 145298 72115
rect 145419 72044 145485 72045
rect 145419 71980 145420 72044
rect 145484 71980 145485 72044
rect 145419 71979 145485 71980
rect 145235 29612 145301 29613
rect 145235 29548 145236 29612
rect 145300 29548 145301 29612
rect 145235 29547 145301 29548
rect 145422 17645 145482 71979
rect 145603 71908 145669 71909
rect 145603 71844 145604 71908
rect 145668 71844 145669 71908
rect 145603 71843 145669 71844
rect 145419 17644 145485 17645
rect 145419 17580 145420 17644
rect 145484 17580 145485 17644
rect 145419 17579 145485 17580
rect 145606 14925 145666 71843
rect 145794 39454 146414 73000
rect 148363 72860 148429 72861
rect 148363 72796 148364 72860
rect 148428 72796 148429 72860
rect 148363 72795 148429 72796
rect 149651 72860 149717 72861
rect 149651 72796 149652 72860
rect 149716 72796 149717 72860
rect 149651 72795 149717 72796
rect 146891 72316 146957 72317
rect 146891 72252 146892 72316
rect 146956 72252 146957 72316
rect 146891 72251 146957 72252
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145603 14924 145669 14925
rect 145603 14860 145604 14924
rect 145668 14860 145669 14924
rect 145603 14859 145669 14860
rect 144683 9076 144749 9077
rect 144683 9012 144684 9076
rect 144748 9012 144749 9076
rect 144683 9011 144749 9012
rect 143395 7852 143461 7853
rect 143395 7788 143396 7852
rect 143460 7788 143461 7852
rect 143395 7787 143461 7788
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 3454 146414 38898
rect 146894 35189 146954 72251
rect 147075 72180 147141 72181
rect 147075 72116 147076 72180
rect 147140 72116 147141 72180
rect 147075 72115 147141 72116
rect 146891 35188 146957 35189
rect 146891 35124 146892 35188
rect 146956 35124 146957 35188
rect 146891 35123 146957 35124
rect 147078 14789 147138 72115
rect 147259 72044 147325 72045
rect 147259 71980 147260 72044
rect 147324 71980 147325 72044
rect 147259 71979 147325 71980
rect 147075 14788 147141 14789
rect 147075 14724 147076 14788
rect 147140 14724 147141 14788
rect 147075 14723 147141 14724
rect 147262 10301 147322 71979
rect 147443 71908 147509 71909
rect 147443 71844 147444 71908
rect 147508 71844 147509 71908
rect 147443 71843 147509 71844
rect 147446 10437 147506 71843
rect 148366 21453 148426 72795
rect 148731 72724 148797 72725
rect 148731 72660 148732 72724
rect 148796 72660 148797 72724
rect 148731 72659 148797 72660
rect 148915 72724 148981 72725
rect 148915 72660 148916 72724
rect 148980 72660 148981 72724
rect 148915 72659 148981 72660
rect 148547 72452 148613 72453
rect 148547 72388 148548 72452
rect 148612 72388 148613 72452
rect 148547 72387 148613 72388
rect 148363 21452 148429 21453
rect 148363 21388 148364 21452
rect 148428 21388 148429 21452
rect 148363 21387 148429 21388
rect 148550 16149 148610 72387
rect 148547 16148 148613 16149
rect 148547 16084 148548 16148
rect 148612 16084 148613 16148
rect 148547 16083 148613 16084
rect 148734 12069 148794 72659
rect 148731 12068 148797 12069
rect 148731 12004 148732 12068
rect 148796 12004 148797 12068
rect 148731 12003 148797 12004
rect 148918 11933 148978 72659
rect 149467 72588 149533 72589
rect 149467 72524 149468 72588
rect 149532 72524 149533 72588
rect 149467 72523 149533 72524
rect 149470 26893 149530 72523
rect 149467 26892 149533 26893
rect 149467 26828 149468 26892
rect 149532 26828 149533 26892
rect 149467 26827 149533 26828
rect 149654 13293 149714 72795
rect 150019 72724 150085 72725
rect 150019 72660 150020 72724
rect 150084 72660 150085 72724
rect 150019 72659 150085 72660
rect 149835 72452 149901 72453
rect 149835 72388 149836 72452
rect 149900 72388 149901 72452
rect 149835 72387 149901 72388
rect 149838 13429 149898 72387
rect 149835 13428 149901 13429
rect 149835 13364 149836 13428
rect 149900 13364 149901 13428
rect 149835 13363 149901 13364
rect 149651 13292 149717 13293
rect 149651 13228 149652 13292
rect 149716 13228 149717 13292
rect 149651 13227 149717 13228
rect 148915 11932 148981 11933
rect 148915 11868 148916 11932
rect 148980 11868 148981 11932
rect 148915 11867 148981 11868
rect 150022 11797 150082 72659
rect 150294 43954 150914 73000
rect 152411 72996 152477 72997
rect 152411 72932 152412 72996
rect 152476 72932 152477 72996
rect 152411 72931 152477 72932
rect 151307 72860 151373 72861
rect 151307 72796 151308 72860
rect 151372 72796 151373 72860
rect 151307 72795 151373 72796
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150019 11796 150085 11797
rect 150019 11732 150020 11796
rect 150084 11732 150085 11796
rect 150019 11731 150085 11732
rect 147443 10436 147509 10437
rect 147443 10372 147444 10436
rect 147508 10372 147509 10436
rect 147443 10371 147509 10372
rect 147259 10300 147325 10301
rect 147259 10236 147260 10300
rect 147324 10236 147325 10300
rect 147259 10235 147325 10236
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 7954 150914 43398
rect 151310 24445 151370 72795
rect 151675 72724 151741 72725
rect 151675 72660 151676 72724
rect 151740 72660 151741 72724
rect 151675 72659 151741 72660
rect 151491 72452 151557 72453
rect 151491 72388 151492 72452
rect 151556 72388 151557 72452
rect 151491 72387 151557 72388
rect 151307 24444 151373 24445
rect 151307 24380 151308 24444
rect 151372 24380 151373 24444
rect 151307 24379 151373 24380
rect 151494 14653 151554 72387
rect 151491 14652 151557 14653
rect 151491 14588 151492 14652
rect 151556 14588 151557 14652
rect 151491 14587 151557 14588
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 151678 6629 151738 72659
rect 152414 16013 152474 72931
rect 152779 72860 152845 72861
rect 152779 72796 152780 72860
rect 152844 72796 152845 72860
rect 152779 72795 152845 72796
rect 154435 72860 154501 72861
rect 154435 72796 154436 72860
rect 154500 72796 154501 72860
rect 154435 72795 154501 72796
rect 152595 72588 152661 72589
rect 152595 72524 152596 72588
rect 152660 72524 152661 72588
rect 152595 72523 152661 72524
rect 152411 16012 152477 16013
rect 152411 15948 152412 16012
rect 152476 15948 152477 16012
rect 152411 15947 152477 15948
rect 152598 14517 152658 72523
rect 152595 14516 152661 14517
rect 152595 14452 152596 14516
rect 152660 14452 152661 14516
rect 152595 14451 152661 14452
rect 152782 11661 152842 72795
rect 152963 72724 153029 72725
rect 152963 72660 152964 72724
rect 153028 72660 153029 72724
rect 152963 72659 153029 72660
rect 154251 72724 154317 72725
rect 154251 72660 154252 72724
rect 154316 72660 154317 72724
rect 154251 72659 154317 72660
rect 152779 11660 152845 11661
rect 152779 11596 152780 11660
rect 152844 11596 152845 11660
rect 152779 11595 152845 11596
rect 151675 6628 151741 6629
rect 151675 6564 151676 6628
rect 151740 6564 151741 6628
rect 151675 6563 151741 6564
rect 152966 5541 153026 72659
rect 153883 72588 153949 72589
rect 153883 72524 153884 72588
rect 153948 72524 153949 72588
rect 153883 72523 153949 72524
rect 153886 17373 153946 72523
rect 154067 72452 154133 72453
rect 154067 72388 154068 72452
rect 154132 72388 154133 72452
rect 154067 72387 154133 72388
rect 154070 17509 154130 72387
rect 154067 17508 154133 17509
rect 154067 17444 154068 17508
rect 154132 17444 154133 17508
rect 154067 17443 154133 17444
rect 153883 17372 153949 17373
rect 153883 17308 153884 17372
rect 153948 17308 153949 17372
rect 153883 17307 153949 17308
rect 154254 15877 154314 72659
rect 154251 15876 154317 15877
rect 154251 15812 154252 15876
rect 154316 15812 154317 15876
rect 154251 15811 154317 15812
rect 154438 13157 154498 72795
rect 154794 48454 155414 73000
rect 157011 72860 157077 72861
rect 157011 72796 157012 72860
rect 157076 72796 157077 72860
rect 157011 72795 157077 72796
rect 158483 72860 158549 72861
rect 158483 72796 158484 72860
rect 158548 72796 158549 72860
rect 158483 72795 158549 72796
rect 158851 72860 158917 72861
rect 158851 72796 158852 72860
rect 158916 72796 158917 72860
rect 158851 72795 158917 72796
rect 155723 72724 155789 72725
rect 155723 72660 155724 72724
rect 155788 72660 155789 72724
rect 155723 72659 155789 72660
rect 156827 72724 156893 72725
rect 156827 72660 156828 72724
rect 156892 72660 156893 72724
rect 156827 72659 156893 72660
rect 155539 72452 155605 72453
rect 155539 72388 155540 72452
rect 155604 72388 155605 72452
rect 155539 72387 155605 72388
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154435 13156 154501 13157
rect 154435 13092 154436 13156
rect 154500 13092 154501 13156
rect 154435 13091 154501 13092
rect 154794 12454 155414 47898
rect 155542 22949 155602 72387
rect 155539 22948 155605 22949
rect 155539 22884 155540 22948
rect 155604 22884 155605 22948
rect 155539 22883 155605 22884
rect 155726 17237 155786 72659
rect 156643 72588 156709 72589
rect 156643 72524 156644 72588
rect 156708 72524 156709 72588
rect 156643 72523 156709 72524
rect 156646 25533 156706 72523
rect 156643 25532 156709 25533
rect 156643 25468 156644 25532
rect 156708 25468 156709 25532
rect 156643 25467 156709 25468
rect 156830 22813 156890 72659
rect 156827 22812 156893 22813
rect 156827 22748 156828 22812
rect 156892 22748 156893 22812
rect 156827 22747 156893 22748
rect 157014 18869 157074 72795
rect 157195 72724 157261 72725
rect 157195 72660 157196 72724
rect 157260 72660 157261 72724
rect 157195 72659 157261 72660
rect 157011 18868 157077 18869
rect 157011 18804 157012 18868
rect 157076 18804 157077 18868
rect 157011 18803 157077 18804
rect 157198 18733 157258 72659
rect 158299 72588 158365 72589
rect 158299 72524 158300 72588
rect 158364 72524 158365 72588
rect 158299 72523 158365 72524
rect 158115 72452 158181 72453
rect 158115 72388 158116 72452
rect 158180 72388 158181 72452
rect 158115 72387 158181 72388
rect 158118 31109 158178 72387
rect 158115 31108 158181 31109
rect 158115 31044 158116 31108
rect 158180 31044 158181 31108
rect 158115 31043 158181 31044
rect 158302 21317 158362 72523
rect 158299 21316 158365 21317
rect 158299 21252 158300 21316
rect 158364 21252 158365 21316
rect 158299 21251 158365 21252
rect 158486 19957 158546 72795
rect 158667 72724 158733 72725
rect 158667 72660 158668 72724
rect 158732 72660 158733 72724
rect 158667 72659 158733 72660
rect 158670 65517 158730 72659
rect 158667 65516 158733 65517
rect 158667 65452 158668 65516
rect 158732 65452 158733 65516
rect 158667 65451 158733 65452
rect 158854 30973 158914 72795
rect 159035 72724 159101 72725
rect 159035 72660 159036 72724
rect 159100 72660 159101 72724
rect 159035 72659 159101 72660
rect 158851 30972 158917 30973
rect 158851 30908 158852 30972
rect 158916 30908 158917 30972
rect 158851 30907 158917 30908
rect 158483 19956 158549 19957
rect 158483 19892 158484 19956
rect 158548 19892 158549 19956
rect 158483 19891 158549 19892
rect 157195 18732 157261 18733
rect 157195 18668 157196 18732
rect 157260 18668 157261 18732
rect 157195 18667 157261 18668
rect 155723 17236 155789 17237
rect 155723 17172 155724 17236
rect 155788 17172 155789 17236
rect 155723 17171 155789 17172
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 152963 5540 153029 5541
rect 152963 5476 152964 5540
rect 153028 5476 153029 5540
rect 152963 5475 153029 5476
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 -2266 155414 11898
rect 159038 3909 159098 72659
rect 159294 52954 159914 73000
rect 160875 72860 160941 72861
rect 160875 72796 160876 72860
rect 160940 72796 160941 72860
rect 160875 72795 160941 72796
rect 160691 72588 160757 72589
rect 160691 72524 160692 72588
rect 160756 72524 160757 72588
rect 160691 72523 160757 72524
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 160694 22677 160754 72523
rect 160691 22676 160757 22677
rect 160691 22612 160692 22676
rect 160756 22612 160757 22676
rect 160691 22611 160757 22612
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159035 3908 159101 3909
rect 159035 3844 159036 3908
rect 159100 3844 159101 3908
rect 159035 3843 159101 3844
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 -3226 159914 16398
rect 160878 13021 160938 72795
rect 161059 72724 161125 72725
rect 161059 72660 161060 72724
rect 161124 72660 161125 72724
rect 161059 72659 161125 72660
rect 161243 72724 161309 72725
rect 161243 72660 161244 72724
rect 161308 72660 161309 72724
rect 161243 72659 161309 72660
rect 160875 13020 160941 13021
rect 160875 12956 160876 13020
rect 160940 12956 160941 13020
rect 160875 12955 160941 12956
rect 161062 5405 161122 72659
rect 161059 5404 161125 5405
rect 161059 5340 161060 5404
rect 161124 5340 161125 5404
rect 161059 5339 161125 5340
rect 161246 5269 161306 72659
rect 161614 72589 161674 74699
rect 162347 72860 162413 72861
rect 162347 72796 162348 72860
rect 162412 72796 162413 72860
rect 162347 72795 162413 72796
rect 163451 72860 163517 72861
rect 163451 72796 163452 72860
rect 163516 72796 163517 72860
rect 163451 72795 163517 72796
rect 161611 72588 161677 72589
rect 161611 72524 161612 72588
rect 161676 72524 161677 72588
rect 161611 72523 161677 72524
rect 162163 72452 162229 72453
rect 162163 72388 162164 72452
rect 162228 72388 162229 72452
rect 162163 72387 162229 72388
rect 162166 24309 162226 72387
rect 162163 24308 162229 24309
rect 162163 24244 162164 24308
rect 162228 24244 162229 24308
rect 162163 24243 162229 24244
rect 162350 18597 162410 72795
rect 162531 72724 162597 72725
rect 162531 72660 162532 72724
rect 162596 72660 162597 72724
rect 162531 72659 162597 72660
rect 162715 72724 162781 72725
rect 162715 72660 162716 72724
rect 162780 72660 162781 72724
rect 162715 72659 162781 72660
rect 162347 18596 162413 18597
rect 162347 18532 162348 18596
rect 162412 18532 162413 18596
rect 162347 18531 162413 18532
rect 162534 6493 162594 72659
rect 162531 6492 162597 6493
rect 162531 6428 162532 6492
rect 162596 6428 162597 6492
rect 162531 6427 162597 6428
rect 162718 6357 162778 72659
rect 163267 72588 163333 72589
rect 163267 72524 163268 72588
rect 163332 72524 163333 72588
rect 163267 72523 163333 72524
rect 163270 31245 163330 72523
rect 163267 31244 163333 31245
rect 163267 31180 163268 31244
rect 163332 31180 163333 31244
rect 163267 31179 163333 31180
rect 163454 24173 163514 72795
rect 163635 72724 163701 72725
rect 163635 72660 163636 72724
rect 163700 72660 163701 72724
rect 163635 72659 163701 72660
rect 163451 24172 163517 24173
rect 163451 24108 163452 24172
rect 163516 24108 163517 24172
rect 163451 24107 163517 24108
rect 162715 6356 162781 6357
rect 162715 6292 162716 6356
rect 162780 6292 162781 6356
rect 162715 6291 162781 6292
rect 161243 5268 161309 5269
rect 161243 5204 161244 5268
rect 161308 5204 161309 5268
rect 161243 5203 161309 5204
rect 163638 5133 163698 72659
rect 163794 57454 164414 73000
rect 164742 71365 164802 74699
rect 164923 74220 164989 74221
rect 164923 74156 164924 74220
rect 164988 74156 164989 74220
rect 164923 74155 164989 74156
rect 164926 72861 164986 74155
rect 166763 73404 166829 73405
rect 166763 73340 166764 73404
rect 166828 73340 166829 73404
rect 166763 73339 166829 73340
rect 165843 73132 165909 73133
rect 165843 73068 165844 73132
rect 165908 73068 165909 73132
rect 165843 73067 165909 73068
rect 164923 72860 164989 72861
rect 164923 72796 164924 72860
rect 164988 72796 164989 72860
rect 164923 72795 164989 72796
rect 165291 72860 165357 72861
rect 165291 72796 165292 72860
rect 165356 72796 165357 72860
rect 165291 72795 165357 72796
rect 164923 72724 164989 72725
rect 164923 72660 164924 72724
rect 164988 72660 164989 72724
rect 164923 72659 164989 72660
rect 164739 71364 164805 71365
rect 164739 71300 164740 71364
rect 164804 71300 164805 71364
rect 164739 71299 164805 71300
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163635 5132 163701 5133
rect 163635 5068 163636 5132
rect 163700 5068 163701 5132
rect 163635 5067 163701 5068
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 -4186 164414 20898
rect 164926 7717 164986 72659
rect 165107 72588 165173 72589
rect 165107 72524 165108 72588
rect 165172 72524 165173 72588
rect 165107 72523 165173 72524
rect 164923 7716 164989 7717
rect 164923 7652 164924 7716
rect 164988 7652 164989 7716
rect 164923 7651 164989 7652
rect 165110 7581 165170 72523
rect 165107 7580 165173 7581
rect 165107 7516 165108 7580
rect 165172 7516 165173 7580
rect 165107 7515 165173 7516
rect 165294 4997 165354 72795
rect 165475 72724 165541 72725
rect 165475 72660 165476 72724
rect 165540 72660 165541 72724
rect 165475 72659 165541 72660
rect 165291 4996 165357 4997
rect 165291 4932 165292 4996
rect 165356 4932 165357 4996
rect 165291 4931 165357 4932
rect 165478 4861 165538 72659
rect 165846 71229 165906 73067
rect 166579 72860 166645 72861
rect 166579 72796 166580 72860
rect 166644 72796 166645 72860
rect 166579 72795 166645 72796
rect 166395 72724 166461 72725
rect 166395 72660 166396 72724
rect 166460 72660 166461 72724
rect 166395 72659 166461 72660
rect 165843 71228 165909 71229
rect 165843 71164 165844 71228
rect 165908 71164 165909 71228
rect 165843 71163 165909 71164
rect 166398 8941 166458 72659
rect 166395 8940 166461 8941
rect 166395 8876 166396 8940
rect 166460 8876 166461 8940
rect 166395 8875 166461 8876
rect 166582 6221 166642 72795
rect 166579 6220 166645 6221
rect 166579 6156 166580 6220
rect 166644 6156 166645 6220
rect 166579 6155 166645 6156
rect 165475 4860 165541 4861
rect 165475 4796 165476 4860
rect 165540 4796 165541 4860
rect 165475 4795 165541 4796
rect 166766 3365 166826 73339
rect 167502 4045 167562 74835
rect 169526 74765 169586 75243
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 169523 74764 169589 74765
rect 169523 74700 169524 74764
rect 169588 74700 169589 74764
rect 169523 74699 169589 74700
rect 167867 71228 167933 71229
rect 167867 71164 167868 71228
rect 167932 71164 167933 71228
rect 167867 71163 167933 71164
rect 167683 70140 167749 70141
rect 167683 70076 167684 70140
rect 167748 70076 167749 70140
rect 167683 70075 167749 70076
rect 167499 4044 167565 4045
rect 167499 3980 167500 4044
rect 167564 3980 167565 4044
rect 167499 3979 167565 3980
rect 167686 3501 167746 70075
rect 167870 3637 167930 71163
rect 168294 61954 168914 73000
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 167867 3636 167933 3637
rect 167867 3572 167868 3636
rect 167932 3572 167933 3636
rect 167867 3571 167933 3572
rect 167683 3500 167749 3501
rect 167683 3436 167684 3500
rect 167748 3436 167749 3500
rect 167683 3435 167749 3436
rect 166763 3364 166829 3365
rect 166763 3300 166764 3364
rect 166828 3300 166829 3364
rect 166763 3299 166829 3300
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 66454 173414 73000
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 70954 177914 73000
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 223954 186914 228484
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 228453 191414 228484
rect 190794 228217 190826 228453
rect 191062 228217 191146 228453
rect 191382 228217 191414 228453
rect 190794 228133 191414 228217
rect 190794 227897 190826 228133
rect 191062 227897 191146 228133
rect 191382 227897 191414 228133
rect 190794 192454 191414 227897
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 196954 195914 228484
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 201454 200414 228484
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 205954 204914 228484
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 210454 209414 228484
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 214954 213914 228484
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 219454 218414 228484
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 223954 222914 228484
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 228453 227414 228484
rect 226794 228217 226826 228453
rect 227062 228217 227146 228453
rect 227382 228217 227414 228453
rect 226794 228133 227414 228217
rect 226794 227897 226826 228133
rect 227062 227897 227146 228133
rect 227382 227897 227414 228133
rect 226794 192454 227414 227897
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 196954 231914 228484
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 201454 236414 228484
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 205954 240914 228484
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 210454 245414 228484
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 214954 249914 228484
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 219454 254414 228484
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 223954 258914 228484
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 228453 263414 228484
rect 262794 228217 262826 228453
rect 263062 228217 263146 228453
rect 263382 228217 263414 228453
rect 262794 228133 263414 228217
rect 262794 227897 262826 228133
rect 263062 227897 263146 228133
rect 263382 227897 263414 228133
rect 262794 192454 263414 227897
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 196954 267914 228484
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 201454 272414 228484
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 205954 276914 228484
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 210454 281414 228484
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 214954 285914 228484
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 219454 290414 228484
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 223954 294914 228484
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 228453 299414 228484
rect 298794 228217 298826 228453
rect 299062 228217 299146 228453
rect 299382 228217 299414 228453
rect 298794 228133 299414 228217
rect 298794 227897 298826 228133
rect 299062 227897 299146 228133
rect 299382 227897 299414 228133
rect 298794 192454 299414 227897
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 196954 303914 228484
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 201454 308414 228484
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 205954 312914 228484
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 210454 317414 228484
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 214954 321914 228484
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 219454 326414 228484
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 223954 330914 228484
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 228453 335414 228484
rect 334794 228217 334826 228453
rect 335062 228217 335146 228453
rect 335382 228217 335414 228453
rect 334794 228133 335414 228217
rect 334794 227897 334826 228133
rect 335062 227897 335146 228133
rect 335382 227897 335414 228133
rect 334794 192454 335414 227897
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 196954 339914 228484
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 201454 344414 228484
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 205954 348914 228484
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 210454 353414 228484
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 214954 357914 228484
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 219454 362414 228484
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 223954 366914 228484
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 228453 371414 228484
rect 370794 228217 370826 228453
rect 371062 228217 371146 228453
rect 371382 228217 371414 228453
rect 370794 228133 371414 228217
rect 370794 227897 370826 228133
rect 371062 227897 371146 228133
rect 371382 227897 371414 228133
rect 370794 192454 371414 227897
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 196954 375914 228484
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 201454 380414 228484
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 205954 384914 228484
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 210454 389414 228484
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 214954 393914 228484
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 396582 138685 396642 418235
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 248684 398414 254898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 396763 240140 396829 240141
rect 396763 240076 396764 240140
rect 396828 240076 396829 240140
rect 396763 240075 396829 240076
rect 396766 232389 396826 240075
rect 396947 240004 397013 240005
rect 396947 239940 396948 240004
rect 397012 239940 397013 240004
rect 396947 239939 397013 239940
rect 396763 232388 396829 232389
rect 396763 232324 396764 232388
rect 396828 232324 396829 232388
rect 396763 232323 396829 232324
rect 396950 231165 397010 239939
rect 396947 231164 397013 231165
rect 396947 231100 396948 231164
rect 397012 231100 397013 231164
rect 396947 231099 397013 231100
rect 397794 219454 398414 228484
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 396579 138684 396645 138685
rect 396579 138620 396580 138684
rect 396644 138620 396645 138684
rect 396579 138619 396645 138620
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 542675 699820 542741 699821
rect 542675 699756 542676 699820
rect 542740 699756 542741 699820
rect 542675 699755 542741 699756
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 542678 683130 542738 699755
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 320800 542414 326898
rect 542494 683070 542738 683130
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 291454 542414 300000
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 542494 151830 542554 683070
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 320800 546914 331398
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 320800 551414 335898
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 320800 555914 340398
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 320800 560414 344898
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 320800 564914 349398
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 320800 569414 353898
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 561300 318361 566100 318486
rect 561300 318125 561342 318361
rect 561578 318125 561662 318361
rect 561898 318125 561982 318361
rect 562218 318125 562302 318361
rect 562538 318125 562622 318361
rect 562858 318125 562942 318361
rect 563178 318125 563262 318361
rect 563498 318125 563582 318361
rect 563818 318125 563902 318361
rect 564138 318125 564222 318361
rect 564458 318125 564542 318361
rect 564778 318125 564862 318361
rect 565098 318125 565182 318361
rect 565418 318125 565502 318361
rect 565738 318125 565822 318361
rect 566058 318125 566100 318361
rect 561300 318000 566100 318125
rect 561300 313954 567300 313986
rect 561300 313718 561462 313954
rect 561698 313718 561782 313954
rect 562018 313718 562102 313954
rect 562338 313718 562422 313954
rect 562658 313718 562742 313954
rect 562978 313718 563062 313954
rect 563298 313718 563382 313954
rect 563618 313718 563702 313954
rect 563938 313718 564022 313954
rect 564258 313718 564342 313954
rect 564578 313718 564662 313954
rect 564898 313718 564982 313954
rect 565218 313718 565302 313954
rect 565538 313718 565622 313954
rect 565858 313718 565942 313954
rect 566178 313718 566262 313954
rect 566498 313718 566582 313954
rect 566818 313718 566902 313954
rect 567138 313718 567300 313954
rect 561300 313634 567300 313718
rect 561300 313398 561462 313634
rect 561698 313398 561782 313634
rect 562018 313398 562102 313634
rect 562338 313398 562422 313634
rect 562658 313398 562742 313634
rect 562978 313398 563062 313634
rect 563298 313398 563382 313634
rect 563618 313398 563702 313634
rect 563938 313398 564022 313634
rect 564258 313398 564342 313634
rect 564578 313398 564662 313634
rect 564898 313398 564982 313634
rect 565218 313398 565302 313634
rect 565538 313398 565622 313634
rect 565858 313398 565942 313634
rect 566178 313398 566262 313634
rect 566498 313398 566582 313634
rect 566818 313398 566902 313634
rect 567138 313398 567300 313634
rect 561300 313366 567300 313398
rect 546294 295954 546914 300000
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 542494 151770 542738 151830
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 542678 137325 542738 151770
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 542675 137324 542741 137325
rect 542675 137260 542676 137324
rect 542740 137260 542741 137324
rect 542675 137259 542741 137260
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 264454 551414 300000
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 268954 555914 300000
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 273454 560414 300000
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 277954 564914 300000
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 282454 569414 300000
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 580211 697236 580277 697237
rect 580211 697172 580212 697236
rect 580276 697172 580277 697236
rect 580211 697171 580277 697172
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 580214 74901 580274 697171
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 577794 39454 578414 74898
rect 580211 74900 580277 74901
rect 580211 74836 580212 74900
rect 580276 74836 580277 74900
rect 580211 74835 580277 74836
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 65342 246067 65578 246303
rect 65662 246067 65898 246303
rect 65982 246067 66218 246303
rect 66302 246067 66538 246303
rect 66622 246067 66858 246303
rect 66942 246067 67178 246303
rect 67262 246067 67498 246303
rect 67582 246067 67818 246303
rect 67902 246067 68138 246303
rect 68222 246067 68458 246303
rect 68542 246067 68778 246303
rect 68862 246067 69098 246303
rect 69182 246067 69418 246303
rect 69502 246067 69738 246303
rect 69822 246067 70058 246303
rect 65462 241717 65698 241953
rect 65782 241717 66018 241953
rect 66102 241717 66338 241953
rect 66422 241717 66658 241953
rect 66742 241717 66978 241953
rect 67062 241717 67298 241953
rect 67382 241717 67618 241953
rect 67702 241717 67938 241953
rect 68022 241717 68258 241953
rect 68342 241717 68578 241953
rect 68662 241717 68898 241953
rect 68982 241717 69218 241953
rect 69302 241717 69538 241953
rect 69622 241717 69858 241953
rect 69942 241717 70178 241953
rect 70262 241717 70498 241953
rect 70582 241717 70818 241953
rect 70902 241717 71138 241953
rect 65462 241397 65698 241633
rect 65782 241397 66018 241633
rect 66102 241397 66338 241633
rect 66422 241397 66658 241633
rect 66742 241397 66978 241633
rect 67062 241397 67298 241633
rect 67382 241397 67618 241633
rect 67702 241397 67938 241633
rect 68022 241397 68258 241633
rect 68342 241397 68578 241633
rect 68662 241397 68898 241633
rect 68982 241397 69218 241633
rect 69302 241397 69538 241633
rect 69622 241397 69858 241633
rect 69942 241397 70178 241633
rect 70262 241397 70498 241633
rect 70582 241397 70818 241633
rect 70902 241397 71138 241633
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 228217 47062 228453
rect 47146 228217 47382 228453
rect 46826 227897 47062 228133
rect 47146 227897 47382 228133
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 228217 83062 228453
rect 83146 228217 83382 228453
rect 82826 227897 83062 228133
rect 83146 227897 83382 228133
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 118826 228217 119062 228453
rect 119146 228217 119382 228453
rect 118826 227897 119062 228133
rect 119146 227897 119382 228133
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 136036 205625 136272 205861
rect 136356 205625 136592 205861
rect 136676 205625 136912 205861
rect 136996 205625 137232 205861
rect 137316 205625 137552 205861
rect 137636 205625 137872 205861
rect 137956 205625 138192 205861
rect 138276 205625 138512 205861
rect 138596 205625 138832 205861
rect 138916 205625 139152 205861
rect 139236 205625 139472 205861
rect 139556 205625 139792 205861
rect 139876 205625 140112 205861
rect 140196 205625 140432 205861
rect 140516 205625 140752 205861
rect 140836 205625 141072 205861
rect 141156 205625 141392 205861
rect 141476 205625 141712 205861
rect 141796 205625 142032 205861
rect 142116 205625 142352 205861
rect 142436 205625 142672 205861
rect 142756 205625 142992 205861
rect 143076 205625 143312 205861
rect 143396 205625 143632 205861
rect 143716 205625 143952 205861
rect 144036 205625 144272 205861
rect 144356 205625 144592 205861
rect 144676 205625 144912 205861
rect 144996 205625 145232 205861
rect 145316 205625 145552 205861
rect 145636 205625 145872 205861
rect 145956 205625 146192 205861
rect 146276 205625 146512 205861
rect 146596 205625 146832 205861
rect 146916 205625 147152 205861
rect 147236 205625 147472 205861
rect 147556 205625 147792 205861
rect 147876 205625 148112 205861
rect 148196 205625 148432 205861
rect 148516 205625 148752 205861
rect 148836 205625 149072 205861
rect 149156 205625 149392 205861
rect 149476 205625 149712 205861
rect 149796 205625 150032 205861
rect 150116 205625 150352 205861
rect 150436 205625 150672 205861
rect 150756 205625 150992 205861
rect 151076 205625 151312 205861
rect 151396 205625 151632 205861
rect 151716 205625 151952 205861
rect 152036 205625 152272 205861
rect 152356 205625 152592 205861
rect 152676 205625 152912 205861
rect 152996 205625 153232 205861
rect 153316 205625 153552 205861
rect 153636 205625 153872 205861
rect 153956 205625 154192 205861
rect 154276 205625 154512 205861
rect 154596 205625 154832 205861
rect 154916 205625 155152 205861
rect 155236 205625 155472 205861
rect 155556 205625 155792 205861
rect 155876 205625 156112 205861
rect 156196 205625 156432 205861
rect 156516 205625 156752 205861
rect 156836 205625 157072 205861
rect 157156 205625 157392 205861
rect 157476 205625 157712 205861
rect 157796 205625 158032 205861
rect 158116 205625 158352 205861
rect 158436 205625 158672 205861
rect 158756 205625 158992 205861
rect 159076 205625 159312 205861
rect 159396 205625 159632 205861
rect 159716 205625 159952 205861
rect 160036 205625 160272 205861
rect 160356 205625 160592 205861
rect 160676 205625 160912 205861
rect 160996 205625 161232 205861
rect 161316 205625 161552 205861
rect 161636 205625 161872 205861
rect 161956 205625 162192 205861
rect 162276 205625 162512 205861
rect 162596 205625 162832 205861
rect 162916 205625 163152 205861
rect 163236 205625 163472 205861
rect 163556 205625 163792 205861
rect 163876 205625 164112 205861
rect 164196 205625 164432 205861
rect 164516 205625 164752 205861
rect 164836 205625 165072 205861
rect 165156 205625 165392 205861
rect 137376 201175 137612 201411
rect 137696 201175 137932 201411
rect 138016 201175 138252 201411
rect 138336 201175 138572 201411
rect 138656 201175 138892 201411
rect 138976 201175 139212 201411
rect 139296 201175 139532 201411
rect 139616 201175 139852 201411
rect 139936 201175 140172 201411
rect 140256 201175 140492 201411
rect 140576 201175 140812 201411
rect 140896 201175 141132 201411
rect 141216 201175 141452 201411
rect 141536 201175 141772 201411
rect 141856 201175 142092 201411
rect 142176 201175 142412 201411
rect 142496 201175 142732 201411
rect 142816 201175 143052 201411
rect 143136 201175 143372 201411
rect 143456 201175 143692 201411
rect 143776 201175 144012 201411
rect 144096 201175 144332 201411
rect 144416 201175 144652 201411
rect 144736 201175 144972 201411
rect 145056 201175 145292 201411
rect 145376 201175 145612 201411
rect 145696 201175 145932 201411
rect 146016 201175 146252 201411
rect 146336 201175 146572 201411
rect 146656 201175 146892 201411
rect 146976 201175 147212 201411
rect 147296 201175 147532 201411
rect 147616 201175 147852 201411
rect 147936 201175 148172 201411
rect 148256 201175 148492 201411
rect 148576 201175 148812 201411
rect 148896 201175 149132 201411
rect 149216 201175 149452 201411
rect 149536 201175 149772 201411
rect 149856 201175 150092 201411
rect 150176 201175 150412 201411
rect 150496 201175 150732 201411
rect 150816 201175 151052 201411
rect 151136 201175 151372 201411
rect 151456 201175 151692 201411
rect 151776 201175 152012 201411
rect 152096 201175 152332 201411
rect 152416 201175 152652 201411
rect 152736 201175 152972 201411
rect 153056 201175 153292 201411
rect 153376 201175 153612 201411
rect 153696 201175 153932 201411
rect 154016 201175 154252 201411
rect 154336 201175 154572 201411
rect 154656 201175 154892 201411
rect 154976 201175 155212 201411
rect 155296 201175 155532 201411
rect 155616 201175 155852 201411
rect 155936 201175 156172 201411
rect 156256 201175 156492 201411
rect 156576 201175 156812 201411
rect 156896 201175 157132 201411
rect 157216 201175 157452 201411
rect 157536 201175 157772 201411
rect 157856 201175 158092 201411
rect 158176 201175 158412 201411
rect 158496 201175 158732 201411
rect 158816 201175 159052 201411
rect 159136 201175 159372 201411
rect 159456 201175 159692 201411
rect 159776 201175 160012 201411
rect 160096 201175 160332 201411
rect 160416 201175 160652 201411
rect 160736 201175 160972 201411
rect 161056 201175 161292 201411
rect 161376 201175 161612 201411
rect 161696 201175 161932 201411
rect 162016 201175 162252 201411
rect 162336 201175 162572 201411
rect 162656 201175 162892 201411
rect 162976 201175 163212 201411
rect 163296 201175 163532 201411
rect 163616 201175 163852 201411
rect 163936 201175 164172 201411
rect 164256 201175 164492 201411
rect 164576 201175 164812 201411
rect 164896 201175 165132 201411
rect 165216 201175 165452 201411
rect 137066 174218 137302 174454
rect 137386 174218 137622 174454
rect 137706 174218 137942 174454
rect 138026 174218 138262 174454
rect 138346 174218 138582 174454
rect 138666 174218 138902 174454
rect 138986 174218 139222 174454
rect 139306 174218 139542 174454
rect 139626 174218 139862 174454
rect 139946 174218 140182 174454
rect 140266 174218 140502 174454
rect 140586 174218 140822 174454
rect 140906 174218 141142 174454
rect 141226 174218 141462 174454
rect 137066 173898 137302 174134
rect 137386 173898 137622 174134
rect 137706 173898 137942 174134
rect 138026 173898 138262 174134
rect 138346 173898 138582 174134
rect 138666 173898 138902 174134
rect 138986 173898 139222 174134
rect 139306 173898 139542 174134
rect 139626 173898 139862 174134
rect 139946 173898 140182 174134
rect 140266 173898 140502 174134
rect 140586 173898 140822 174134
rect 140906 173898 141142 174134
rect 141226 173898 141462 174134
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 135610 115718 135846 115954
rect 135610 115398 135846 115634
rect 166330 115718 166566 115954
rect 166330 115398 166566 115634
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 120250 111218 120486 111454
rect 120250 110898 120486 111134
rect 150970 111218 151206 111454
rect 150970 110898 151206 111134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 135610 79718 135846 79954
rect 135610 79398 135846 79634
rect 166330 79718 166566 79954
rect 166330 79398 166566 79634
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 228217 191062 228453
rect 191146 228217 191382 228453
rect 190826 227897 191062 228133
rect 191146 227897 191382 228133
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 228217 227062 228453
rect 227146 228217 227382 228453
rect 226826 227897 227062 228133
rect 227146 227897 227382 228133
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 228217 263062 228453
rect 263146 228217 263382 228453
rect 262826 227897 263062 228133
rect 263146 227897 263382 228133
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 228217 299062 228453
rect 299146 228217 299382 228453
rect 298826 227897 299062 228133
rect 299146 227897 299382 228133
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 228217 335062 228453
rect 335146 228217 335382 228453
rect 334826 227897 335062 228133
rect 335146 227897 335382 228133
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 228217 371062 228453
rect 371146 228217 371382 228453
rect 370826 227897 371062 228133
rect 371146 227897 371382 228133
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 561342 318125 561578 318361
rect 561662 318125 561898 318361
rect 561982 318125 562218 318361
rect 562302 318125 562538 318361
rect 562622 318125 562858 318361
rect 562942 318125 563178 318361
rect 563262 318125 563498 318361
rect 563582 318125 563818 318361
rect 563902 318125 564138 318361
rect 564222 318125 564458 318361
rect 564542 318125 564778 318361
rect 564862 318125 565098 318361
rect 565182 318125 565418 318361
rect 565502 318125 565738 318361
rect 565822 318125 566058 318361
rect 561462 313718 561698 313954
rect 561782 313718 562018 313954
rect 562102 313718 562338 313954
rect 562422 313718 562658 313954
rect 562742 313718 562978 313954
rect 563062 313718 563298 313954
rect 563382 313718 563618 313954
rect 563702 313718 563938 313954
rect 564022 313718 564258 313954
rect 564342 313718 564578 313954
rect 564662 313718 564898 313954
rect 564982 313718 565218 313954
rect 565302 313718 565538 313954
rect 565622 313718 565858 313954
rect 565942 313718 566178 313954
rect 566262 313718 566498 313954
rect 566582 313718 566818 313954
rect 566902 313718 567138 313954
rect 561462 313398 561698 313634
rect 561782 313398 562018 313634
rect 562102 313398 562338 313634
rect 562422 313398 562658 313634
rect 562742 313398 562978 313634
rect 563062 313398 563298 313634
rect 563382 313398 563618 313634
rect 563702 313398 563938 313634
rect 564022 313398 564258 313634
rect 564342 313398 564578 313634
rect 564662 313398 564898 313634
rect 564982 313398 565218 313634
rect 565302 313398 565538 313634
rect 565622 313398 565858 313634
rect 565942 313398 566178 313634
rect 566262 313398 566498 313634
rect 566582 313398 566818 313634
rect 566902 313398 567138 313634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318361 591102 318454
rect 533382 318218 561342 318361
rect -8726 318134 561342 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 318125 561342 318134
rect 561578 318125 561662 318361
rect 561898 318125 561982 318361
rect 562218 318125 562302 318361
rect 562538 318125 562622 318361
rect 562858 318125 562942 318361
rect 563178 318125 563262 318361
rect 563498 318125 563582 318361
rect 563818 318125 563902 318361
rect 564138 318125 564222 318361
rect 564458 318125 564542 318361
rect 564778 318125 564862 318361
rect 565098 318125 565182 318361
rect 565418 318125 565502 318361
rect 565738 318125 565822 318361
rect 566058 318218 591102 318361
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect 566058 318134 592650 318218
rect 566058 318125 591102 318134
rect 533382 317898 591102 318125
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 561462 313954
rect 561698 313718 561782 313954
rect 562018 313718 562102 313954
rect 562338 313718 562422 313954
rect 562658 313718 562742 313954
rect 562978 313718 563062 313954
rect 563298 313718 563382 313954
rect 563618 313718 563702 313954
rect 563938 313718 564022 313954
rect 564258 313718 564342 313954
rect 564578 313718 564662 313954
rect 564898 313718 564982 313954
rect 565218 313718 565302 313954
rect 565538 313718 565622 313954
rect 565858 313718 565942 313954
rect 566178 313718 566262 313954
rect 566498 313718 566582 313954
rect 566818 313718 566902 313954
rect 567138 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 561462 313634
rect 561698 313398 561782 313634
rect 562018 313398 562102 313634
rect 562338 313398 562422 313634
rect 562658 313398 562742 313634
rect 562978 313398 563062 313634
rect 563298 313398 563382 313634
rect 563618 313398 563702 313634
rect 563938 313398 564022 313634
rect 564258 313398 564342 313634
rect 564578 313398 564662 313634
rect 564898 313398 564982 313634
rect 565218 313398 565302 313634
rect 565538 313398 565622 313634
rect 565858 313398 565942 313634
rect 566178 313398 566262 313634
rect 566498 313398 566582 313634
rect 566818 313398 566902 313634
rect 567138 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246303 424826 246454
rect 29382 246218 65342 246303
rect -8726 246134 65342 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 246067 65342 246134
rect 65578 246067 65662 246303
rect 65898 246067 65982 246303
rect 66218 246067 66302 246303
rect 66538 246067 66622 246303
rect 66858 246067 66942 246303
rect 67178 246067 67262 246303
rect 67498 246067 67582 246303
rect 67818 246067 67902 246303
rect 68138 246067 68222 246303
rect 68458 246067 68542 246303
rect 68778 246067 68862 246303
rect 69098 246067 69182 246303
rect 69418 246067 69502 246303
rect 69738 246067 69822 246303
rect 70058 246218 424826 246303
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect 70058 246134 592650 246218
rect 70058 246067 424826 246134
rect 29382 245898 424826 246067
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241953 420326 241954
rect 24882 241718 65462 241953
rect -8726 241717 65462 241718
rect 65698 241717 65782 241953
rect 66018 241717 66102 241953
rect 66338 241717 66422 241953
rect 66658 241717 66742 241953
rect 66978 241717 67062 241953
rect 67298 241717 67382 241953
rect 67618 241717 67702 241953
rect 67938 241717 68022 241953
rect 68258 241717 68342 241953
rect 68578 241717 68662 241953
rect 68898 241717 68982 241953
rect 69218 241717 69302 241953
rect 69538 241717 69622 241953
rect 69858 241717 69942 241953
rect 70178 241717 70262 241953
rect 70498 241717 70582 241953
rect 70818 241717 70902 241953
rect 71138 241718 420326 241953
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect 71138 241717 592650 241718
rect -8726 241634 592650 241717
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241633 420326 241634
rect 24882 241398 65462 241633
rect -8726 241397 65462 241398
rect 65698 241397 65782 241633
rect 66018 241397 66102 241633
rect 66338 241397 66422 241633
rect 66658 241397 66742 241633
rect 66978 241397 67062 241633
rect 67298 241397 67382 241633
rect 67618 241397 67702 241633
rect 67938 241397 68022 241633
rect 68258 241397 68342 241633
rect 68578 241397 68662 241633
rect 68898 241397 68982 241633
rect 69218 241397 69302 241633
rect 69538 241397 69622 241633
rect 69858 241397 69942 241633
rect 70178 241397 70262 241633
rect 70498 241397 70582 241633
rect 70818 241397 70902 241633
rect 71138 241398 420326 241633
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect 71138 241397 592650 241398
rect -8726 241366 592650 241397
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228453 406826 228454
rect 11382 228218 46826 228453
rect -8726 228217 46826 228218
rect 47062 228217 47146 228453
rect 47382 228217 82826 228453
rect 83062 228217 83146 228453
rect 83382 228217 118826 228453
rect 119062 228217 119146 228453
rect 119382 228217 190826 228453
rect 191062 228217 191146 228453
rect 191382 228217 226826 228453
rect 227062 228217 227146 228453
rect 227382 228217 262826 228453
rect 263062 228217 263146 228453
rect 263382 228217 298826 228453
rect 299062 228217 299146 228453
rect 299382 228217 334826 228453
rect 335062 228217 335146 228453
rect 335382 228217 370826 228453
rect 371062 228217 371146 228453
rect 371382 228218 406826 228453
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect 371382 228217 592650 228218
rect -8726 228134 592650 228217
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 228133 406826 228134
rect 11382 227898 46826 228133
rect -8726 227897 46826 227898
rect 47062 227897 47146 228133
rect 47382 227897 82826 228133
rect 83062 227897 83146 228133
rect 83382 227897 118826 228133
rect 119062 227897 119146 228133
rect 119382 227897 190826 228133
rect 191062 227897 191146 228133
rect 191382 227897 226826 228133
rect 227062 227897 227146 228133
rect 227382 227897 262826 228133
rect 263062 227897 263146 228133
rect 263382 227897 298826 228133
rect 299062 227897 299146 228133
rect 299382 227897 334826 228133
rect 335062 227897 335146 228133
rect 335382 227897 370826 228133
rect 371062 227897 371146 228133
rect 371382 227898 406826 228133
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect 371382 227897 592650 227898
rect -8726 227866 592650 227897
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205861 204326 205954
rect 132882 205718 136036 205861
rect -8726 205634 136036 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205625 136036 205634
rect 136272 205625 136356 205861
rect 136592 205625 136676 205861
rect 136912 205625 136996 205861
rect 137232 205625 137316 205861
rect 137552 205625 137636 205861
rect 137872 205625 137956 205861
rect 138192 205625 138276 205861
rect 138512 205625 138596 205861
rect 138832 205625 138916 205861
rect 139152 205625 139236 205861
rect 139472 205625 139556 205861
rect 139792 205625 139876 205861
rect 140112 205625 140196 205861
rect 140432 205625 140516 205861
rect 140752 205625 140836 205861
rect 141072 205625 141156 205861
rect 141392 205625 141476 205861
rect 141712 205625 141796 205861
rect 142032 205625 142116 205861
rect 142352 205625 142436 205861
rect 142672 205625 142756 205861
rect 142992 205625 143076 205861
rect 143312 205625 143396 205861
rect 143632 205625 143716 205861
rect 143952 205625 144036 205861
rect 144272 205625 144356 205861
rect 144592 205625 144676 205861
rect 144912 205625 144996 205861
rect 145232 205625 145316 205861
rect 145552 205625 145636 205861
rect 145872 205625 145956 205861
rect 146192 205625 146276 205861
rect 146512 205625 146596 205861
rect 146832 205625 146916 205861
rect 147152 205625 147236 205861
rect 147472 205625 147556 205861
rect 147792 205625 147876 205861
rect 148112 205625 148196 205861
rect 148432 205625 148516 205861
rect 148752 205625 148836 205861
rect 149072 205625 149156 205861
rect 149392 205625 149476 205861
rect 149712 205625 149796 205861
rect 150032 205625 150116 205861
rect 150352 205625 150436 205861
rect 150672 205625 150756 205861
rect 150992 205625 151076 205861
rect 151312 205625 151396 205861
rect 151632 205625 151716 205861
rect 151952 205625 152036 205861
rect 152272 205625 152356 205861
rect 152592 205625 152676 205861
rect 152912 205625 152996 205861
rect 153232 205625 153316 205861
rect 153552 205625 153636 205861
rect 153872 205625 153956 205861
rect 154192 205625 154276 205861
rect 154512 205625 154596 205861
rect 154832 205625 154916 205861
rect 155152 205625 155236 205861
rect 155472 205625 155556 205861
rect 155792 205625 155876 205861
rect 156112 205625 156196 205861
rect 156432 205625 156516 205861
rect 156752 205625 156836 205861
rect 157072 205625 157156 205861
rect 157392 205625 157476 205861
rect 157712 205625 157796 205861
rect 158032 205625 158116 205861
rect 158352 205625 158436 205861
rect 158672 205625 158756 205861
rect 158992 205625 159076 205861
rect 159312 205625 159396 205861
rect 159632 205625 159716 205861
rect 159952 205625 160036 205861
rect 160272 205625 160356 205861
rect 160592 205625 160676 205861
rect 160912 205625 160996 205861
rect 161232 205625 161316 205861
rect 161552 205625 161636 205861
rect 161872 205625 161956 205861
rect 162192 205625 162276 205861
rect 162512 205625 162596 205861
rect 162832 205625 162916 205861
rect 163152 205625 163236 205861
rect 163472 205625 163556 205861
rect 163792 205625 163876 205861
rect 164112 205625 164196 205861
rect 164432 205625 164516 205861
rect 164752 205625 164836 205861
rect 165072 205625 165156 205861
rect 165392 205718 204326 205861
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect 165392 205634 592650 205718
rect 165392 205625 204326 205634
rect 132882 205398 204326 205625
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201411 199826 201454
rect 128382 201218 137376 201411
rect -8726 201175 137376 201218
rect 137612 201175 137696 201411
rect 137932 201175 138016 201411
rect 138252 201175 138336 201411
rect 138572 201175 138656 201411
rect 138892 201175 138976 201411
rect 139212 201175 139296 201411
rect 139532 201175 139616 201411
rect 139852 201175 139936 201411
rect 140172 201175 140256 201411
rect 140492 201175 140576 201411
rect 140812 201175 140896 201411
rect 141132 201175 141216 201411
rect 141452 201175 141536 201411
rect 141772 201175 141856 201411
rect 142092 201175 142176 201411
rect 142412 201175 142496 201411
rect 142732 201175 142816 201411
rect 143052 201175 143136 201411
rect 143372 201175 143456 201411
rect 143692 201175 143776 201411
rect 144012 201175 144096 201411
rect 144332 201175 144416 201411
rect 144652 201175 144736 201411
rect 144972 201175 145056 201411
rect 145292 201175 145376 201411
rect 145612 201175 145696 201411
rect 145932 201175 146016 201411
rect 146252 201175 146336 201411
rect 146572 201175 146656 201411
rect 146892 201175 146976 201411
rect 147212 201175 147296 201411
rect 147532 201175 147616 201411
rect 147852 201175 147936 201411
rect 148172 201175 148256 201411
rect 148492 201175 148576 201411
rect 148812 201175 148896 201411
rect 149132 201175 149216 201411
rect 149452 201175 149536 201411
rect 149772 201175 149856 201411
rect 150092 201175 150176 201411
rect 150412 201175 150496 201411
rect 150732 201175 150816 201411
rect 151052 201175 151136 201411
rect 151372 201175 151456 201411
rect 151692 201175 151776 201411
rect 152012 201175 152096 201411
rect 152332 201175 152416 201411
rect 152652 201175 152736 201411
rect 152972 201175 153056 201411
rect 153292 201175 153376 201411
rect 153612 201175 153696 201411
rect 153932 201175 154016 201411
rect 154252 201175 154336 201411
rect 154572 201175 154656 201411
rect 154892 201175 154976 201411
rect 155212 201175 155296 201411
rect 155532 201175 155616 201411
rect 155852 201175 155936 201411
rect 156172 201175 156256 201411
rect 156492 201175 156576 201411
rect 156812 201175 156896 201411
rect 157132 201175 157216 201411
rect 157452 201175 157536 201411
rect 157772 201175 157856 201411
rect 158092 201175 158176 201411
rect 158412 201175 158496 201411
rect 158732 201175 158816 201411
rect 159052 201175 159136 201411
rect 159372 201175 159456 201411
rect 159692 201175 159776 201411
rect 160012 201175 160096 201411
rect 160332 201175 160416 201411
rect 160652 201175 160736 201411
rect 160972 201175 161056 201411
rect 161292 201175 161376 201411
rect 161612 201175 161696 201411
rect 161932 201175 162016 201411
rect 162252 201175 162336 201411
rect 162572 201175 162656 201411
rect 162892 201175 162976 201411
rect 163212 201175 163296 201411
rect 163532 201175 163616 201411
rect 163852 201175 163936 201411
rect 164172 201175 164256 201411
rect 164492 201175 164576 201411
rect 164812 201175 164896 201411
rect 165132 201175 165216 201411
rect 165452 201218 199826 201411
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect 165452 201175 592650 201218
rect -8726 201134 592650 201175
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 137066 174454
rect 137302 174218 137386 174454
rect 137622 174218 137706 174454
rect 137942 174218 138026 174454
rect 138262 174218 138346 174454
rect 138582 174218 138666 174454
rect 138902 174218 138986 174454
rect 139222 174218 139306 174454
rect 139542 174218 139626 174454
rect 139862 174218 139946 174454
rect 140182 174218 140266 174454
rect 140502 174218 140586 174454
rect 140822 174218 140906 174454
rect 141142 174218 141226 174454
rect 141462 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 137066 174134
rect 137302 173898 137386 174134
rect 137622 173898 137706 174134
rect 137942 173898 138026 174134
rect 138262 173898 138346 174134
rect 138582 173898 138666 174134
rect 138902 173898 138986 174134
rect 139222 173898 139306 174134
rect 139542 173898 139626 174134
rect 139862 173898 139946 174134
rect 140182 173898 140266 174134
rect 140502 173898 140586 174134
rect 140822 173898 140906 174134
rect 141142 173898 141226 174134
rect 141462 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 135610 115954
rect 135846 115718 166330 115954
rect 166566 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 135610 115634
rect 135846 115398 166330 115634
rect 166566 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 120250 111454
rect 120486 111218 150970 111454
rect 151206 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 120250 111134
rect 120486 110898 150970 111134
rect 151206 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 135610 79954
rect 135846 79718 166330 79954
rect 166566 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 135610 79634
rect 135846 79398 166330 79634
rect 166566 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use APS  APS_macro0
timestamp 0
transform 1 0 512000 0 1 304600
box 30000 -2600 55300 14200
use PD_M1_M2  PD_M1_M2_macro0
timestamp 0
transform 1 0 16000 0 1 232484
box 30000 -2000 380500 14200
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 116000 0 1 75000
box 0 0 60000 60000
use SystemLevel  sl_macro0
timestamp 0
transform 1 0 148914 0 1 188300
box -13000 -15200 17500 18000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 248684 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 248684 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 73000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 248684 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 248684 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 248684 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 248684 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 248684 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 248684 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 248684 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 248684 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 300000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 320800 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 248684 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 248684 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 73000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 137000 119414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 248684 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 73000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 248684 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 248684 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 248684 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 248684 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 248684 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 248684 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 248684 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 300000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 320800 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 248684 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 248684 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 73000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 137000 128414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 248684 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 73000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 248684 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 248684 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 248684 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 248684 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 248684 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 248684 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 248684 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 300000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 320800 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 248684 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 248684 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 73000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 248684 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 73000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 137000 173414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 248684 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 248684 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 248684 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 248684 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 248684 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 248684 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 248684 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 300000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 320800 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 248684 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 248684 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 73000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 137000 132914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 248684 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 73000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 248684 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 248684 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 248684 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 248684 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 248684 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 248684 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 248684 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 300000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 320800 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 248684 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 248684 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 73000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 248684 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 73000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 137000 177914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 248684 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 248684 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 248684 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 248684 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 248684 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 248684 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 248684 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 248684 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 73000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 137000 114914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 248684 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 73000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 248684 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 248684 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 248684 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 248684 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 248684 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 248684 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 248684 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 300000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 320800 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 248684 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 248684 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 73000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 137000 123914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 248684 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 73000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 248684 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 248684 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 248684 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 248684 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 248684 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 248684 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 248684 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 300000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 320800 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
